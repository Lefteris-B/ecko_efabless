magic
tech sky130A
magscale 1 2
timestamp 1715980349
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 934 2128 68894 67504
<< metal2 >>
rect 3882 69200 3938 70000
rect 12898 69200 12954 70000
rect 21270 69200 21326 70000
rect 30286 69200 30342 70000
rect 39302 69200 39358 70000
rect 47674 69200 47730 70000
rect 56690 69200 56746 70000
rect 65706 69200 65762 70000
rect 18 0 74 800
rect 8390 0 8446 800
rect 17406 0 17462 800
rect 26422 0 26478 800
rect 34794 0 34850 800
rect 43810 0 43866 800
rect 52826 0 52882 800
rect 61198 0 61254 800
<< obsm2 >>
rect 938 69144 3826 69306
rect 3994 69144 12842 69306
rect 13010 69144 21214 69306
rect 21382 69144 30230 69306
rect 30398 69144 39246 69306
rect 39414 69144 47618 69306
rect 47786 69144 56634 69306
rect 56802 69144 65650 69306
rect 65818 69144 68890 69306
rect 938 856 68890 69144
rect 938 31 8334 856
rect 8502 31 17350 856
rect 17518 31 26366 856
rect 26534 31 34738 856
rect 34906 31 43754 856
rect 43922 31 52770 856
rect 52938 31 61142 856
rect 61310 31 68890 856
<< metal3 >>
rect 69200 65288 70000 65408
rect 0 64608 800 64728
rect 0 55768 800 55888
rect 69200 55768 70000 55888
rect 0 46248 800 46368
rect 69200 46248 70000 46368
rect 69200 37408 70000 37528
rect 0 36728 800 36848
rect 0 27888 800 28008
rect 69200 27888 70000 28008
rect 0 18368 800 18488
rect 69200 18368 70000 18488
rect 69200 9528 70000 9648
rect 0 8848 800 8968
rect 69200 8 70000 128
<< obsm3 >>
rect 798 65488 69200 67489
rect 798 65208 69120 65488
rect 798 64808 69200 65208
rect 880 64528 69200 64808
rect 798 55968 69200 64528
rect 880 55688 69120 55968
rect 798 46448 69200 55688
rect 880 46168 69120 46448
rect 798 37608 69200 46168
rect 798 37328 69120 37608
rect 798 36928 69200 37328
rect 880 36648 69200 36928
rect 798 28088 69200 36648
rect 880 27808 69120 28088
rect 798 18568 69200 27808
rect 880 18288 69120 18568
rect 798 9728 69200 18288
rect 798 9448 69120 9728
rect 798 9048 69200 9448
rect 880 8768 69200 9048
rect 798 208 69200 8768
rect 798 35 69120 208
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< labels >>
rlabel metal3 s 69200 46248 70000 46368 6 audio_sample[0]
port 1 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 audio_sample[10]
port 2 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 audio_sample[11]
port 3 nsew signal input
rlabel metal3 s 69200 37408 70000 37528 6 audio_sample[12]
port 4 nsew signal input
rlabel metal2 s 47674 69200 47730 70000 6 audio_sample[13]
port 5 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 audio_sample[14]
port 6 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 audio_sample[15]
port 7 nsew signal input
rlabel metal3 s 69200 65288 70000 65408 6 audio_sample[1]
port 8 nsew signal input
rlabel metal2 s 56690 69200 56746 70000 6 audio_sample[2]
port 9 nsew signal input
rlabel metal3 s 69200 18368 70000 18488 6 audio_sample[3]
port 10 nsew signal input
rlabel metal2 s 18 0 74 800 6 audio_sample[4]
port 11 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 audio_sample[5]
port 12 nsew signal input
rlabel metal2 s 65706 69200 65762 70000 6 audio_sample[6]
port 13 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 audio_sample[7]
port 14 nsew signal input
rlabel metal2 s 21270 69200 21326 70000 6 audio_sample[8]
port 15 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 audio_sample[9]
port 16 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 clk
port 17 nsew signal input
rlabel metal3 s 69200 8 70000 128 6 done
port 18 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 psram_ce_n
port 19 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 psram_d[0]
port 20 nsew signal bidirectional
rlabel metal2 s 12898 69200 12954 70000 6 psram_d[1]
port 21 nsew signal bidirectional
rlabel metal3 s 69200 9528 70000 9648 6 psram_d[2]
port 22 nsew signal bidirectional
rlabel metal2 s 26422 0 26478 800 6 psram_d[3]
port 23 nsew signal bidirectional
rlabel metal3 s 0 64608 800 64728 6 psram_douten[0]
port 24 nsew signal output
rlabel metal3 s 69200 55768 70000 55888 6 psram_douten[1]
port 25 nsew signal output
rlabel metal2 s 30286 69200 30342 70000 6 psram_douten[2]
port 26 nsew signal output
rlabel metal2 s 39302 69200 39358 70000 6 psram_douten[3]
port 27 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 psram_sck
port 28 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 rst
port 29 nsew signal input
rlabel metal2 s 3882 69200 3938 70000 6 sample_valid
port 30 nsew signal input
rlabel metal3 s 69200 27888 70000 28008 6 start
port 31 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 33 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3412756
string GDS_FILE /home/iamme/asic_tools/caravel_user_project/openlane/cnn_kws_accel/runs/24_05_17_23_52/results/signoff/cnn_kws_accel.magic.gds
string GDS_START 483518
<< end >>

