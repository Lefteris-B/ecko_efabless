VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cnn_kws_accel
  CLASS BLOCK ;
  FOREIGN cnn_kws_accel ;
  ORIGIN 0.000 0.000 ;
  SIZE 138.205 BY 148.925 ;
  PIN audio_sample[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.205 98.640 138.205 99.240 ;
    END
  END audio_sample[0]
  PIN audio_sample[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END audio_sample[10]
  PIN audio_sample[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END audio_sample[11]
  PIN audio_sample[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.205 81.640 138.205 82.240 ;
    END
  END audio_sample[12]
  PIN audio_sample[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 144.925 90.530 148.925 ;
    END
  END audio_sample[13]
  PIN audio_sample[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END audio_sample[14]
  PIN audio_sample[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END audio_sample[15]
  PIN audio_sample[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.205 139.440 138.205 140.040 ;
    END
  END audio_sample[1]
  PIN audio_sample[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 144.925 109.850 148.925 ;
    END
  END audio_sample[2]
  PIN audio_sample[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.205 44.240 138.205 44.840 ;
    END
  END audio_sample[3]
  PIN audio_sample[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END audio_sample[4]
  PIN audio_sample[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END audio_sample[5]
  PIN audio_sample[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 144.925 129.170 148.925 ;
    END
  END audio_sample[6]
  PIN audio_sample[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END audio_sample[7]
  PIN audio_sample[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 144.925 39.010 148.925 ;
    END
  END audio_sample[8]
  PIN audio_sample[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END audio_sample[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 134.205 3.440 138.205 4.040 ;
    END
  END done
  PIN psram_ce_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END psram_ce_n
  PIN psram_d[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.484000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END psram_d[0]
  PIN psram_d[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 144.925 19.690 148.925 ;
    END
  END psram_d[1]
  PIN psram_d[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.205 23.840 138.205 24.440 ;
    END
  END psram_d[2]
  PIN psram_d[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END psram_d[3]
  PIN psram_douten[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END psram_douten[0]
  PIN psram_douten[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.205 119.040 138.205 119.640 ;
    END
  END psram_douten[1]
  PIN psram_douten[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 144.925 55.110 148.925 ;
    END
  END psram_douten[2]
  PIN psram_douten[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 144.925 74.430 148.925 ;
    END
  END psram_douten[3]
  PIN psram_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END psram_sck
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END rst_n
  PIN sample_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 144.925 0.370 148.925 ;
    END
  END sample_valid
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 134.205 61.240 138.205 61.840 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.590 10.640 22.190 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 52.330 10.640 53.930 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.070 10.640 85.670 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.810 10.640 117.410 136.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 36.460 10.640 38.060 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.200 10.640 69.800 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.940 10.640 101.540 136.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.680 10.640 133.280 136.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 132.480 136.085 ;
      LAYER met1 ;
        RECT 4.670 10.640 133.280 136.240 ;
      LAYER met2 ;
        RECT 4.690 144.645 19.130 144.925 ;
        RECT 19.970 144.645 38.450 144.925 ;
        RECT 39.290 144.645 54.550 144.925 ;
        RECT 55.390 144.645 73.870 144.925 ;
        RECT 74.710 144.645 89.970 144.925 ;
        RECT 90.810 144.645 109.290 144.925 ;
        RECT 110.130 144.645 128.610 144.925 ;
        RECT 129.450 144.645 133.250 144.925 ;
        RECT 4.690 4.280 133.250 144.645 ;
        RECT 4.690 3.555 15.910 4.280 ;
        RECT 16.750 3.555 35.230 4.280 ;
        RECT 36.070 3.555 51.330 4.280 ;
        RECT 52.170 3.555 70.650 4.280 ;
        RECT 71.490 3.555 89.970 4.280 ;
        RECT 90.810 3.555 106.070 4.280 ;
        RECT 106.910 3.555 125.390 4.280 ;
        RECT 126.230 3.555 133.250 4.280 ;
      LAYER met3 ;
        RECT 3.990 133.640 134.930 136.165 ;
        RECT 4.400 132.240 134.930 133.640 ;
        RECT 3.990 120.040 134.930 132.240 ;
        RECT 3.990 118.640 133.805 120.040 ;
        RECT 3.990 113.240 134.930 118.640 ;
        RECT 4.400 111.840 134.930 113.240 ;
        RECT 3.990 99.640 134.930 111.840 ;
        RECT 3.990 98.240 133.805 99.640 ;
        RECT 3.990 96.240 134.930 98.240 ;
        RECT 4.400 94.840 134.930 96.240 ;
        RECT 3.990 82.640 134.930 94.840 ;
        RECT 3.990 81.240 133.805 82.640 ;
        RECT 3.990 75.840 134.930 81.240 ;
        RECT 4.400 74.440 134.930 75.840 ;
        RECT 3.990 62.240 134.930 74.440 ;
        RECT 3.990 60.840 133.805 62.240 ;
        RECT 3.990 55.440 134.930 60.840 ;
        RECT 4.400 54.040 134.930 55.440 ;
        RECT 3.990 45.240 134.930 54.040 ;
        RECT 3.990 43.840 133.805 45.240 ;
        RECT 3.990 38.440 134.930 43.840 ;
        RECT 4.400 37.040 134.930 38.440 ;
        RECT 3.990 24.840 134.930 37.040 ;
        RECT 3.990 23.440 133.805 24.840 ;
        RECT 3.990 18.040 134.930 23.440 ;
        RECT 4.400 16.640 134.930 18.040 ;
        RECT 3.990 4.440 134.930 16.640 ;
        RECT 3.990 3.575 133.805 4.440 ;
  END
END cnn_kws_accel
END LIBRARY

