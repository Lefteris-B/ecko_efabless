magic
tech sky130A
magscale 1 2
timestamp 1715939643
<< viali >>
rect 56149 67337 56183 67371
rect 1593 67201 1627 67235
rect 2237 67201 2271 67235
rect 4813 67201 4847 67235
rect 7389 67201 7423 67235
rect 9965 67201 9999 67235
rect 12541 67201 12575 67235
rect 15117 67201 15151 67235
rect 17693 67201 17727 67235
rect 20269 67201 20303 67235
rect 22845 67201 22879 67235
rect 25421 67201 25455 67235
rect 27997 67201 28031 67235
rect 30573 67201 30607 67235
rect 33149 67201 33183 67235
rect 38301 67201 38335 67235
rect 40877 67201 40911 67235
rect 46029 67201 46063 67235
rect 53757 67201 53791 67235
rect 58909 67201 58943 67235
rect 61485 67201 61519 67235
rect 64061 67201 64095 67235
rect 68477 67201 68511 67235
rect 68477 65977 68511 66011
rect 1593 64889 1627 64923
rect 68477 63325 68511 63359
rect 67833 60673 67867 60707
rect 68201 60673 68235 60707
rect 68385 60537 68419 60571
rect 1593 59381 1627 59415
rect 68477 57885 68511 57919
rect 1593 56797 1627 56831
rect 68477 55097 68511 55131
rect 68477 52445 68511 52479
rect 1593 51357 1627 51391
rect 68477 49725 68511 49759
rect 1593 48501 1627 48535
rect 68477 47005 68511 47039
rect 1593 45917 1627 45951
rect 68477 44217 68511 44251
rect 1593 43061 1627 43095
rect 68477 41565 68511 41599
rect 1593 37621 1627 37655
rect 68477 36125 68511 36159
rect 1593 35037 1627 35071
rect 68293 33473 68327 33507
rect 68385 33269 68419 33303
rect 1593 32181 1627 32215
rect 68477 30685 68511 30719
rect 1593 29597 1627 29631
rect 68477 27897 68511 27931
rect 1593 26741 1627 26775
rect 28733 25245 28767 25279
rect 28917 25245 28951 25279
rect 31217 25245 31251 25279
rect 68477 25245 68511 25279
rect 28825 25109 28859 25143
rect 31769 25109 31803 25143
rect 31401 24905 31435 24939
rect 28448 24837 28482 24871
rect 30288 24769 30322 24803
rect 33977 24769 34011 24803
rect 34244 24769 34278 24803
rect 35449 24769 35483 24803
rect 35716 24769 35750 24803
rect 28181 24701 28215 24735
rect 30021 24701 30055 24735
rect 37289 24701 37323 24735
rect 29561 24565 29595 24599
rect 35357 24565 35391 24599
rect 36829 24565 36863 24599
rect 37933 24565 37967 24599
rect 28825 24361 28859 24395
rect 30297 24361 30331 24395
rect 33241 24361 33275 24395
rect 36001 24293 36035 24327
rect 30665 24225 30699 24259
rect 31217 24225 31251 24259
rect 31861 24225 31895 24259
rect 35357 24225 35391 24259
rect 36369 24225 36403 24259
rect 1593 24157 1627 24191
rect 29009 24157 29043 24191
rect 29101 24157 29135 24191
rect 29561 24157 29595 24191
rect 30481 24157 30515 24191
rect 30573 24157 30607 24191
rect 30757 24157 30791 24191
rect 36093 24157 36127 24191
rect 36185 24157 36219 24191
rect 36737 24157 36771 24191
rect 37381 24157 37415 24191
rect 28825 24089 28859 24123
rect 30205 24089 30239 24123
rect 32106 24089 32140 24123
rect 37648 24089 37682 24123
rect 31769 24021 31803 24055
rect 36369 24021 36403 24055
rect 37289 24021 37323 24055
rect 38761 24021 38795 24055
rect 30389 23817 30423 23851
rect 36185 23817 36219 23851
rect 36737 23817 36771 23851
rect 28365 23749 28399 23783
rect 28825 23749 28859 23783
rect 29561 23749 29595 23783
rect 31125 23749 31159 23783
rect 31309 23749 31343 23783
rect 34253 23749 34287 23783
rect 34469 23749 34503 23783
rect 36921 23749 36955 23783
rect 38025 23749 38059 23783
rect 38255 23715 38289 23749
rect 27169 23681 27203 23715
rect 28273 23681 28307 23715
rect 28457 23681 28491 23715
rect 28595 23681 28629 23715
rect 29009 23681 29043 23715
rect 29193 23681 29227 23715
rect 29285 23681 29319 23715
rect 29377 23681 29411 23715
rect 29653 23681 29687 23715
rect 30573 23681 30607 23715
rect 31033 23681 31067 23715
rect 31217 23681 31251 23715
rect 31493 23681 31527 23715
rect 31769 23681 31803 23715
rect 32321 23681 32355 23715
rect 32597 23681 32631 23715
rect 32781 23681 32815 23715
rect 34897 23681 34931 23715
rect 35173 23681 35207 23715
rect 35357 23681 35391 23715
rect 36093 23681 36127 23715
rect 36277 23681 36311 23715
rect 36829 23681 36863 23715
rect 38844 23681 38878 23715
rect 46673 23681 46707 23715
rect 28733 23613 28767 23647
rect 30849 23613 30883 23647
rect 32137 23613 32171 23647
rect 34713 23613 34747 23647
rect 35449 23613 35483 23647
rect 35633 23613 35667 23647
rect 35725 23613 35759 23647
rect 35817 23613 35851 23647
rect 35909 23613 35943 23647
rect 36553 23613 36587 23647
rect 37381 23613 37415 23647
rect 38577 23613 38611 23647
rect 46029 23613 46063 23647
rect 29469 23545 29503 23579
rect 32597 23545 32631 23579
rect 34621 23545 34655 23579
rect 26985 23477 27019 23511
rect 28089 23477 28123 23511
rect 30757 23477 30791 23511
rect 31677 23477 31711 23511
rect 32505 23477 32539 23511
rect 34437 23477 34471 23511
rect 37105 23477 37139 23511
rect 37933 23477 37967 23511
rect 38209 23477 38243 23511
rect 38393 23477 38427 23511
rect 39957 23477 39991 23511
rect 46581 23477 46615 23511
rect 46765 23477 46799 23511
rect 29101 23273 29135 23307
rect 31033 23273 31067 23307
rect 35081 23273 35115 23307
rect 36461 23273 36495 23307
rect 37013 23273 37047 23307
rect 37289 23273 37323 23307
rect 37749 23273 37783 23307
rect 39313 23273 39347 23307
rect 27997 23205 28031 23239
rect 31217 23205 31251 23239
rect 32045 23205 32079 23239
rect 37841 23205 37875 23239
rect 38301 23205 38335 23239
rect 28733 23137 28767 23171
rect 28825 23137 28859 23171
rect 31861 23137 31895 23171
rect 32413 23137 32447 23171
rect 34437 23137 34471 23171
rect 35173 23137 35207 23171
rect 36001 23137 36035 23171
rect 36093 23137 36127 23171
rect 36829 23137 36863 23171
rect 38485 23137 38519 23171
rect 38577 23137 38611 23171
rect 45569 23137 45603 23171
rect 47685 23137 47719 23171
rect 26617 23069 26651 23103
rect 28917 23069 28951 23103
rect 29101 23069 29135 23103
rect 29285 23069 29319 23103
rect 29561 23069 29595 23103
rect 29653 23069 29687 23103
rect 29837 23069 29871 23103
rect 30205 23069 30239 23103
rect 30941 23069 30975 23103
rect 31033 23069 31067 23103
rect 31493 23069 31527 23103
rect 31677 23069 31711 23103
rect 32321 23069 32355 23103
rect 34345 23069 34379 23103
rect 34529 23069 34563 23103
rect 34897 23069 34931 23103
rect 35449 23069 35483 23103
rect 36277 23063 36311 23097
rect 36645 23069 36679 23103
rect 37013 23069 37047 23103
rect 37749 23069 37783 23103
rect 38209 23069 38243 23103
rect 39589 23069 39623 23103
rect 45017 23069 45051 23103
rect 49525 23069 49559 23103
rect 26884 23001 26918 23035
rect 30021 23001 30055 23035
rect 30113 23001 30147 23035
rect 30573 23001 30607 23035
rect 31309 23001 31343 23035
rect 32045 23001 32079 23035
rect 32229 23001 32263 23035
rect 32680 23001 32714 23035
rect 37105 23001 37139 23035
rect 37321 23001 37355 23035
rect 38025 23001 38059 23035
rect 38485 23001 38519 23035
rect 39313 23001 39347 23035
rect 45845 23001 45879 23035
rect 47961 23001 47995 23035
rect 49617 23001 49651 23035
rect 28549 22933 28583 22967
rect 30389 22933 30423 22967
rect 31585 22933 31619 22967
rect 33793 22933 33827 22967
rect 34713 22933 34747 22967
rect 36737 22933 36771 22967
rect 37473 22933 37507 22967
rect 39221 22933 39255 22967
rect 39497 22933 39531 22967
rect 45109 22933 45143 22967
rect 47317 22933 47351 22967
rect 49433 22933 49467 22967
rect 27353 22729 27387 22763
rect 31693 22729 31727 22763
rect 32965 22729 32999 22763
rect 35449 22729 35483 22763
rect 46029 22729 46063 22763
rect 46397 22729 46431 22763
rect 31493 22661 31527 22695
rect 38853 22661 38887 22695
rect 46489 22661 46523 22695
rect 27169 22593 27203 22627
rect 30297 22593 30331 22627
rect 31033 22593 31067 22627
rect 31125 22593 31159 22627
rect 32413 22593 32447 22627
rect 33057 22593 33091 22627
rect 34069 22593 34103 22627
rect 34336 22593 34370 22627
rect 38485 22593 38519 22627
rect 38577 22593 38611 22627
rect 46857 22593 46891 22627
rect 47041 22593 47075 22627
rect 48881 22593 48915 22627
rect 26985 22525 27019 22559
rect 30941 22525 30975 22559
rect 31217 22525 31251 22559
rect 33333 22525 33367 22559
rect 37841 22525 37875 22559
rect 44097 22525 44131 22559
rect 44373 22525 44407 22559
rect 46673 22525 46707 22559
rect 47593 22525 47627 22559
rect 33241 22457 33275 22491
rect 38669 22457 38703 22491
rect 45845 22457 45879 22491
rect 68477 22457 68511 22491
rect 30113 22389 30147 22423
rect 30757 22389 30791 22423
rect 31677 22389 31711 22423
rect 31861 22389 31895 22423
rect 33149 22389 33183 22423
rect 38761 22389 38795 22423
rect 46857 22389 46891 22423
rect 48237 22389 48271 22423
rect 49433 22389 49467 22423
rect 28917 22185 28951 22219
rect 29193 22185 29227 22219
rect 31585 22185 31619 22219
rect 37473 22185 37507 22219
rect 44649 22185 44683 22219
rect 47317 22185 47351 22219
rect 47869 22185 47903 22219
rect 48605 22185 48639 22219
rect 29837 22117 29871 22151
rect 46397 22117 46431 22151
rect 48789 22117 48823 22151
rect 29561 22049 29595 22083
rect 35081 22049 35115 22083
rect 35909 22049 35943 22083
rect 37841 22049 37875 22083
rect 48881 22049 48915 22083
rect 27353 21981 27387 22015
rect 28733 21981 28767 22015
rect 30205 21981 30239 22015
rect 30472 21981 30506 22015
rect 35265 21981 35299 22015
rect 35449 21981 35483 22015
rect 35725 21981 35759 22015
rect 37749 21981 37783 22015
rect 38108 21981 38142 22015
rect 44833 21981 44867 22015
rect 45753 21981 45787 22015
rect 46489 21981 46523 22015
rect 46673 21981 46707 22015
rect 46765 21981 46799 22015
rect 46857 21981 46891 22015
rect 47501 21981 47535 22015
rect 47685 21981 47719 22015
rect 47777 21981 47811 22015
rect 48053 21981 48087 22015
rect 48237 21981 48271 22015
rect 48329 21981 48363 22015
rect 49065 21981 49099 22015
rect 49617 21981 49651 22015
rect 36154 21913 36188 21947
rect 37473 21913 37507 21947
rect 48421 21913 48455 21947
rect 27905 21845 27939 21879
rect 30021 21845 30055 21879
rect 35541 21845 35575 21879
rect 37289 21845 37323 21879
rect 37657 21845 37691 21879
rect 39221 21845 39255 21879
rect 47041 21845 47075 21879
rect 48621 21845 48655 21879
rect 49249 21845 49283 21879
rect 49709 21845 49743 21879
rect 29101 21641 29135 21675
rect 30865 21641 30899 21675
rect 31033 21641 31067 21675
rect 35541 21641 35575 21675
rect 35909 21641 35943 21675
rect 38485 21641 38519 21675
rect 46121 21641 46155 21675
rect 47041 21641 47075 21675
rect 47869 21641 47903 21675
rect 30665 21573 30699 21607
rect 36369 21573 36403 21607
rect 38577 21573 38611 21607
rect 38777 21573 38811 21607
rect 43913 21573 43947 21607
rect 46489 21573 46523 21607
rect 46581 21573 46615 21607
rect 1501 21505 1535 21539
rect 25688 21505 25722 21539
rect 26985 21505 27019 21539
rect 27169 21505 27203 21539
rect 27445 21505 27479 21539
rect 27629 21505 27663 21539
rect 27988 21505 28022 21539
rect 29469 21505 29503 21539
rect 32321 21505 32355 21539
rect 32588 21505 32622 21539
rect 34529 21505 34563 21539
rect 36553 21505 36587 21539
rect 36645 21505 36679 21539
rect 36737 21505 36771 21539
rect 36875 21505 36909 21539
rect 37933 21505 37967 21539
rect 42441 21505 42475 21539
rect 43637 21505 43671 21539
rect 46397 21505 46431 21539
rect 46699 21505 46733 21539
rect 46857 21505 46891 21539
rect 46949 21505 46983 21539
rect 47133 21505 47167 21539
rect 47225 21505 47259 21539
rect 47409 21505 47443 21539
rect 47777 21505 47811 21539
rect 48789 21505 48823 21539
rect 51549 21505 51583 21539
rect 25421 21437 25455 21471
rect 27721 21437 27755 21471
rect 33793 21437 33827 21471
rect 36001 21437 36035 21471
rect 36185 21437 36219 21471
rect 37013 21437 37047 21471
rect 45385 21437 45419 21471
rect 45569 21437 45603 21471
rect 46213 21437 46247 21471
rect 47317 21437 47351 21471
rect 49065 21437 49099 21471
rect 49341 21437 49375 21471
rect 50905 21437 50939 21471
rect 33701 21369 33735 21403
rect 1777 21301 1811 21335
rect 26801 21301 26835 21335
rect 30113 21301 30147 21335
rect 30849 21301 30883 21335
rect 34437 21301 34471 21335
rect 35173 21301 35207 21335
rect 38761 21301 38795 21335
rect 38945 21301 38979 21335
rect 42533 21301 42567 21335
rect 48881 21301 48915 21335
rect 50813 21301 50847 21335
rect 26617 21097 26651 21131
rect 29561 21097 29595 21131
rect 33425 21097 33459 21131
rect 36921 21097 36955 21131
rect 44557 21097 44591 21131
rect 46213 21097 46247 21131
rect 46397 21097 46431 21131
rect 47225 21097 47259 21131
rect 47409 21097 47443 21131
rect 47685 21097 47719 21131
rect 49157 21097 49191 21131
rect 49249 21097 49283 21131
rect 38577 21029 38611 21063
rect 38761 21029 38795 21063
rect 39589 21029 39623 21063
rect 25513 20961 25547 20995
rect 25697 20961 25731 20995
rect 33517 20961 33551 20995
rect 34713 20961 34747 20995
rect 39865 20961 39899 20995
rect 47593 20961 47627 20995
rect 49893 20961 49927 20995
rect 25421 20893 25455 20927
rect 25605 20893 25639 20927
rect 26801 20893 26835 20927
rect 26893 20893 26927 20927
rect 27077 20893 27111 20927
rect 27169 20893 27203 20927
rect 29745 20893 29779 20927
rect 29837 20893 29871 20927
rect 30021 20893 30055 20927
rect 30113 20893 30147 20927
rect 31677 20893 31711 20927
rect 33609 20893 33643 20927
rect 33885 20893 33919 20927
rect 33977 20893 34011 20927
rect 34969 20893 35003 20927
rect 36829 20893 36863 20927
rect 37013 20893 37047 20927
rect 38301 20893 38335 20927
rect 39037 20893 39071 20927
rect 39405 20893 39439 20927
rect 39681 20893 39715 20927
rect 41337 20893 41371 20927
rect 42809 20893 42843 20927
rect 43453 20893 43487 20927
rect 43729 20893 43763 20927
rect 43821 20893 43855 20927
rect 44005 20893 44039 20927
rect 44097 20893 44131 20927
rect 44465 20893 44499 20927
rect 46029 20893 46063 20927
rect 46673 20893 46707 20927
rect 46765 20893 46799 20927
rect 47501 20893 47535 20927
rect 49433 20893 49467 20927
rect 49525 20893 49559 20927
rect 49617 20893 49651 20927
rect 50353 20893 50387 20927
rect 50445 20893 50479 20927
rect 50537 20893 50571 20927
rect 50629 20893 50663 20927
rect 31944 20825 31978 20859
rect 38025 20825 38059 20859
rect 38209 20825 38243 20859
rect 38761 20825 38795 20859
rect 39221 20825 39255 20859
rect 40110 20825 40144 20859
rect 41604 20825 41638 20859
rect 43545 20825 43579 20859
rect 45845 20825 45879 20859
rect 46305 20825 46339 20859
rect 47041 20825 47075 20859
rect 48605 20825 48639 20859
rect 49755 20825 49789 20859
rect 26341 20757 26375 20791
rect 33057 20757 33091 20791
rect 33149 20757 33183 20791
rect 33793 20757 33827 20791
rect 34069 20757 34103 20791
rect 36093 20757 36127 20791
rect 38393 20757 38427 20791
rect 38945 20757 38979 20791
rect 41245 20757 41279 20791
rect 42717 20757 42751 20791
rect 46949 20757 46983 20791
rect 47251 20757 47285 20791
rect 47869 20757 47903 20791
rect 48789 20757 48823 20791
rect 48881 20757 48915 20791
rect 48973 20757 49007 20791
rect 50169 20757 50203 20791
rect 26801 20553 26835 20587
rect 28089 20553 28123 20587
rect 28273 20553 28307 20587
rect 32781 20553 32815 20587
rect 33073 20553 33107 20587
rect 33977 20553 34011 20587
rect 39497 20553 39531 20587
rect 40233 20553 40267 20587
rect 40509 20553 40543 20587
rect 40969 20553 41003 20587
rect 41153 20553 41187 20587
rect 45293 20553 45327 20587
rect 47409 20553 47443 20587
rect 48329 20553 48363 20587
rect 25228 20485 25262 20519
rect 32873 20485 32907 20519
rect 34805 20485 34839 20519
rect 37657 20485 37691 20519
rect 37873 20485 37907 20519
rect 50261 20485 50295 20519
rect 24961 20417 24995 20451
rect 26617 20417 26651 20451
rect 28549 20417 28583 20451
rect 28733 20417 28767 20451
rect 28825 20417 28859 20451
rect 29092 20417 29126 20451
rect 30564 20417 30598 20451
rect 32229 20417 32263 20451
rect 33333 20417 33367 20451
rect 34069 20417 34103 20451
rect 35173 20417 35207 20451
rect 36277 20417 36311 20451
rect 36461 20417 36495 20451
rect 38209 20417 38243 20451
rect 39681 20417 39715 20451
rect 40325 20417 40359 20451
rect 40601 20417 40635 20451
rect 40693 20417 40727 20451
rect 40877 20417 40911 20451
rect 41150 20417 41184 20451
rect 42533 20417 42567 20451
rect 45109 20417 45143 20451
rect 46765 20417 46799 20451
rect 47133 20417 47167 20451
rect 47225 20417 47259 20451
rect 48053 20417 48087 20451
rect 48421 20417 48455 20451
rect 48697 20417 48731 20451
rect 50077 20417 50111 20451
rect 50353 20439 50387 20473
rect 26433 20349 26467 20383
rect 27077 20349 27111 20383
rect 30297 20349 30331 20383
rect 38853 20349 38887 20383
rect 41613 20349 41647 20383
rect 42809 20349 42843 20383
rect 44373 20349 44407 20383
rect 48789 20349 48823 20383
rect 26341 20281 26375 20315
rect 27721 20281 27755 20315
rect 35725 20281 35759 20315
rect 38761 20281 38795 20315
rect 40325 20281 40359 20315
rect 47685 20281 47719 20315
rect 48145 20281 48179 20315
rect 49065 20281 49099 20315
rect 27629 20213 27663 20247
rect 28089 20213 28123 20247
rect 28641 20213 28675 20247
rect 30205 20213 30239 20247
rect 31677 20213 31711 20247
rect 33057 20213 33091 20247
rect 33241 20213 33275 20247
rect 36369 20213 36403 20247
rect 37841 20213 37875 20247
rect 38025 20213 38059 20247
rect 40693 20213 40727 20247
rect 41521 20213 41555 20247
rect 44281 20213 44315 20247
rect 45017 20213 45051 20247
rect 46949 20213 46983 20247
rect 47961 20213 47995 20247
rect 50169 20213 50203 20247
rect 26525 20009 26559 20043
rect 29745 20009 29779 20043
rect 30665 20009 30699 20043
rect 32045 20009 32079 20043
rect 32597 20009 32631 20043
rect 32965 20009 32999 20043
rect 41429 20009 41463 20043
rect 42441 20009 42475 20043
rect 43545 20009 43579 20043
rect 31033 19941 31067 19975
rect 33425 19941 33459 19975
rect 33701 19941 33735 19975
rect 34253 19941 34287 19975
rect 38853 19941 38887 19975
rect 44741 19941 44775 19975
rect 46765 19941 46799 19975
rect 48237 19941 48271 19975
rect 26617 19873 26651 19907
rect 27353 19873 27387 19907
rect 27905 19873 27939 19907
rect 29193 19873 29227 19907
rect 31125 19873 31159 19907
rect 31493 19873 31527 19907
rect 33241 19873 33275 19907
rect 33793 19873 33827 19907
rect 35633 19873 35667 19907
rect 37473 19873 37507 19907
rect 39865 19873 39899 19907
rect 46489 19873 46523 19907
rect 46857 19873 46891 19907
rect 47593 19873 47627 19907
rect 47869 19873 47903 19907
rect 49341 19873 49375 19907
rect 50445 19873 50479 19907
rect 52193 19873 52227 19907
rect 26341 19805 26375 19839
rect 26433 19805 26467 19839
rect 27169 19805 27203 19839
rect 27261 19805 27295 19839
rect 27445 19805 27479 19839
rect 28089 19805 28123 19839
rect 30849 19805 30883 19839
rect 32321 19805 32355 19839
rect 32781 19805 32815 19839
rect 32873 19805 32907 19839
rect 33149 19805 33183 19839
rect 33333 19805 33367 19839
rect 33609 19805 33643 19839
rect 33885 19805 33919 19839
rect 34253 19805 34287 19839
rect 34437 19805 34471 19839
rect 34989 19805 35023 19839
rect 37105 19805 37139 19839
rect 37197 19805 37231 19839
rect 39221 19805 39255 19839
rect 40132 19805 40166 19839
rect 41337 19805 41371 19839
rect 42625 19805 42659 19839
rect 43453 19805 43487 19839
rect 44557 19805 44591 19839
rect 44833 19805 44867 19839
rect 45017 19805 45051 19839
rect 46673 19805 46707 19839
rect 46949 19805 46983 19839
rect 47133 19805 47167 19839
rect 47501 19805 47535 19839
rect 47685 19805 47719 19839
rect 49525 19805 49559 19839
rect 49617 19805 49651 19839
rect 49985 19805 50019 19839
rect 50169 19805 50203 19839
rect 68477 19805 68511 19839
rect 28457 19737 28491 19771
rect 29561 19737 29595 19771
rect 35900 19737 35934 19771
rect 37381 19737 37415 19771
rect 37718 19737 37752 19771
rect 39405 19737 39439 19771
rect 44373 19737 44407 19771
rect 45262 19737 45296 19771
rect 49709 19737 49743 19771
rect 49847 19737 49881 19771
rect 26985 19669 27019 19703
rect 28273 19669 28307 19703
rect 29761 19669 29795 19703
rect 29929 19669 29963 19703
rect 32413 19669 32447 19703
rect 34805 19669 34839 19703
rect 37013 19669 37047 19703
rect 37105 19669 37139 19703
rect 41245 19669 41279 19703
rect 46397 19669 46431 19703
rect 48329 19669 48363 19703
rect 27629 19465 27663 19499
rect 29009 19465 29043 19499
rect 33793 19465 33827 19499
rect 35633 19465 35667 19499
rect 36645 19465 36679 19499
rect 42993 19465 43027 19499
rect 46029 19465 46063 19499
rect 46765 19465 46799 19499
rect 50169 19465 50203 19499
rect 31861 19397 31895 19431
rect 33977 19397 34011 19431
rect 34520 19397 34554 19431
rect 42073 19397 42107 19431
rect 42717 19397 42751 19431
rect 43913 19397 43947 19431
rect 47593 19397 47627 19431
rect 50537 19397 50571 19431
rect 26157 19329 26191 19363
rect 26985 19329 27019 19363
rect 27261 19329 27295 19363
rect 27445 19329 27479 19363
rect 27905 19329 27939 19363
rect 27997 19329 28031 19363
rect 28089 19329 28123 19363
rect 28549 19329 28583 19363
rect 28733 19329 28767 19363
rect 29193 19329 29227 19363
rect 31585 19329 31619 19363
rect 32137 19329 32171 19363
rect 32393 19329 32427 19363
rect 33885 19329 33919 19363
rect 34253 19329 34287 19363
rect 39681 19329 39715 19363
rect 41337 19329 41371 19363
rect 42441 19329 42475 19363
rect 43361 19329 43395 19363
rect 43821 19329 43855 19363
rect 44005 19329 44039 19363
rect 46305 19329 46339 19363
rect 46949 19329 46983 19363
rect 47041 19329 47075 19363
rect 47317 19329 47351 19363
rect 47777 19329 47811 19363
rect 50353 19329 50387 19363
rect 50629 19329 50663 19363
rect 28825 19261 28859 19295
rect 36093 19261 36127 19295
rect 37289 19261 37323 19295
rect 42533 19261 42567 19295
rect 43453 19261 43487 19295
rect 43545 19261 43579 19295
rect 45477 19261 45511 19295
rect 46121 19261 46155 19295
rect 27721 19193 27755 19227
rect 31585 19193 31619 19227
rect 31677 19193 31711 19227
rect 33517 19193 33551 19227
rect 33609 19193 33643 19227
rect 46489 19193 46523 19227
rect 26249 19125 26283 19159
rect 27445 19125 27479 19159
rect 28273 19125 28307 19159
rect 28365 19125 28399 19159
rect 34161 19125 34195 19159
rect 37933 19125 37967 19159
rect 39773 19125 39807 19159
rect 42625 19125 42659 19159
rect 47225 19125 47259 19159
rect 47961 19125 47995 19159
rect 27445 18921 27479 18955
rect 27629 18921 27663 18955
rect 31677 18921 31711 18955
rect 32873 18921 32907 18955
rect 34161 18921 34195 18955
rect 34345 18921 34379 18955
rect 36645 18921 36679 18955
rect 36829 18921 36863 18955
rect 43269 18921 43303 18955
rect 45937 18921 45971 18955
rect 46121 18921 46155 18955
rect 47409 18921 47443 18955
rect 51089 18921 51123 18955
rect 42165 18853 42199 18887
rect 33333 18785 33367 18819
rect 42625 18785 42659 18819
rect 43821 18785 43855 18819
rect 44281 18785 44315 18819
rect 45017 18785 45051 18819
rect 46857 18785 46891 18819
rect 50629 18785 50663 18819
rect 50813 18785 50847 18819
rect 1593 18717 1627 18751
rect 25605 18717 25639 18751
rect 25872 18717 25906 18751
rect 27077 18717 27111 18751
rect 29561 18717 29595 18751
rect 33149 18717 33183 18751
rect 34713 18717 34747 18751
rect 36001 18717 36035 18751
rect 36149 18717 36183 18751
rect 36277 18717 36311 18751
rect 36369 18717 36403 18751
rect 36507 18717 36541 18751
rect 37089 18727 37123 18761
rect 37197 18717 37231 18751
rect 37933 18717 37967 18751
rect 38081 18717 38115 18751
rect 38398 18717 38432 18751
rect 38945 18717 38979 18751
rect 40141 18717 40175 18751
rect 40785 18717 40819 18751
rect 43269 18717 43303 18751
rect 43545 18717 43579 18751
rect 43729 18717 43763 18751
rect 43913 18717 43947 18751
rect 44189 18717 44223 18751
rect 44373 18717 44407 18751
rect 44649 18717 44683 18751
rect 46305 18717 46339 18751
rect 47041 18717 47075 18751
rect 47225 18717 47259 18751
rect 47317 18717 47351 18751
rect 48697 18717 48731 18751
rect 48881 18717 48915 18751
rect 48973 18717 49007 18751
rect 50537 18717 50571 18751
rect 50997 18717 51031 18751
rect 28457 18649 28491 18683
rect 29193 18649 29227 18683
rect 29828 18649 29862 18683
rect 31401 18649 31435 18683
rect 32873 18649 32907 18683
rect 33885 18649 33919 18683
rect 33977 18649 34011 18683
rect 35449 18649 35483 18683
rect 36829 18649 36863 18683
rect 38209 18649 38243 18683
rect 38301 18649 38335 18683
rect 41052 18649 41086 18683
rect 45753 18649 45787 18683
rect 45953 18649 45987 18683
rect 47685 18649 47719 18683
rect 48421 18649 48455 18683
rect 26985 18581 27019 18615
rect 27445 18581 27479 18615
rect 30941 18581 30975 18615
rect 33057 18581 33091 18615
rect 34177 18581 34211 18615
rect 37013 18581 37047 18615
rect 37841 18581 37875 18615
rect 38577 18581 38611 18615
rect 39497 18581 39531 18615
rect 40693 18581 40727 18615
rect 43177 18581 43211 18615
rect 43453 18581 43487 18615
rect 44741 18581 44775 18615
rect 45661 18581 45695 18615
rect 46489 18581 46523 18615
rect 48789 18581 48823 18615
rect 49065 18581 49099 18615
rect 50169 18581 50203 18615
rect 30113 18377 30147 18411
rect 33425 18377 33459 18411
rect 33517 18377 33551 18411
rect 33701 18377 33735 18411
rect 34003 18377 34037 18411
rect 38393 18377 38427 18411
rect 40233 18377 40267 18411
rect 41153 18377 41187 18411
rect 44925 18377 44959 18411
rect 45017 18377 45051 18411
rect 46581 18377 46615 18411
rect 29193 18309 29227 18343
rect 29653 18309 29687 18343
rect 30021 18309 30055 18343
rect 31309 18309 31343 18343
rect 33149 18309 33183 18343
rect 33793 18309 33827 18343
rect 37381 18309 37415 18343
rect 37597 18309 37631 18343
rect 42073 18309 42107 18343
rect 47134 18309 47168 18343
rect 47251 18309 47285 18343
rect 51733 18309 51767 18343
rect 27629 18241 27663 18275
rect 29469 18241 29503 18275
rect 30665 18241 30699 18275
rect 31493 18241 31527 18275
rect 31585 18241 31619 18275
rect 32873 18241 32907 18275
rect 33333 18241 33367 18275
rect 35265 18241 35299 18275
rect 35532 18241 35566 18275
rect 36829 18241 36863 18275
rect 37841 18241 37875 18275
rect 38117 18241 38151 18275
rect 38669 18241 38703 18275
rect 38853 18241 38887 18275
rect 39109 18241 39143 18275
rect 41061 18241 41095 18275
rect 41245 18241 41279 18275
rect 41337 18241 41371 18275
rect 42441 18241 42475 18275
rect 42697 18241 42731 18275
rect 44373 18241 44407 18275
rect 45293 18241 45327 18275
rect 45385 18241 45419 18275
rect 45477 18241 45511 18275
rect 45661 18241 45695 18275
rect 46489 18241 46523 18275
rect 46673 18241 46707 18275
rect 46949 18241 46983 18275
rect 47041 18241 47075 18275
rect 47593 18241 47627 18275
rect 49709 18241 49743 18275
rect 32137 18173 32171 18207
rect 33701 18173 33735 18207
rect 36921 18173 36955 18207
rect 37105 18173 37139 18207
rect 45753 18173 45787 18207
rect 47409 18173 47443 18207
rect 47869 18173 47903 18207
rect 49617 18173 49651 18207
rect 49985 18173 50019 18207
rect 28825 18105 28859 18139
rect 29837 18105 29871 18139
rect 30481 18105 30515 18139
rect 32965 18105 32999 18139
rect 34161 18105 34195 18139
rect 36645 18105 36679 18139
rect 43821 18105 43855 18139
rect 28273 18037 28307 18071
rect 29193 18037 29227 18071
rect 29377 18037 29411 18071
rect 31309 18037 31343 18071
rect 32781 18037 32815 18071
rect 32873 18037 32907 18071
rect 33977 18037 34011 18071
rect 37013 18037 37047 18071
rect 37565 18037 37599 18071
rect 37749 18037 37783 18071
rect 46397 18037 46431 18071
rect 46765 18037 46799 18071
rect 27445 17833 27479 17867
rect 30573 17833 30607 17867
rect 32137 17833 32171 17867
rect 32229 17833 32263 17867
rect 34437 17833 34471 17867
rect 35817 17833 35851 17867
rect 38577 17833 38611 17867
rect 39313 17833 39347 17867
rect 43361 17833 43395 17867
rect 46489 17833 46523 17867
rect 47317 17833 47351 17867
rect 49249 17833 49283 17867
rect 50629 17833 50663 17867
rect 28089 17765 28123 17799
rect 44189 17765 44223 17799
rect 44281 17765 44315 17799
rect 27813 17697 27847 17731
rect 32689 17697 32723 17731
rect 34529 17697 34563 17731
rect 35357 17697 35391 17731
rect 38669 17697 38703 17731
rect 48145 17697 48179 17731
rect 49065 17697 49099 17731
rect 26065 17629 26099 17663
rect 27721 17629 27755 17663
rect 28181 17629 28215 17663
rect 28365 17629 28399 17663
rect 30297 17629 30331 17663
rect 30757 17629 30791 17663
rect 31024 17629 31058 17663
rect 32413 17629 32447 17663
rect 32505 17629 32539 17663
rect 33425 17629 33459 17663
rect 34069 17629 34103 17663
rect 34253 17629 34287 17663
rect 34713 17629 34747 17663
rect 36001 17629 36035 17663
rect 36277 17629 36311 17663
rect 36461 17629 36495 17663
rect 36737 17629 36771 17663
rect 36829 17629 36863 17663
rect 37013 17629 37047 17663
rect 37105 17629 37139 17663
rect 37197 17629 37231 17663
rect 37453 17629 37487 17663
rect 39405 17629 39439 17663
rect 39589 17629 39623 17663
rect 43545 17629 43579 17663
rect 43821 17629 43855 17663
rect 44097 17629 44131 17663
rect 44373 17629 44407 17663
rect 45109 17629 45143 17663
rect 46673 17629 46707 17663
rect 47409 17629 47443 17663
rect 49433 17629 49467 17663
rect 50537 17629 50571 17663
rect 26332 17561 26366 17595
rect 28273 17561 28307 17595
rect 29009 17561 29043 17595
rect 29745 17561 29779 17595
rect 30113 17561 30147 17595
rect 32229 17561 32263 17595
rect 36553 17561 36587 17595
rect 43729 17561 43763 17595
rect 45376 17561 45410 17595
rect 29101 17493 29135 17527
rect 33241 17493 33275 17527
rect 33977 17493 34011 17527
rect 39497 17493 39531 17527
rect 43913 17493 43947 17527
rect 48421 17493 48455 17527
rect 48789 17493 48823 17527
rect 48881 17493 48915 17527
rect 29377 17289 29411 17323
rect 31861 17289 31895 17323
rect 33609 17289 33643 17323
rect 35081 17289 35115 17323
rect 36277 17289 36311 17323
rect 41613 17289 41647 17323
rect 44189 17289 44223 17323
rect 46857 17289 46891 17323
rect 36093 17221 36127 17255
rect 50169 17221 50203 17255
rect 26157 17153 26191 17187
rect 28172 17153 28206 17187
rect 29561 17153 29595 17187
rect 30481 17153 30515 17187
rect 31585 17153 31619 17187
rect 31677 17153 31711 17187
rect 32229 17153 32263 17187
rect 32496 17153 32530 17187
rect 33701 17153 33735 17187
rect 33968 17153 34002 17187
rect 35725 17153 35759 17187
rect 35909 17153 35943 17187
rect 36369 17153 36403 17187
rect 38853 17153 38887 17187
rect 39129 17153 39163 17187
rect 39313 17153 39347 17187
rect 39497 17153 39531 17187
rect 39753 17153 39787 17187
rect 43076 17153 43110 17187
rect 46397 17153 46431 17187
rect 46765 17153 46799 17187
rect 50077 17153 50111 17187
rect 27905 17085 27939 17119
rect 31861 17085 31895 17119
rect 38669 17085 38703 17119
rect 40969 17085 41003 17119
rect 42809 17085 42843 17119
rect 44373 17085 44407 17119
rect 46673 17085 46707 17119
rect 48237 17085 48271 17119
rect 48513 17085 48547 17119
rect 36093 17017 36127 17051
rect 46581 17017 46615 17051
rect 68477 17017 68511 17051
rect 25973 16949 26007 16983
rect 29285 16949 29319 16983
rect 30297 16949 30331 16983
rect 35725 16949 35759 16983
rect 40877 16949 40911 16983
rect 44925 16949 44959 16983
rect 46213 16949 46247 16983
rect 49985 16949 50019 16983
rect 28181 16745 28215 16779
rect 37841 16745 37875 16779
rect 39497 16745 39531 16779
rect 44833 16745 44867 16779
rect 48237 16745 48271 16779
rect 49157 16745 49191 16779
rect 36737 16677 36771 16711
rect 39681 16677 39715 16711
rect 39865 16677 39899 16711
rect 41521 16677 41555 16711
rect 44189 16677 44223 16711
rect 45017 16677 45051 16711
rect 48145 16677 48179 16711
rect 27537 16609 27571 16643
rect 28457 16609 28491 16643
rect 29745 16609 29779 16643
rect 37197 16609 37231 16643
rect 38669 16609 38703 16643
rect 39129 16609 39163 16643
rect 41613 16609 41647 16643
rect 42809 16609 42843 16643
rect 43637 16609 43671 16643
rect 46121 16609 46155 16643
rect 48513 16609 48547 16643
rect 49249 16609 49283 16643
rect 25513 16541 25547 16575
rect 25780 16541 25814 16575
rect 27813 16541 27847 16575
rect 27997 16541 28031 16575
rect 29285 16541 29319 16575
rect 29377 16541 29411 16575
rect 30012 16541 30046 16575
rect 35357 16541 35391 16575
rect 35624 16541 35658 16575
rect 38117 16541 38151 16575
rect 38853 16541 38887 16575
rect 40049 16541 40083 16575
rect 40141 16541 40175 16575
rect 42441 16541 42475 16575
rect 42717 16541 42751 16575
rect 44281 16541 44315 16575
rect 44649 16541 44683 16575
rect 45293 16541 45327 16575
rect 45385 16541 45419 16575
rect 45569 16541 45603 16575
rect 46765 16541 46799 16575
rect 48421 16541 48455 16575
rect 51273 16541 51307 16575
rect 51825 16541 51859 16575
rect 27445 16473 27479 16507
rect 29009 16473 29043 16507
rect 29101 16473 29135 16507
rect 38209 16473 38243 16507
rect 40386 16473 40420 16507
rect 44465 16473 44499 16507
rect 44557 16473 44591 16507
rect 45017 16473 45051 16507
rect 45477 16473 45511 16507
rect 46673 16473 46707 16507
rect 47010 16473 47044 16507
rect 26893 16405 26927 16439
rect 26985 16405 27019 16439
rect 27353 16405 27387 16439
rect 29199 16405 29233 16439
rect 31125 16405 31159 16439
rect 39037 16405 39071 16439
rect 39497 16405 39531 16439
rect 42257 16405 42291 16439
rect 42539 16405 42573 16439
rect 42625 16405 42659 16439
rect 43453 16405 43487 16439
rect 45201 16405 45235 16439
rect 49893 16405 49927 16439
rect 51365 16405 51399 16439
rect 52377 16405 52411 16439
rect 26617 16201 26651 16235
rect 29193 16201 29227 16235
rect 32505 16201 32539 16235
rect 40877 16201 40911 16235
rect 44005 16201 44039 16235
rect 51917 16201 51951 16235
rect 25973 16133 26007 16167
rect 30849 16133 30883 16167
rect 37565 16133 37599 16167
rect 40693 16133 40727 16167
rect 44741 16133 44775 16167
rect 25789 16065 25823 16099
rect 26065 16065 26099 16099
rect 26433 16065 26467 16099
rect 27804 16065 27838 16099
rect 29101 16065 29135 16099
rect 29285 16065 29319 16099
rect 29469 16065 29503 16099
rect 30573 16065 30607 16099
rect 30757 16065 30791 16099
rect 30941 16065 30975 16099
rect 32321 16065 32355 16099
rect 33333 16065 33367 16099
rect 33425 16065 33459 16099
rect 33609 16065 33643 16099
rect 33701 16065 33735 16099
rect 34437 16065 34471 16099
rect 39129 16065 39163 16099
rect 39396 16065 39430 16099
rect 40969 16065 41003 16099
rect 42441 16065 42475 16099
rect 42708 16065 42742 16099
rect 43913 16065 43947 16099
rect 44097 16065 44131 16099
rect 46489 16065 46523 16099
rect 47041 16065 47075 16099
rect 47225 16065 47259 16099
rect 26249 15997 26283 16031
rect 27537 15997 27571 16031
rect 31217 15997 31251 16031
rect 32137 15997 32171 16031
rect 33793 15997 33827 16031
rect 37289 15997 37323 16031
rect 44465 15997 44499 16031
rect 46765 15997 46799 16031
rect 50169 15997 50203 16031
rect 50445 15997 50479 16031
rect 30113 15929 30147 15963
rect 31125 15929 31159 15963
rect 40693 15929 40727 15963
rect 1593 15861 1627 15895
rect 25789 15861 25823 15895
rect 28917 15861 28951 15895
rect 31861 15861 31895 15895
rect 33149 15861 33183 15895
rect 39037 15861 39071 15895
rect 40509 15861 40543 15895
rect 43821 15861 43855 15895
rect 46213 15861 46247 15895
rect 46305 15861 46339 15895
rect 46673 15861 46707 15895
rect 47041 15861 47075 15895
rect 27445 15657 27479 15691
rect 29837 15657 29871 15691
rect 32137 15657 32171 15691
rect 38117 15657 38151 15691
rect 39313 15657 39347 15691
rect 42901 15657 42935 15691
rect 45753 15657 45787 15691
rect 51365 15657 51399 15691
rect 27537 15589 27571 15623
rect 42073 15589 42107 15623
rect 28641 15521 28675 15555
rect 40693 15521 40727 15555
rect 42257 15521 42291 15555
rect 42993 15521 43027 15555
rect 43361 15521 43395 15555
rect 44787 15521 44821 15555
rect 45109 15521 45143 15555
rect 46121 15521 46155 15555
rect 46765 15521 46799 15555
rect 52101 15521 52135 15555
rect 25145 15453 25179 15487
rect 26065 15453 26099 15487
rect 26801 15453 26835 15487
rect 27445 15453 27479 15487
rect 27905 15453 27939 15487
rect 29745 15453 29779 15487
rect 29837 15453 29871 15487
rect 30021 15453 30055 15487
rect 30757 15453 30791 15487
rect 32597 15453 32631 15487
rect 34713 15453 34747 15487
rect 37473 15453 37507 15487
rect 38025 15453 38059 15487
rect 38853 15453 38887 15487
rect 39497 15453 39531 15487
rect 40325 15453 40359 15487
rect 40417 15453 40451 15487
rect 40509 15453 40543 15487
rect 48237 15453 48271 15487
rect 49801 15453 49835 15487
rect 50813 15453 50847 15487
rect 51457 15453 51491 15487
rect 51650 15463 51684 15497
rect 51825 15453 51859 15487
rect 51963 15453 51997 15487
rect 52561 15453 52595 15487
rect 52653 15453 52687 15487
rect 52837 15453 52871 15487
rect 53389 15453 53423 15487
rect 27721 15385 27755 15419
rect 29193 15385 29227 15419
rect 31024 15385 31058 15419
rect 32864 15385 32898 15419
rect 34958 15385 34992 15419
rect 37749 15385 37783 15419
rect 39221 15385 39255 15419
rect 40141 15385 40175 15419
rect 40938 15385 40972 15419
rect 46673 15385 46707 15419
rect 47010 15385 47044 15419
rect 51734 15385 51768 15419
rect 52193 15385 52227 15419
rect 52377 15385 52411 15419
rect 52745 15385 52779 15419
rect 25697 15317 25731 15351
rect 26617 15317 26651 15351
rect 27353 15317 27387 15351
rect 28457 15317 28491 15351
rect 29561 15317 29595 15351
rect 33977 15317 34011 15351
rect 36093 15317 36127 15351
rect 48145 15317 48179 15351
rect 48329 15317 48363 15351
rect 49893 15317 49927 15351
rect 53941 15317 53975 15351
rect 26617 15113 26651 15147
rect 27077 15113 27111 15147
rect 28641 15113 28675 15147
rect 29101 15113 29135 15147
rect 30849 15113 30883 15147
rect 31677 15113 31711 15147
rect 33701 15113 33735 15147
rect 34437 15113 34471 15147
rect 42441 15113 42475 15147
rect 44557 15113 44591 15147
rect 45385 15113 45419 15147
rect 54493 15113 54527 15147
rect 25504 15045 25538 15079
rect 29714 15045 29748 15079
rect 38485 15045 38519 15079
rect 41245 15045 41279 15079
rect 51273 15045 51307 15079
rect 51503 15011 51537 15045
rect 23765 14977 23799 15011
rect 24032 14977 24066 15011
rect 26985 14977 27019 15011
rect 27169 14977 27203 15011
rect 27353 14977 27387 15011
rect 28089 14977 28123 15011
rect 28733 14977 28767 15011
rect 28917 14977 28951 15011
rect 29193 14977 29227 15011
rect 29469 14977 29503 15011
rect 31769 14977 31803 15011
rect 32588 14977 32622 15011
rect 34434 14977 34468 15011
rect 34897 14977 34931 15011
rect 34989 14977 35023 15011
rect 35364 14977 35398 15011
rect 35624 14977 35658 15011
rect 36829 14977 36863 15011
rect 37013 14977 37047 15011
rect 39497 14977 39531 15011
rect 39957 14977 39991 15011
rect 40233 14977 40267 15011
rect 40417 14977 40451 15011
rect 40509 14977 40543 15011
rect 40601 14977 40635 15011
rect 40969 14977 41003 15011
rect 42625 14977 42659 15011
rect 42717 14977 42751 15011
rect 42901 14977 42935 15011
rect 42993 14977 43027 15011
rect 44465 14977 44499 15011
rect 45017 14977 45051 15011
rect 45201 14977 45235 15011
rect 45937 14977 45971 15011
rect 46204 14977 46238 15011
rect 48421 14977 48455 15011
rect 48513 14977 48547 15011
rect 48881 14977 48915 15011
rect 51733 14977 51767 15011
rect 51917 14977 51951 15011
rect 52009 14977 52043 15011
rect 52101 14977 52135 15011
rect 52377 14977 52411 15011
rect 52561 14977 52595 15011
rect 52745 14977 52779 15011
rect 25237 14909 25271 14943
rect 31033 14909 31067 14943
rect 32321 14909 32355 14943
rect 34805 14909 34839 14943
rect 39773 14909 39807 14943
rect 43821 14909 43855 14943
rect 44373 14909 44407 14943
rect 47593 14909 47627 14943
rect 48697 14909 48731 14943
rect 49157 14909 49191 14943
rect 53021 14909 53055 14943
rect 47317 14841 47351 14875
rect 51641 14841 51675 14875
rect 52285 14841 52319 14875
rect 25145 14773 25179 14807
rect 27905 14773 27939 14807
rect 29285 14773 29319 14807
rect 31861 14773 31895 14807
rect 34253 14773 34287 14807
rect 35081 14773 35115 14807
rect 36737 14773 36771 14807
rect 36829 14773 36863 14807
rect 38761 14773 38795 14807
rect 39589 14773 39623 14807
rect 40141 14773 40175 14807
rect 40785 14773 40819 14807
rect 48237 14773 48271 14807
rect 50629 14773 50663 14807
rect 51457 14773 51491 14807
rect 52377 14773 52411 14807
rect 26341 14569 26375 14603
rect 26893 14569 26927 14603
rect 31033 14569 31067 14603
rect 33149 14569 33183 14603
rect 34529 14569 34563 14603
rect 34713 14569 34747 14603
rect 36461 14569 36495 14603
rect 42165 14569 42199 14603
rect 42901 14569 42935 14603
rect 46949 14569 46983 14603
rect 47777 14569 47811 14603
rect 49525 14569 49559 14603
rect 51089 14569 51123 14603
rect 52837 14569 52871 14603
rect 29929 14501 29963 14535
rect 42349 14501 42383 14535
rect 43729 14501 43763 14535
rect 47317 14501 47351 14535
rect 47409 14501 47443 14535
rect 49249 14501 49283 14535
rect 25973 14433 26007 14467
rect 27261 14433 27295 14467
rect 33977 14433 34011 14467
rect 36737 14433 36771 14467
rect 40601 14433 40635 14467
rect 25789 14365 25823 14399
rect 25881 14365 25915 14399
rect 26249 14365 26283 14399
rect 26893 14365 26927 14399
rect 27169 14365 27203 14399
rect 28825 14365 28859 14399
rect 29561 14365 29595 14399
rect 29745 14365 29779 14399
rect 29837 14365 29871 14399
rect 30021 14365 30055 14399
rect 30205 14365 30239 14399
rect 31217 14365 31251 14399
rect 31309 14365 31343 14399
rect 31493 14365 31527 14399
rect 31585 14365 31619 14399
rect 31953 14365 31987 14399
rect 32597 14365 32631 14399
rect 33333 14365 33367 14399
rect 34897 14365 34931 14399
rect 35199 14365 35233 14399
rect 35357 14365 35391 14399
rect 36185 14365 36219 14399
rect 36277 14365 36311 14399
rect 37289 14365 37323 14399
rect 39865 14365 39899 14399
rect 41613 14365 41647 14399
rect 42530 14365 42564 14399
rect 42993 14365 43027 14399
rect 43085 14365 43119 14399
rect 43269 14365 43303 14399
rect 43637 14365 43671 14399
rect 46397 14365 46431 14399
rect 47041 14365 47075 14399
rect 47225 14365 47259 14399
rect 47501 14365 47535 14399
rect 47685 14365 47719 14399
rect 48145 14365 48179 14399
rect 48329 14365 48363 14399
rect 48421 14365 48455 14399
rect 48605 14365 48639 14399
rect 49065 14365 49099 14399
rect 49709 14365 49743 14399
rect 50997 14365 51031 14399
rect 51089 14365 51123 14399
rect 51549 14365 51583 14399
rect 51733 14365 51767 14399
rect 52745 14365 52779 14399
rect 68477 14365 68511 14399
rect 27528 14297 27562 14331
rect 29377 14297 29411 14331
rect 32873 14297 32907 14331
rect 34989 14297 35023 14331
rect 35081 14297 35115 14331
rect 37473 14297 37507 14331
rect 50629 14297 50663 14331
rect 25421 14229 25455 14263
rect 27077 14229 27111 14263
rect 28641 14229 28675 14263
rect 32505 14229 32539 14263
rect 35817 14229 35851 14263
rect 38761 14229 38795 14263
rect 40509 14229 40543 14263
rect 41245 14229 41279 14263
rect 42533 14229 42567 14263
rect 43177 14229 43211 14263
rect 48237 14229 48271 14263
rect 48605 14229 48639 14263
rect 51273 14229 51307 14263
rect 51641 14229 51675 14263
rect 33517 14025 33551 14059
rect 33609 14025 33643 14059
rect 34345 14025 34379 14059
rect 38669 14025 38703 14059
rect 40233 14025 40267 14059
rect 42257 14025 42291 14059
rect 44741 14025 44775 14059
rect 45569 14025 45603 14059
rect 50721 14025 50755 14059
rect 51917 14025 51951 14059
rect 52377 14025 52411 14059
rect 36553 13957 36587 13991
rect 37534 13957 37568 13991
rect 39120 13957 39154 13991
rect 42708 13957 42742 13991
rect 27813 13889 27847 13923
rect 27997 13889 28031 13923
rect 28089 13889 28123 13923
rect 29736 13889 29770 13923
rect 32137 13889 32171 13923
rect 32404 13889 32438 13923
rect 33793 13889 33827 13923
rect 33885 13889 33919 13923
rect 34069 13889 34103 13923
rect 34253 13889 34287 13923
rect 34437 13889 34471 13923
rect 36369 13889 36403 13923
rect 36645 13889 36679 13923
rect 36737 13889 36771 13923
rect 37289 13889 37323 13923
rect 41133 13889 41167 13923
rect 45661 13889 45695 13923
rect 46213 13889 46247 13923
rect 46489 13889 46523 13923
rect 46673 13889 46707 13923
rect 48053 13889 48087 13923
rect 48237 13889 48271 13923
rect 48329 13889 48363 13923
rect 48513 13889 48547 13923
rect 48789 13889 48823 13923
rect 49065 13889 49099 13923
rect 49249 13889 49283 13923
rect 49709 13889 49743 13923
rect 50077 13889 50111 13923
rect 50169 13889 50203 13923
rect 51089 13889 51123 13923
rect 51549 13889 51583 13923
rect 51733 13889 51767 13923
rect 52193 13889 52227 13923
rect 22937 13821 22971 13855
rect 23213 13821 23247 13855
rect 24961 13821 24995 13855
rect 28181 13821 28215 13855
rect 29469 13821 29503 13855
rect 31217 13821 31251 13855
rect 38853 13821 38887 13855
rect 40877 13821 40911 13855
rect 42441 13821 42475 13855
rect 44833 13821 44867 13855
rect 45017 13821 45051 13855
rect 45845 13821 45879 13855
rect 46029 13821 46063 13855
rect 48145 13821 48179 13855
rect 48605 13821 48639 13855
rect 48973 13821 49007 13855
rect 51181 13821 51215 13855
rect 51273 13821 51307 13855
rect 52009 13821 52043 13855
rect 30849 13753 30883 13787
rect 36921 13753 36955 13787
rect 43821 13753 43855 13787
rect 50353 13753 50387 13787
rect 27813 13685 27847 13719
rect 31769 13685 31803 13719
rect 33885 13685 33919 13719
rect 44373 13685 44407 13719
rect 45201 13685 45235 13719
rect 46397 13685 46431 13719
rect 46489 13685 46523 13719
rect 47869 13685 47903 13719
rect 49433 13685 49467 13719
rect 49801 13685 49835 13719
rect 51549 13685 51583 13719
rect 23397 13481 23431 13515
rect 23949 13481 23983 13515
rect 29653 13481 29687 13515
rect 31953 13481 31987 13515
rect 39221 13481 39255 13515
rect 39405 13481 39439 13515
rect 41981 13481 42015 13515
rect 44787 13481 44821 13515
rect 48329 13481 48363 13515
rect 48789 13481 48823 13515
rect 49801 13481 49835 13515
rect 51273 13481 51307 13515
rect 24961 13413 24995 13447
rect 32045 13413 32079 13447
rect 39497 13413 39531 13447
rect 47225 13413 47259 13447
rect 25513 13345 25547 13379
rect 30941 13345 30975 13379
rect 31585 13345 31619 13379
rect 39589 13345 39623 13379
rect 42901 13345 42935 13379
rect 43361 13345 43395 13379
rect 45477 13345 45511 13379
rect 50905 13345 50939 13379
rect 1593 13277 1627 13311
rect 23581 13277 23615 13311
rect 23857 13277 23891 13311
rect 25145 13277 25179 13311
rect 29653 13277 29687 13311
rect 29837 13277 29871 13311
rect 30021 13277 30055 13311
rect 31769 13277 31803 13311
rect 32229 13277 32263 13311
rect 32321 13277 32355 13311
rect 32413 13277 32447 13311
rect 33149 13277 33183 13311
rect 35081 13277 35115 13311
rect 37105 13277 37139 13311
rect 38669 13277 38703 13311
rect 39313 13277 39347 13311
rect 39865 13277 39899 13311
rect 41981 13277 42015 13311
rect 42165 13277 42199 13311
rect 42349 13277 42383 13311
rect 42993 13277 43027 13311
rect 47777 13277 47811 13311
rect 47961 13277 47995 13311
rect 48237 13277 48271 13311
rect 48513 13277 48547 13311
rect 48605 13277 48639 13311
rect 48881 13277 48915 13311
rect 48973 13277 49007 13311
rect 49157 13277 49191 13311
rect 49433 13277 49467 13311
rect 49525 13277 49559 13311
rect 49617 13277 49651 13311
rect 51089 13277 51123 13311
rect 51365 13277 51399 13311
rect 51549 13277 51583 13311
rect 51733 13277 51767 13311
rect 52009 13277 52043 13311
rect 24869 13209 24903 13243
rect 25053 13209 25087 13243
rect 25789 13209 25823 13243
rect 27537 13209 27571 13243
rect 31493 13209 31527 13243
rect 32045 13209 32079 13243
rect 33416 13209 33450 13243
rect 35348 13209 35382 13243
rect 37372 13209 37406 13243
rect 40132 13209 40166 13243
rect 45753 13209 45787 13243
rect 47869 13209 47903 13243
rect 48099 13209 48133 13243
rect 49065 13209 49099 13243
rect 51641 13209 51675 13243
rect 52285 13209 52319 13243
rect 30573 13141 30607 13175
rect 33057 13141 33091 13175
rect 34529 13141 34563 13175
rect 36461 13141 36495 13175
rect 38485 13141 38519 13175
rect 41245 13141 41279 13175
rect 47593 13141 47627 13175
rect 51917 13141 51951 13175
rect 53757 13141 53791 13175
rect 24777 12937 24811 12971
rect 26709 12937 26743 12971
rect 30481 12937 30515 12971
rect 31217 12937 31251 12971
rect 34069 12937 34103 12971
rect 36277 12937 36311 12971
rect 37657 12937 37691 12971
rect 39037 12937 39071 12971
rect 41061 12937 41095 12971
rect 41245 12937 41279 12971
rect 43821 12937 43855 12971
rect 44557 12937 44591 12971
rect 45569 12937 45603 12971
rect 48789 12937 48823 12971
rect 53389 12937 53423 12971
rect 53573 12937 53607 12971
rect 24685 12869 24719 12903
rect 29276 12869 29310 12903
rect 34437 12869 34471 12903
rect 34647 12869 34681 12903
rect 36645 12869 36679 12903
rect 36855 12869 36889 12903
rect 38485 12869 38519 12903
rect 38853 12869 38887 12903
rect 39957 12869 39991 12903
rect 42686 12869 42720 12903
rect 44189 12869 44223 12903
rect 49065 12869 49099 12903
rect 51917 12869 51951 12903
rect 25145 12801 25179 12835
rect 25605 12801 25639 12835
rect 26525 12801 26559 12835
rect 26801 12801 26835 12835
rect 26985 12801 27019 12835
rect 27537 12801 27571 12835
rect 27804 12801 27838 12835
rect 29009 12801 29043 12835
rect 30665 12801 30699 12835
rect 30941 12801 30975 12835
rect 31125 12801 31159 12835
rect 31217 12801 31251 12835
rect 31769 12801 31803 12835
rect 32137 12801 32171 12835
rect 32873 12801 32907 12835
rect 33057 12801 33091 12835
rect 34345 12801 34379 12835
rect 34529 12801 34563 12835
rect 36553 12801 36587 12835
rect 36737 12801 36771 12835
rect 37013 12801 37047 12835
rect 37289 12801 37323 12835
rect 37473 12801 37507 12835
rect 37565 12801 37599 12835
rect 37841 12801 37875 12835
rect 37933 12801 37967 12835
rect 38117 12801 38151 12835
rect 38945 12801 38979 12835
rect 39129 12801 39163 12835
rect 39865 12801 39899 12835
rect 40050 12801 40084 12835
rect 40167 12801 40201 12835
rect 40325 12801 40359 12835
rect 41429 12801 41463 12835
rect 43913 12801 43947 12835
rect 44465 12801 44499 12835
rect 45753 12801 45787 12835
rect 46029 12801 46063 12835
rect 49617 12801 49651 12835
rect 49801 12801 49835 12835
rect 50077 12801 50111 12835
rect 52101 12801 52135 12835
rect 52837 12801 52871 12835
rect 53481 12801 53515 12835
rect 22661 12733 22695 12767
rect 22937 12733 22971 12767
rect 25237 12733 25271 12767
rect 25421 12733 25455 12767
rect 31493 12733 31527 12767
rect 31585 12733 31619 12767
rect 33517 12733 33551 12767
rect 34161 12733 34195 12767
rect 34805 12733 34839 12767
rect 35725 12733 35759 12767
rect 36369 12733 36403 12767
rect 40417 12733 40451 12767
rect 42441 12733 42475 12767
rect 45937 12733 45971 12767
rect 48237 12733 48271 12767
rect 49341 12733 49375 12767
rect 49433 12733 49467 12767
rect 49985 12733 50019 12767
rect 51273 12733 51307 12767
rect 52285 12733 52319 12767
rect 30389 12665 30423 12699
rect 30757 12665 30791 12699
rect 30849 12665 30883 12699
rect 31309 12665 31343 12699
rect 39681 12665 39715 12699
rect 50445 12665 50479 12699
rect 26249 12597 26283 12631
rect 26341 12597 26375 12631
rect 27077 12597 27111 12631
rect 27445 12597 27479 12631
rect 28917 12597 28951 12631
rect 31953 12597 31987 12631
rect 32781 12597 32815 12631
rect 33241 12597 33275 12631
rect 37289 12597 37323 12631
rect 37933 12597 37967 12631
rect 49525 12597 49559 12631
rect 51825 12597 51859 12631
rect 23673 12393 23707 12427
rect 24501 12393 24535 12427
rect 26617 12393 26651 12427
rect 38393 12393 38427 12427
rect 38853 12393 38887 12427
rect 47961 12393 47995 12427
rect 51273 12393 51307 12427
rect 51457 12393 51491 12427
rect 25145 12257 25179 12291
rect 26985 12257 27019 12291
rect 29561 12257 29595 12291
rect 32597 12257 32631 12291
rect 33057 12257 33091 12291
rect 33149 12257 33183 12291
rect 37105 12257 37139 12291
rect 40969 12257 41003 12291
rect 43085 12257 43119 12291
rect 46213 12257 46247 12291
rect 46489 12257 46523 12291
rect 50445 12257 50479 12291
rect 50537 12257 50571 12291
rect 23581 12189 23615 12223
rect 24685 12189 24719 12223
rect 24777 12189 24811 12223
rect 26525 12189 26559 12223
rect 27445 12189 27479 12223
rect 29193 12189 29227 12223
rect 29377 12189 29411 12223
rect 30389 12189 30423 12223
rect 31033 12189 31067 12223
rect 32045 12189 32079 12223
rect 32873 12189 32907 12223
rect 32965 12189 32999 12223
rect 33609 12189 33643 12223
rect 33793 12189 33827 12223
rect 34713 12189 34747 12223
rect 36277 12189 36311 12223
rect 37841 12189 37875 12223
rect 39221 12189 39255 12223
rect 40601 12189 40635 12223
rect 40693 12189 40727 12223
rect 40877 12189 40911 12223
rect 41705 12189 41739 12223
rect 42533 12189 42567 12223
rect 45017 12189 45051 12223
rect 50353 12189 50387 12223
rect 50629 12189 50663 12223
rect 51549 12189 51583 12223
rect 24869 12121 24903 12155
rect 25007 12121 25041 12155
rect 30941 12121 30975 12155
rect 34980 12121 35014 12155
rect 37657 12121 37691 12155
rect 38577 12121 38611 12155
rect 40325 12121 40359 12155
rect 42349 12121 42383 12155
rect 42809 12121 42843 12155
rect 43361 12121 43395 12155
rect 45109 12121 45143 12155
rect 51089 12121 51123 12155
rect 27261 12053 27295 12087
rect 27353 12053 27387 12087
rect 29285 12053 29319 12087
rect 30205 12053 30239 12087
rect 31677 12053 31711 12087
rect 32689 12053 32723 12087
rect 33701 12053 33735 12087
rect 36093 12053 36127 12087
rect 36921 12053 36955 12087
rect 39037 12053 39071 12087
rect 40423 12053 40457 12087
rect 40509 12053 40543 12087
rect 40785 12053 40819 12087
rect 41613 12053 41647 12087
rect 44833 12053 44867 12087
rect 50169 12053 50203 12087
rect 51289 12053 51323 12087
rect 51641 12053 51675 12087
rect 25973 11849 26007 11883
rect 27353 11849 27387 11883
rect 31039 11849 31073 11883
rect 31125 11849 31159 11883
rect 35173 11849 35207 11883
rect 38669 11849 38703 11883
rect 40233 11849 40267 11883
rect 42165 11849 42199 11883
rect 44189 11849 44223 11883
rect 47133 11849 47167 11883
rect 49341 11849 49375 11883
rect 26249 11781 26283 11815
rect 26341 11781 26375 11815
rect 26985 11781 27019 11815
rect 29714 11781 29748 11815
rect 30941 11781 30975 11815
rect 33324 11781 33358 11815
rect 49893 11781 49927 11815
rect 50031 11781 50065 11815
rect 51641 11781 51675 11815
rect 51759 11781 51793 11815
rect 52009 11781 52043 11815
rect 24777 11713 24811 11747
rect 26157 11713 26191 11747
rect 26459 11713 26493 11747
rect 26617 11713 26651 11747
rect 27169 11713 27203 11747
rect 28089 11713 28123 11747
rect 31217 11713 31251 11747
rect 31309 11713 31343 11747
rect 31493 11713 31527 11747
rect 31585 11713 31619 11747
rect 31677 11713 31711 11747
rect 32413 11713 32447 11747
rect 35081 11713 35115 11747
rect 35265 11713 35299 11747
rect 35633 11713 35667 11747
rect 35909 11713 35943 11747
rect 36093 11713 36127 11747
rect 36277 11713 36311 11747
rect 37289 11713 37323 11747
rect 37556 11713 37590 11747
rect 38853 11713 38887 11747
rect 39120 11713 39154 11747
rect 40417 11713 40451 11747
rect 41061 11713 41095 11747
rect 41797 11713 41831 11747
rect 41981 11713 42015 11747
rect 44373 11713 44407 11747
rect 44925 11713 44959 11747
rect 45201 11713 45235 11747
rect 45385 11713 45419 11747
rect 47041 11713 47075 11747
rect 49709 11713 49743 11747
rect 49801 11713 49835 11747
rect 50169 11713 50203 11747
rect 51181 11713 51215 11747
rect 51457 11713 51491 11747
rect 51549 11713 51583 11747
rect 51917 11713 51951 11747
rect 52193 11713 52227 11747
rect 52745 11713 52779 11747
rect 52929 11713 52963 11747
rect 29469 11645 29503 11679
rect 33057 11645 33091 11679
rect 35449 11645 35483 11679
rect 36461 11645 36495 11679
rect 42441 11645 42475 11679
rect 44649 11645 44683 11679
rect 44741 11645 44775 11679
rect 47593 11645 47627 11679
rect 47869 11645 47903 11679
rect 50537 11645 50571 11679
rect 52377 11645 52411 11679
rect 40969 11577 41003 11611
rect 45201 11577 45235 11611
rect 52837 11577 52871 11611
rect 68477 11577 68511 11611
rect 24869 11509 24903 11543
rect 28273 11509 28307 11543
rect 30849 11509 30883 11543
rect 31309 11509 31343 11543
rect 32965 11509 32999 11543
rect 34437 11509 34471 11543
rect 35817 11509 35851 11543
rect 37013 11509 37047 11543
rect 41705 11509 41739 11543
rect 43085 11509 43119 11543
rect 44557 11509 44591 11543
rect 45109 11509 45143 11543
rect 49525 11509 49559 11543
rect 51273 11509 51307 11543
rect 26617 11305 26651 11339
rect 27169 11305 27203 11339
rect 27629 11305 27663 11339
rect 28365 11305 28399 11339
rect 36185 11305 36219 11339
rect 38761 11305 38795 11339
rect 39221 11305 39255 11339
rect 41245 11305 41279 11339
rect 45937 11305 45971 11339
rect 47317 11305 47351 11339
rect 49893 11305 49927 11339
rect 50800 11305 50834 11339
rect 26433 11237 26467 11271
rect 28733 11237 28767 11271
rect 30021 11237 30055 11271
rect 31125 11237 31159 11271
rect 46213 11237 46247 11271
rect 47777 11237 47811 11271
rect 47961 11237 47995 11271
rect 22385 11169 22419 11203
rect 22661 11169 22695 11203
rect 25605 11169 25639 11203
rect 25697 11169 25731 11203
rect 26249 11169 26283 11203
rect 29745 11169 29779 11203
rect 30113 11169 30147 11203
rect 30205 11169 30239 11203
rect 36369 11169 36403 11203
rect 37749 11169 37783 11203
rect 38209 11169 38243 11203
rect 38393 11169 38427 11203
rect 39865 11169 39899 11203
rect 46305 11169 46339 11203
rect 48421 11169 48455 11203
rect 48605 11169 48639 11203
rect 49525 11169 49559 11203
rect 52561 11169 52595 11203
rect 24777 11101 24811 11135
rect 25789 11101 25823 11135
rect 25881 11101 25915 11135
rect 26065 11101 26099 11135
rect 26157 11101 26191 11135
rect 26433 11101 26467 11135
rect 26525 11101 26559 11135
rect 26700 11101 26734 11135
rect 27353 11101 27387 11135
rect 27445 11101 27479 11135
rect 27905 11101 27939 11135
rect 28181 11101 28215 11135
rect 28457 11101 28491 11135
rect 28549 11101 28583 11135
rect 29929 11101 29963 11135
rect 30389 11101 30423 11135
rect 30573 11101 30607 11135
rect 31585 11101 31619 11135
rect 34805 11101 34839 11135
rect 37105 11101 37139 11135
rect 37933 11101 37967 11135
rect 38025 11101 38059 11135
rect 38117 11101 38151 11135
rect 38577 11101 38611 11135
rect 39221 11101 39255 11135
rect 39405 11101 39439 11135
rect 41521 11101 41555 11135
rect 41797 11101 41831 11135
rect 46121 11101 46155 11135
rect 46397 11101 46431 11135
rect 46581 11101 46615 11135
rect 47501 11101 47535 11135
rect 47685 11101 47719 11135
rect 49709 11101 49743 11135
rect 50537 11101 50571 11135
rect 27169 11033 27203 11067
rect 27721 11033 27755 11067
rect 28273 11033 28307 11067
rect 31852 11033 31886 11067
rect 35072 11033 35106 11067
rect 36921 11033 36955 11067
rect 40132 11033 40166 11067
rect 42064 11033 42098 11067
rect 48329 11033 48363 11067
rect 24133 10965 24167 10999
rect 25329 10965 25363 10999
rect 25421 10965 25455 10999
rect 28089 10965 28123 10999
rect 32965 10965 32999 10999
rect 37657 10965 37691 10999
rect 41613 10965 41647 10999
rect 43177 10965 43211 10999
rect 23581 10761 23615 10795
rect 24409 10761 24443 10795
rect 25329 10761 25363 10795
rect 25513 10761 25547 10795
rect 25697 10761 25731 10795
rect 25881 10761 25915 10795
rect 26801 10761 26835 10795
rect 27353 10761 27387 10795
rect 43085 10761 43119 10795
rect 44189 10761 44223 10795
rect 45017 10761 45051 10795
rect 50997 10761 51031 10795
rect 51457 10761 51491 10795
rect 24685 10693 24719 10727
rect 25421 10693 25455 10727
rect 27537 10693 27571 10727
rect 28365 10693 28399 10727
rect 29101 10693 29135 10727
rect 33977 10693 34011 10727
rect 40693 10693 40727 10727
rect 40785 10693 40819 10727
rect 41521 10693 41555 10727
rect 44281 10693 44315 10727
rect 49525 10693 49559 10727
rect 51181 10693 51215 10727
rect 23489 10625 23523 10659
rect 24593 10625 24627 10659
rect 24777 10625 24811 10659
rect 24915 10625 24949 10659
rect 25789 10625 25823 10659
rect 26617 10625 26651 10659
rect 26985 10625 27019 10659
rect 29745 10625 29779 10659
rect 33057 10625 33091 10659
rect 33333 10625 33367 10659
rect 33517 10625 33551 10659
rect 35357 10625 35391 10659
rect 36369 10625 36403 10659
rect 37381 10625 37415 10659
rect 37565 10625 37599 10659
rect 37657 10625 37691 10659
rect 37933 10625 37967 10659
rect 40233 10625 40267 10659
rect 40509 10625 40543 10659
rect 41889 10625 41923 10659
rect 41981 10631 42015 10665
rect 49249 10625 49283 10659
rect 51089 10625 51123 10659
rect 51365 10625 51399 10659
rect 25053 10557 25087 10591
rect 25145 10557 25179 10591
rect 26433 10557 26467 10591
rect 27261 10557 27295 10591
rect 27353 10557 27387 10591
rect 29193 10557 29227 10591
rect 29285 10557 29319 10591
rect 32873 10557 32907 10591
rect 34069 10557 34103 10591
rect 34253 10557 34287 10591
rect 35633 10557 35667 10591
rect 35817 10557 35851 10591
rect 36461 10557 36495 10591
rect 40325 10557 40359 10591
rect 42441 10557 42475 10591
rect 44465 10557 44499 10591
rect 45109 10557 45143 10591
rect 45293 10557 45327 10591
rect 28733 10489 28767 10523
rect 35449 10489 35483 10523
rect 40049 10489 40083 10523
rect 1593 10421 1627 10455
rect 27077 10421 27111 10455
rect 29561 10421 29595 10455
rect 33241 10421 33275 10455
rect 33333 10421 33367 10455
rect 33609 10421 33643 10455
rect 35357 10421 35391 10455
rect 37105 10421 37139 10455
rect 37841 10421 37875 10455
rect 42165 10421 42199 10455
rect 43821 10421 43855 10455
rect 44649 10421 44683 10455
rect 25697 10217 25731 10251
rect 32919 10217 32953 10251
rect 33425 10217 33459 10251
rect 38669 10217 38703 10251
rect 42073 10217 42107 10251
rect 44787 10217 44821 10251
rect 46121 10217 46155 10251
rect 46305 10217 46339 10251
rect 25881 10149 25915 10183
rect 34713 10149 34747 10183
rect 42349 10149 42383 10183
rect 42441 10149 42475 10183
rect 24685 10081 24719 10115
rect 26985 10081 27019 10115
rect 30389 10081 30423 10115
rect 31493 10081 31527 10115
rect 34345 10081 34379 10115
rect 35357 10081 35391 10115
rect 38393 10081 38427 10115
rect 39221 10081 39255 10115
rect 41061 10081 41095 10115
rect 42993 10081 43027 10115
rect 45293 10081 45327 10115
rect 45569 10081 45603 10115
rect 45937 10081 45971 10115
rect 47777 10081 47811 10115
rect 23949 10013 23983 10047
rect 24225 10013 24259 10047
rect 25973 10013 26007 10047
rect 26157 10013 26191 10047
rect 26709 10013 26743 10047
rect 26893 10013 26927 10047
rect 27169 10013 27203 10047
rect 27537 10013 27571 10047
rect 28549 10013 28583 10047
rect 28733 10013 28767 10047
rect 31125 10013 31159 10047
rect 33241 10013 33275 10047
rect 33517 10013 33551 10047
rect 33609 10013 33643 10047
rect 35817 10013 35851 10047
rect 37289 10013 37323 10047
rect 38209 10013 38243 10047
rect 40785 10013 40819 10047
rect 40877 10013 40911 10047
rect 40969 10013 41003 10047
rect 41337 10013 41371 10047
rect 42257 10013 42291 10047
rect 42533 10013 42567 10047
rect 42717 10013 42751 10047
rect 43361 10013 43395 10047
rect 45201 10013 45235 10047
rect 45661 10013 45695 10047
rect 46121 10013 46155 10047
rect 48237 10013 48271 10047
rect 50169 10013 50203 10047
rect 25513 9945 25547 9979
rect 28273 9945 28307 9979
rect 35081 9945 35115 9979
rect 36084 9945 36118 9979
rect 41981 9945 42015 9979
rect 47041 9945 47075 9979
rect 48053 9945 48087 9979
rect 23765 9877 23799 9911
rect 24133 9877 24167 9911
rect 25237 9877 25271 9911
rect 25713 9877 25747 9911
rect 26065 9877 26099 9911
rect 27353 9877 27387 9911
rect 28641 9877 28675 9911
rect 31033 9877 31067 9911
rect 33057 9877 33091 9911
rect 35173 9877 35207 9911
rect 37197 9877 37231 9911
rect 37381 9877 37415 9911
rect 37841 9877 37875 9911
rect 38301 9877 38335 9911
rect 39037 9877 39071 9911
rect 39129 9877 39163 9911
rect 40601 9877 40635 9911
rect 48421 9877 48455 9911
rect 50813 9877 50847 9911
rect 30757 9673 30791 9707
rect 30941 9673 30975 9707
rect 34529 9673 34563 9707
rect 36737 9673 36771 9707
rect 43361 9673 43395 9707
rect 50997 9673 51031 9707
rect 24685 9605 24719 9639
rect 25697 9605 25731 9639
rect 25897 9605 25931 9639
rect 26249 9605 26283 9639
rect 26617 9605 26651 9639
rect 29285 9605 29319 9639
rect 33057 9605 33091 9639
rect 35538 9605 35572 9639
rect 40500 9605 40534 9639
rect 44005 9605 44039 9639
rect 46305 9605 46339 9639
rect 48053 9605 48087 9639
rect 48191 9605 48225 9639
rect 51181 9605 51215 9639
rect 24501 9537 24535 9571
rect 24777 9537 24811 9571
rect 24869 9537 24903 9571
rect 25145 9537 25179 9571
rect 25329 9537 25363 9571
rect 25513 9537 25547 9571
rect 25605 9537 25639 9571
rect 26157 9537 26191 9571
rect 26341 9537 26375 9571
rect 26525 9537 26559 9571
rect 26709 9537 26743 9571
rect 27261 9537 27295 9571
rect 27445 9537 27479 9571
rect 27905 9537 27939 9571
rect 30849 9537 30883 9571
rect 31033 9537 31067 9571
rect 31125 9537 31159 9571
rect 32137 9537 32171 9571
rect 32229 9537 32263 9571
rect 34713 9537 34747 9571
rect 35725 9537 35759 9571
rect 35817 9537 35851 9571
rect 38025 9537 38059 9571
rect 38761 9537 38795 9571
rect 38945 9537 38979 9571
rect 39221 9537 39255 9571
rect 39589 9537 39623 9571
rect 39773 9537 39807 9571
rect 41705 9537 41739 9571
rect 41797 9537 41831 9571
rect 42441 9537 42475 9571
rect 43269 9537 43303 9571
rect 43453 9537 43487 9571
rect 43913 9537 43947 9571
rect 44925 9537 44959 9571
rect 45109 9537 45143 9571
rect 45845 9537 45879 9571
rect 46489 9537 46523 9571
rect 46581 9537 46615 9571
rect 47225 9537 47259 9571
rect 47869 9537 47903 9571
rect 47961 9537 47995 9571
rect 48329 9537 48363 9571
rect 49065 9537 49099 9571
rect 49249 9537 49283 9571
rect 51089 9537 51123 9571
rect 22569 9469 22603 9503
rect 22845 9469 22879 9503
rect 29009 9469 29043 9503
rect 31217 9469 31251 9503
rect 32781 9469 32815 9503
rect 34989 9469 35023 9503
rect 36093 9469 36127 9503
rect 38209 9469 38243 9503
rect 38853 9469 38887 9503
rect 39497 9469 39531 9503
rect 40233 9469 40267 9503
rect 41981 9469 42015 9503
rect 44281 9469 44315 9503
rect 45293 9469 45327 9503
rect 48421 9469 48455 9503
rect 25053 9401 25087 9435
rect 26065 9401 26099 9435
rect 41613 9401 41647 9435
rect 44833 9401 44867 9435
rect 46765 9401 46799 9435
rect 24317 9333 24351 9367
rect 25881 9333 25915 9367
rect 27261 9333 27295 9367
rect 27721 9333 27755 9367
rect 35541 9333 35575 9367
rect 39037 9333 39071 9367
rect 39405 9333 39439 9367
rect 39957 9333 39991 9367
rect 41705 9333 41739 9367
rect 43085 9333 43119 9367
rect 46029 9333 46063 9367
rect 46581 9333 46615 9367
rect 47317 9333 47351 9367
rect 47685 9333 47719 9367
rect 49506 9333 49540 9367
rect 23673 9129 23707 9163
rect 25513 9129 25547 9163
rect 25973 9129 26007 9163
rect 26157 9129 26191 9163
rect 26801 9129 26835 9163
rect 34437 9129 34471 9163
rect 36093 9129 36127 9163
rect 40122 9129 40156 9163
rect 46660 9129 46694 9163
rect 48145 9129 48179 9163
rect 49157 9129 49191 9163
rect 31677 9061 31711 9095
rect 36461 9061 36495 9095
rect 39267 9061 39301 9095
rect 43177 9061 43211 9095
rect 49709 9061 49743 9095
rect 24961 8993 24995 9027
rect 27445 8993 27479 9027
rect 27905 8993 27939 9027
rect 32137 8993 32171 9027
rect 39865 8993 39899 9027
rect 41797 8993 41831 9027
rect 43729 8993 43763 9027
rect 43913 8993 43947 9027
rect 44097 8993 44131 9027
rect 46397 8993 46431 9027
rect 23581 8925 23615 8959
rect 26433 8925 26467 8959
rect 26709 8925 26743 8959
rect 27169 8925 27203 8959
rect 27629 8925 27663 8959
rect 29561 8925 29595 8959
rect 30297 8925 30331 8959
rect 30564 8925 30598 8959
rect 33149 8925 33183 8959
rect 34345 8925 34379 8959
rect 35449 8925 35483 8959
rect 36277 8925 36311 8959
rect 36369 8925 36403 8959
rect 36553 8925 36587 8959
rect 36737 8925 36771 8959
rect 37473 8925 37507 8959
rect 37841 8925 37875 8959
rect 45109 8925 45143 8959
rect 45293 8925 45327 8959
rect 45569 8925 45603 8959
rect 45753 8925 45787 8959
rect 48605 8925 48639 8959
rect 48789 8925 48823 8959
rect 48881 8925 48915 8959
rect 48973 8925 49007 8959
rect 49617 8925 49651 8959
rect 49709 8925 49743 8959
rect 49893 8925 49927 8959
rect 68477 8925 68511 8959
rect 25789 8857 25823 8891
rect 26005 8857 26039 8891
rect 26249 8857 26283 8891
rect 27261 8857 27295 8891
rect 29653 8857 29687 8891
rect 33977 8857 34011 8891
rect 42064 8857 42098 8891
rect 43637 8857 43671 8891
rect 44741 8857 44775 8891
rect 49249 8857 49283 8891
rect 49433 8857 49467 8891
rect 26617 8789 26651 8823
rect 29377 8789 29411 8823
rect 32781 8789 32815 8823
rect 36001 8789 36035 8823
rect 41613 8789 41647 8823
rect 43269 8789 43303 8823
rect 45477 8789 45511 8823
rect 45937 8789 45971 8823
rect 32505 8585 32539 8619
rect 37933 8585 37967 8619
rect 38485 8585 38519 8619
rect 40693 8585 40727 8619
rect 48437 8585 48471 8619
rect 48605 8585 48639 8619
rect 48789 8585 48823 8619
rect 51273 8585 51307 8619
rect 23489 8517 23523 8551
rect 26617 8517 26651 8551
rect 27629 8517 27663 8551
rect 27905 8517 27939 8551
rect 28089 8517 28123 8551
rect 32597 8517 32631 8551
rect 39681 8517 39715 8551
rect 40877 8517 40911 8551
rect 41981 8517 42015 8551
rect 43361 8517 43395 8551
rect 45017 8517 45051 8551
rect 46397 8517 46431 8551
rect 48237 8517 48271 8551
rect 51549 8517 51583 8551
rect 23213 8449 23247 8483
rect 26433 8449 26467 8483
rect 26709 8449 26743 8483
rect 26985 8449 27019 8483
rect 27721 8449 27755 8483
rect 31033 8449 31067 8483
rect 33241 8449 33275 8483
rect 33885 8449 33919 8483
rect 34704 8449 34738 8483
rect 35909 8449 35943 8483
rect 36645 8449 36679 8483
rect 36829 8449 36863 8483
rect 37841 8449 37875 8483
rect 38025 8449 38059 8483
rect 38393 8449 38427 8483
rect 40601 8449 40635 8483
rect 41889 8449 41923 8483
rect 42073 8449 42107 8483
rect 42901 8449 42935 8483
rect 44925 8449 44959 8483
rect 45901 8449 45935 8483
rect 46029 8449 46063 8483
rect 46121 8449 46155 8483
rect 46305 8449 46339 8483
rect 48697 8449 48731 8483
rect 48881 8449 48915 8483
rect 51457 8449 51491 8483
rect 32781 8381 32815 8415
rect 33977 8381 34011 8415
rect 34437 8381 34471 8415
rect 39129 8381 39163 8415
rect 41613 8381 41647 8415
rect 43085 8381 43119 8415
rect 47133 8381 47167 8415
rect 49525 8381 49559 8415
rect 49801 8381 49835 8415
rect 24961 8313 24995 8347
rect 32137 8313 32171 8347
rect 35817 8313 35851 8347
rect 42717 8313 42751 8347
rect 44833 8313 44867 8347
rect 26249 8245 26283 8279
rect 30849 8245 30883 8279
rect 33333 8245 33367 8279
rect 36553 8245 36587 8279
rect 36645 8245 36679 8279
rect 48421 8245 48455 8279
rect 24501 8041 24535 8075
rect 27077 8041 27111 8075
rect 32137 8041 32171 8075
rect 34713 8041 34747 8075
rect 45845 8041 45879 8075
rect 46765 8041 46799 8075
rect 48145 8041 48179 8075
rect 48421 8041 48455 8075
rect 49617 8041 49651 8075
rect 37749 7973 37783 8007
rect 42349 7973 42383 8007
rect 46949 7973 46983 8007
rect 48789 7973 48823 8007
rect 25329 7905 25363 7939
rect 27629 7905 27663 7939
rect 29377 7905 29411 7939
rect 30389 7905 30423 7939
rect 32229 7905 32263 7939
rect 36369 7905 36403 7939
rect 38301 7905 38335 7939
rect 38485 7905 38519 7939
rect 38669 7905 38703 7939
rect 41409 7905 41443 7939
rect 41705 7905 41739 7939
rect 44097 7905 44131 7939
rect 47777 7905 47811 7939
rect 49341 7905 49375 7939
rect 1593 7837 1627 7871
rect 24409 7837 24443 7871
rect 29837 7837 29871 7871
rect 30021 7837 30055 7871
rect 32597 7837 32631 7871
rect 34713 7837 34747 7871
rect 34897 7837 34931 7871
rect 34989 7837 35023 7871
rect 35265 7837 35299 7871
rect 35357 7837 35391 7871
rect 36636 7837 36670 7871
rect 39589 7837 39623 7871
rect 41061 7837 41095 7871
rect 41245 7837 41279 7871
rect 41613 7837 41647 7871
rect 42441 7837 42475 7871
rect 43177 7837 43211 7871
rect 43545 7837 43579 7871
rect 46026 7837 46060 7871
rect 46397 7837 46431 7871
rect 46489 7837 46523 7871
rect 47501 7837 47535 7871
rect 47947 7847 47981 7881
rect 49801 7837 49835 7871
rect 25605 7769 25639 7803
rect 27905 7769 27939 7803
rect 30665 7769 30699 7803
rect 38209 7769 38243 7803
rect 39313 7769 39347 7803
rect 41337 7769 41371 7803
rect 41521 7769 41555 7803
rect 43085 7769 43119 7803
rect 46581 7769 46615 7803
rect 46781 7769 46815 7803
rect 47593 7769 47627 7803
rect 48237 7769 48271 7803
rect 48437 7769 48471 7803
rect 49249 7769 49283 7803
rect 29653 7701 29687 7735
rect 30113 7701 30147 7735
rect 34023 7701 34057 7735
rect 35087 7701 35121 7735
rect 35173 7701 35207 7735
rect 36001 7701 36035 7735
rect 37841 7701 37875 7735
rect 39405 7701 39439 7735
rect 41153 7701 41187 7735
rect 43269 7701 43303 7735
rect 46029 7701 46063 7735
rect 48605 7701 48639 7735
rect 49157 7701 49191 7735
rect 26341 7497 26375 7531
rect 28917 7497 28951 7531
rect 29285 7497 29319 7531
rect 31585 7497 31619 7531
rect 31953 7497 31987 7531
rect 32873 7497 32907 7531
rect 33425 7497 33459 7531
rect 33517 7497 33551 7531
rect 40141 7497 40175 7531
rect 42257 7497 42291 7531
rect 43821 7497 43855 7531
rect 44741 7497 44775 7531
rect 46305 7497 46339 7531
rect 47777 7497 47811 7531
rect 49709 7497 49743 7531
rect 30757 7429 30791 7463
rect 35164 7429 35198 7463
rect 38485 7429 38519 7463
rect 44833 7429 44867 7463
rect 45937 7429 45971 7463
rect 48145 7429 48179 7463
rect 48973 7429 49007 7463
rect 49433 7429 49467 7463
rect 46167 7395 46201 7429
rect 26249 7361 26283 7395
rect 28457 7361 28491 7395
rect 29101 7361 29135 7395
rect 29193 7361 29227 7395
rect 29469 7361 29503 7395
rect 29653 7361 29687 7395
rect 30205 7361 30239 7395
rect 30389 7361 30423 7395
rect 31493 7361 31527 7395
rect 31769 7361 31803 7395
rect 31953 7361 31987 7395
rect 38209 7361 38243 7395
rect 40049 7361 40083 7395
rect 40877 7361 40911 7395
rect 41144 7361 41178 7395
rect 42441 7361 42475 7395
rect 42697 7361 42731 7395
rect 46397 7361 46431 7395
rect 46673 7361 46707 7395
rect 46857 7361 46891 7395
rect 47961 7361 47995 7395
rect 48237 7361 48271 7395
rect 49249 7361 49283 7395
rect 49522 7383 49556 7417
rect 49617 7361 49651 7395
rect 49801 7361 49835 7395
rect 28549 7293 28583 7327
rect 28687 7293 28721 7327
rect 32229 7293 32263 7327
rect 33701 7293 33735 7327
rect 34897 7293 34931 7327
rect 36369 7293 36403 7327
rect 45017 7293 45051 7327
rect 48329 7293 48363 7327
rect 28089 7225 28123 7259
rect 44373 7225 44407 7259
rect 33057 7157 33091 7191
rect 36277 7157 36311 7191
rect 37013 7157 37047 7191
rect 39957 7157 39991 7191
rect 46121 7157 46155 7191
rect 46489 7157 46523 7191
rect 46673 7157 46707 7191
rect 49065 7157 49099 7191
rect 25868 6953 25902 6987
rect 29193 6953 29227 6987
rect 29745 6953 29779 6987
rect 36461 6953 36495 6987
rect 41889 6953 41923 6987
rect 43256 6953 43290 6987
rect 45017 6953 45051 6987
rect 48316 6953 48350 6987
rect 49801 6953 49835 6987
rect 27353 6817 27387 6851
rect 27905 6817 27939 6851
rect 29837 6817 29871 6851
rect 31585 6817 31619 6851
rect 35265 6817 35299 6851
rect 37657 6817 37691 6851
rect 42993 6817 43027 6851
rect 44741 6817 44775 6851
rect 45661 6817 45695 6851
rect 46397 6817 46431 6851
rect 46949 6817 46983 6851
rect 25605 6749 25639 6783
rect 27629 6749 27663 6783
rect 27721 6749 27755 6783
rect 28549 6749 28583 6783
rect 28641 6749 28675 6783
rect 28825 6749 28859 6783
rect 29009 6749 29043 6783
rect 29745 6749 29779 6783
rect 31769 6749 31803 6783
rect 33333 6749 33367 6783
rect 33517 6749 33551 6783
rect 33793 6749 33827 6783
rect 36369 6749 36403 6783
rect 37473 6749 37507 6783
rect 37749 6749 37783 6783
rect 38393 6749 38427 6783
rect 39957 6749 39991 6783
rect 40049 6749 40083 6783
rect 40417 6749 40451 6783
rect 40601 6749 40635 6783
rect 41889 6749 41923 6783
rect 42165 6749 42199 6783
rect 45201 6749 45235 6783
rect 45293 6749 45327 6783
rect 45845 6749 45879 6783
rect 46673 6749 46707 6783
rect 46765 6749 46799 6783
rect 46857 6749 46891 6783
rect 48053 6749 48087 6783
rect 27445 6681 27479 6715
rect 28917 6681 28951 6715
rect 35081 6681 35115 6715
rect 40509 6681 40543 6715
rect 42073 6681 42107 6715
rect 45385 6681 45419 6715
rect 45523 6681 45557 6715
rect 27543 6613 27577 6647
rect 30113 6613 30147 6647
rect 31953 6613 31987 6647
rect 33701 6613 33735 6647
rect 33885 6613 33919 6647
rect 34713 6613 34747 6647
rect 35173 6613 35207 6647
rect 37289 6613 37323 6647
rect 38945 6613 38979 6647
rect 40233 6613 40267 6647
rect 46489 6613 46523 6647
rect 26709 6409 26743 6443
rect 28825 6409 28859 6443
rect 29285 6409 29319 6443
rect 36093 6409 36127 6443
rect 38853 6409 38887 6443
rect 39129 6409 39163 6443
rect 40785 6409 40819 6443
rect 44281 6409 44315 6443
rect 45937 6409 45971 6443
rect 48789 6409 48823 6443
rect 28457 6341 28491 6375
rect 28917 6341 28951 6375
rect 29117 6341 29151 6375
rect 30021 6341 30055 6375
rect 38209 6341 38243 6375
rect 40509 6341 40543 6375
rect 41153 6341 41187 6375
rect 45569 6341 45603 6375
rect 46397 6341 46431 6375
rect 46765 6341 46799 6375
rect 46857 6341 46891 6375
rect 48605 6341 48639 6375
rect 26617 6273 26651 6307
rect 28641 6273 28675 6307
rect 29561 6273 29595 6307
rect 29653 6273 29687 6307
rect 29837 6273 29871 6307
rect 29929 6273 29963 6307
rect 30389 6273 30423 6307
rect 30481 6273 30515 6307
rect 30665 6273 30699 6307
rect 30941 6273 30975 6307
rect 31585 6273 31619 6307
rect 31769 6273 31803 6307
rect 35541 6273 35575 6307
rect 35725 6273 35759 6307
rect 35817 6273 35851 6307
rect 35909 6273 35943 6307
rect 36369 6273 36403 6307
rect 36462 6273 36496 6307
rect 36645 6273 36679 6307
rect 36737 6273 36771 6307
rect 36834 6273 36868 6307
rect 37473 6273 37507 6307
rect 38669 6273 38703 6307
rect 38945 6273 38979 6307
rect 40417 6273 40451 6307
rect 40601 6273 40635 6307
rect 44189 6273 44223 6307
rect 45753 6273 45787 6307
rect 46029 6273 46063 6307
rect 46489 6273 46523 6307
rect 46581 6273 46615 6307
rect 46949 6273 46983 6307
rect 48697 6273 48731 6307
rect 30297 6205 30331 6239
rect 31677 6205 31711 6239
rect 32781 6205 32815 6239
rect 33057 6205 33091 6239
rect 36093 6205 36127 6239
rect 37565 6205 37599 6239
rect 38485 6205 38519 6239
rect 41245 6205 41279 6239
rect 41429 6205 41463 6239
rect 48053 6205 48087 6239
rect 30205 6137 30239 6171
rect 35633 6137 35667 6171
rect 68477 6137 68511 6171
rect 29101 6069 29135 6103
rect 29377 6069 29411 6103
rect 31033 6069 31067 6103
rect 34529 6069 34563 6103
rect 37013 6069 37047 6103
rect 37841 6069 37875 6103
rect 38577 6069 38611 6103
rect 46213 6069 46247 6103
rect 47133 6069 47167 6103
rect 29653 5865 29687 5899
rect 30389 5865 30423 5899
rect 31309 5865 31343 5899
rect 33057 5865 33091 5899
rect 33425 5865 33459 5899
rect 36185 5865 36219 5899
rect 37289 5865 37323 5899
rect 37841 5865 37875 5899
rect 38853 5865 38887 5899
rect 39037 5865 39071 5899
rect 39405 5865 39439 5899
rect 40785 5865 40819 5899
rect 41521 5865 41555 5899
rect 46397 5865 46431 5899
rect 46765 5865 46799 5899
rect 48881 5865 48915 5899
rect 30021 5797 30055 5831
rect 38301 5797 38335 5831
rect 39221 5797 39255 5831
rect 40049 5797 40083 5831
rect 27169 5729 27203 5763
rect 27905 5729 27939 5763
rect 29929 5729 29963 5763
rect 30573 5729 30607 5763
rect 30757 5729 30791 5763
rect 31125 5729 31159 5763
rect 33517 5729 33551 5763
rect 33701 5729 33735 5763
rect 37381 5729 37415 5763
rect 38025 5729 38059 5763
rect 41705 5729 41739 5763
rect 45753 5729 45787 5763
rect 46857 5729 46891 5763
rect 47409 5729 47443 5763
rect 25421 5661 25455 5695
rect 28089 5661 28123 5695
rect 28273 5661 28307 5695
rect 28365 5661 28399 5695
rect 28549 5661 28583 5695
rect 29561 5661 29595 5695
rect 29837 5661 29871 5695
rect 30665 5661 30699 5695
rect 30849 5661 30883 5695
rect 31309 5661 31343 5695
rect 31585 5661 31619 5695
rect 31769 5661 31803 5695
rect 32321 5661 32355 5695
rect 32505 5661 32539 5695
rect 32623 5661 32657 5695
rect 32781 5661 32815 5695
rect 33241 5661 33275 5695
rect 33609 5661 33643 5695
rect 33793 5661 33827 5695
rect 36093 5661 36127 5695
rect 36369 5661 36403 5695
rect 37105 5661 37139 5695
rect 38117 5661 38151 5695
rect 38669 5661 38703 5695
rect 38853 5661 38887 5695
rect 39129 5661 39163 5695
rect 39313 5661 39347 5695
rect 39405 5661 39439 5695
rect 39589 5661 39623 5695
rect 40233 5661 40267 5695
rect 40509 5661 40543 5695
rect 43545 5661 43579 5695
rect 45937 5661 45971 5695
rect 46581 5661 46615 5695
rect 47133 5661 47167 5695
rect 48973 5661 49007 5695
rect 25697 5593 25731 5627
rect 27629 5593 27663 5627
rect 28181 5593 28215 5627
rect 31033 5593 31067 5627
rect 32413 5593 32447 5627
rect 36921 5593 36955 5627
rect 37841 5593 37875 5627
rect 40601 5593 40635 5627
rect 40801 5593 40835 5627
rect 41153 5593 41187 5627
rect 41337 5593 41371 5627
rect 41981 5593 42015 5627
rect 43637 5593 43671 5627
rect 49065 5593 49099 5627
rect 27261 5525 27295 5559
rect 27721 5525 27755 5559
rect 28549 5525 28583 5559
rect 31493 5525 31527 5559
rect 31953 5525 31987 5559
rect 32137 5525 32171 5559
rect 36461 5525 36495 5559
rect 40417 5525 40451 5559
rect 40969 5525 41003 5559
rect 43453 5525 43487 5559
rect 46121 5525 46155 5559
rect 25973 5321 26007 5355
rect 26525 5321 26559 5355
rect 29117 5321 29151 5355
rect 29469 5321 29503 5355
rect 30849 5321 30883 5355
rect 31309 5321 31343 5355
rect 31953 5321 31987 5355
rect 32965 5321 32999 5355
rect 33885 5321 33919 5355
rect 40693 5321 40727 5355
rect 41337 5321 41371 5355
rect 45661 5321 45695 5355
rect 27445 5253 27479 5287
rect 28273 5253 28307 5287
rect 28917 5253 28951 5287
rect 31769 5253 31803 5287
rect 36461 5253 36495 5287
rect 41153 5253 41187 5287
rect 43085 5253 43119 5287
rect 45753 5253 45787 5287
rect 47225 5253 47259 5287
rect 26157 5185 26191 5219
rect 26433 5185 26467 5219
rect 27261 5185 27295 5219
rect 27537 5185 27571 5219
rect 28365 5185 28399 5219
rect 28549 5185 28583 5219
rect 28733 5185 28767 5219
rect 28825 5185 28859 5219
rect 29377 5185 29411 5219
rect 30573 5185 30607 5219
rect 30665 5185 30699 5219
rect 31125 5185 31159 5219
rect 31585 5185 31619 5219
rect 32137 5185 32171 5219
rect 32873 5185 32907 5219
rect 33057 5185 33091 5219
rect 36277 5185 36311 5219
rect 39497 5185 39531 5219
rect 40509 5185 40543 5219
rect 40693 5185 40727 5219
rect 40969 5185 41003 5219
rect 41245 5185 41279 5219
rect 41521 5185 41555 5219
rect 46305 5185 46339 5219
rect 46397 5185 46431 5219
rect 46489 5185 46523 5219
rect 46607 5185 46641 5219
rect 46857 5185 46891 5219
rect 47041 5185 47075 5219
rect 47593 5185 47627 5219
rect 48329 5185 48363 5219
rect 48513 5185 48547 5219
rect 27629 5117 27663 5151
rect 30849 5117 30883 5151
rect 33333 5117 33367 5151
rect 34161 5117 34195 5151
rect 34437 5117 34471 5151
rect 36185 5117 36219 5151
rect 39313 5117 39347 5151
rect 42441 5117 42475 5151
rect 43453 5117 43487 5151
rect 43729 5117 43763 5151
rect 45937 5117 45971 5151
rect 46765 5117 46799 5151
rect 29285 5049 29319 5083
rect 45201 5049 45235 5083
rect 48237 5049 48271 5083
rect 27077 4981 27111 5015
rect 29101 4981 29135 5015
rect 32781 4981 32815 5015
rect 36645 4981 36679 5015
rect 39681 4981 39715 5015
rect 40785 4981 40819 5015
rect 45293 4981 45327 5015
rect 46121 4981 46155 5015
rect 48421 4981 48455 5015
rect 26052 4777 26086 4811
rect 27537 4777 27571 4811
rect 28181 4777 28215 4811
rect 30573 4777 30607 4811
rect 32124 4777 32158 4811
rect 33609 4777 33643 4811
rect 35081 4777 35115 4811
rect 36093 4777 36127 4811
rect 39497 4777 39531 4811
rect 42901 4777 42935 4811
rect 44005 4777 44039 4811
rect 44465 4777 44499 4811
rect 45832 4777 45866 4811
rect 28365 4709 28399 4743
rect 38117 4709 38151 4743
rect 25789 4641 25823 4675
rect 31861 4641 31895 4675
rect 37933 4641 37967 4675
rect 41429 4641 41463 4675
rect 45569 4641 45603 4675
rect 47777 4641 47811 4675
rect 30757 4573 30791 4607
rect 30941 4573 30975 4607
rect 31033 4573 31067 4607
rect 34989 4573 35023 4607
rect 35817 4573 35851 4607
rect 36001 4573 36035 4607
rect 36277 4573 36311 4607
rect 36369 4573 36403 4607
rect 36579 4573 36613 4607
rect 36737 4573 36771 4607
rect 36829 4573 36863 4607
rect 38025 4573 38059 4607
rect 38209 4573 38243 4607
rect 39865 4573 39899 4607
rect 40233 4573 40267 4607
rect 41153 4573 41187 4607
rect 42993 4573 43027 4607
rect 44189 4589 44223 4623
rect 44373 4573 44407 4607
rect 47593 4573 47627 4607
rect 47685 4573 47719 4607
rect 27997 4505 28031 4539
rect 28213 4505 28247 4539
rect 36461 4505 36495 4539
rect 37565 4505 37599 4539
rect 37749 4505 37783 4539
rect 39313 4505 39347 4539
rect 40049 4505 40083 4539
rect 40141 4505 40175 4539
rect 43085 4505 43119 4539
rect 36001 4437 36035 4471
rect 37473 4437 37507 4471
rect 39513 4437 39547 4471
rect 39681 4437 39715 4471
rect 40417 4437 40451 4471
rect 27077 4233 27111 4267
rect 38485 4233 38519 4267
rect 39497 4233 39531 4267
rect 30205 4165 30239 4199
rect 30323 4165 30357 4199
rect 36185 4165 36219 4199
rect 36415 4165 36449 4199
rect 37841 4165 37875 4199
rect 40509 4165 40543 4199
rect 40601 4165 40635 4199
rect 40785 4165 40819 4199
rect 26985 4097 27019 4131
rect 28549 4097 28583 4131
rect 30021 4097 30055 4131
rect 30113 4097 30147 4131
rect 32965 4097 32999 4131
rect 33885 4097 33919 4131
rect 36093 4097 36127 4131
rect 36277 4097 36311 4131
rect 36553 4097 36587 4131
rect 37749 4097 37783 4131
rect 37933 4097 37967 4131
rect 38051 4097 38085 4131
rect 38393 4097 38427 4131
rect 38577 4103 38611 4137
rect 39405 4097 39439 4131
rect 41061 4097 41095 4131
rect 28825 4029 28859 4063
rect 30481 4029 30515 4063
rect 30757 4029 30791 4063
rect 33057 4029 33091 4063
rect 34161 4029 34195 4063
rect 35909 4029 35943 4063
rect 38209 4029 38243 4063
rect 38669 4029 38703 4063
rect 39957 4029 39991 4063
rect 28641 3961 28675 3995
rect 31401 3961 31435 3995
rect 35633 3961 35667 3995
rect 39313 3961 39347 3995
rect 28733 3893 28767 3927
rect 29837 3893 29871 3927
rect 37565 3893 37599 3927
rect 40969 3893 41003 3927
rect 41153 3893 41187 3927
rect 30113 3689 30147 3723
rect 30757 3689 30791 3723
rect 31290 3689 31324 3723
rect 34805 3689 34839 3723
rect 38301 3689 38335 3723
rect 41797 3689 41831 3723
rect 30297 3621 30331 3655
rect 30941 3621 30975 3655
rect 38209 3621 38243 3655
rect 28733 3553 28767 3587
rect 31033 3553 31067 3587
rect 36553 3553 36587 3587
rect 37657 3553 37691 3587
rect 38761 3553 38795 3587
rect 40049 3553 40083 3587
rect 28273 3485 28307 3519
rect 28365 3485 28399 3519
rect 28825 3485 28859 3519
rect 29009 3485 29043 3519
rect 30021 3485 30055 3519
rect 30481 3485 30515 3519
rect 34713 3485 34747 3519
rect 36277 3485 36311 3519
rect 38025 3485 38059 3519
rect 38485 3485 38519 3519
rect 38577 3485 38611 3519
rect 38669 3485 38703 3519
rect 39129 3485 39163 3519
rect 68477 3485 68511 3519
rect 28641 3417 28675 3451
rect 30573 3417 30607 3451
rect 30789 3417 30823 3451
rect 33057 3417 33091 3451
rect 36369 3417 36403 3451
rect 37841 3417 37875 3451
rect 37933 3417 37967 3451
rect 40325 3417 40359 3451
rect 28089 3349 28123 3383
rect 29193 3349 29227 3383
rect 35909 3349 35943 3383
rect 39681 3349 39715 3383
rect 31217 3145 31251 3179
rect 31585 3145 31619 3179
rect 31677 3145 31711 3179
rect 32229 3145 32263 3179
rect 39037 3145 39071 3179
rect 27721 3077 27755 3111
rect 29653 3077 29687 3111
rect 37105 3077 37139 3111
rect 27445 3009 27479 3043
rect 29377 3009 29411 3043
rect 32137 3009 32171 3043
rect 32689 3009 32723 3043
rect 39129 3009 39163 3043
rect 39313 3009 39347 3043
rect 39681 3009 39715 3043
rect 47777 3009 47811 3043
rect 31125 2941 31159 2975
rect 31769 2941 31803 2975
rect 35081 2941 35115 2975
rect 35357 2941 35391 2975
rect 37289 2941 37323 2975
rect 37565 2941 37599 2975
rect 39957 2941 39991 2975
rect 29193 2873 29227 2907
rect 32873 2805 32907 2839
rect 39129 2805 39163 2839
rect 41429 2805 41463 2839
rect 47593 2805 47627 2839
rect 28549 2601 28583 2635
rect 30389 2601 30423 2635
rect 35633 2601 35667 2635
rect 36277 2601 36311 2635
rect 38301 2601 38335 2635
rect 39681 2601 39715 2635
rect 40693 2601 40727 2635
rect 1869 2533 1903 2567
rect 36093 2533 36127 2567
rect 68017 2465 68051 2499
rect 1593 2397 1627 2431
rect 2237 2397 2271 2431
rect 4813 2397 4847 2431
rect 7389 2397 7423 2431
rect 9965 2397 9999 2431
rect 17693 2397 17727 2431
rect 25421 2397 25455 2431
rect 28457 2397 28491 2431
rect 30297 2397 30331 2431
rect 30757 2397 30791 2431
rect 33149 2397 33183 2431
rect 35817 2397 35851 2431
rect 36185 2397 36219 2431
rect 38209 2397 38243 2431
rect 38669 2397 38703 2431
rect 39129 2397 39163 2431
rect 39405 2397 39439 2431
rect 39497 2397 39531 2431
rect 40601 2397 40635 2431
rect 43453 2397 43487 2431
rect 46029 2397 46063 2431
rect 48513 2397 48547 2431
rect 51181 2397 51215 2431
rect 53757 2397 53791 2431
rect 56333 2397 56367 2431
rect 58909 2397 58943 2431
rect 66637 2397 66671 2431
rect 68477 2397 68511 2431
rect 12449 2329 12483 2363
rect 39313 2329 39347 2363
rect 12541 2261 12575 2295
rect 48605 2261 48639 2295
<< metal1 >>
rect 1104 67482 68816 67504
rect 1104 67430 19574 67482
rect 19626 67430 19638 67482
rect 19690 67430 19702 67482
rect 19754 67430 19766 67482
rect 19818 67430 19830 67482
rect 19882 67430 50294 67482
rect 50346 67430 50358 67482
rect 50410 67430 50422 67482
rect 50474 67430 50486 67482
rect 50538 67430 50550 67482
rect 50602 67430 68816 67482
rect 1104 67408 68816 67430
rect 56134 67328 56140 67380
rect 56192 67328 56198 67380
rect 934 67192 940 67244
rect 992 67232 998 67244
rect 1581 67235 1639 67241
rect 1581 67232 1593 67235
rect 992 67204 1593 67232
rect 992 67192 998 67204
rect 1581 67201 1593 67204
rect 1627 67201 1639 67235
rect 1581 67195 1639 67201
rect 2222 67192 2228 67244
rect 2280 67192 2286 67244
rect 4798 67192 4804 67244
rect 4856 67192 4862 67244
rect 7374 67192 7380 67244
rect 7432 67192 7438 67244
rect 9950 67192 9956 67244
rect 10008 67192 10014 67244
rect 12434 67192 12440 67244
rect 12492 67232 12498 67244
rect 12529 67235 12587 67241
rect 12529 67232 12541 67235
rect 12492 67204 12541 67232
rect 12492 67192 12498 67204
rect 12529 67201 12541 67204
rect 12575 67201 12587 67235
rect 12529 67195 12587 67201
rect 15102 67192 15108 67244
rect 15160 67192 15166 67244
rect 17678 67192 17684 67244
rect 17736 67192 17742 67244
rect 20254 67192 20260 67244
rect 20312 67192 20318 67244
rect 22830 67192 22836 67244
rect 22888 67192 22894 67244
rect 25406 67192 25412 67244
rect 25464 67192 25470 67244
rect 27982 67192 27988 67244
rect 28040 67192 28046 67244
rect 30374 67192 30380 67244
rect 30432 67232 30438 67244
rect 30561 67235 30619 67241
rect 30561 67232 30573 67235
rect 30432 67204 30573 67232
rect 30432 67192 30438 67204
rect 30561 67201 30573 67204
rect 30607 67201 30619 67235
rect 30561 67195 30619 67201
rect 33134 67192 33140 67244
rect 33192 67192 33198 67244
rect 38286 67192 38292 67244
rect 38344 67192 38350 67244
rect 40862 67192 40868 67244
rect 40920 67192 40926 67244
rect 46014 67192 46020 67244
rect 46072 67192 46078 67244
rect 53742 67192 53748 67244
rect 53800 67192 53806 67244
rect 58894 67192 58900 67244
rect 58952 67192 58958 67244
rect 61470 67192 61476 67244
rect 61528 67192 61534 67244
rect 64046 67192 64052 67244
rect 64104 67192 64110 67244
rect 68465 67235 68523 67241
rect 68465 67201 68477 67235
rect 68511 67232 68523 67235
rect 68922 67232 68928 67244
rect 68511 67204 68928 67232
rect 68511 67201 68523 67204
rect 68465 67195 68523 67201
rect 68922 67192 68928 67204
rect 68980 67192 68986 67244
rect 1104 66938 68816 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 68816 66938
rect 1104 66864 68816 66886
rect 1104 66394 68816 66416
rect 1104 66342 19574 66394
rect 19626 66342 19638 66394
rect 19690 66342 19702 66394
rect 19754 66342 19766 66394
rect 19818 66342 19830 66394
rect 19882 66342 50294 66394
rect 50346 66342 50358 66394
rect 50410 66342 50422 66394
rect 50474 66342 50486 66394
rect 50538 66342 50550 66394
rect 50602 66342 68816 66394
rect 1104 66320 68816 66342
rect 68462 65968 68468 66020
rect 68520 65968 68526 66020
rect 1104 65850 68816 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 68816 65850
rect 1104 65776 68816 65798
rect 1104 65306 68816 65328
rect 1104 65254 19574 65306
rect 19626 65254 19638 65306
rect 19690 65254 19702 65306
rect 19754 65254 19766 65306
rect 19818 65254 19830 65306
rect 19882 65254 50294 65306
rect 50346 65254 50358 65306
rect 50410 65254 50422 65306
rect 50474 65254 50486 65306
rect 50538 65254 50550 65306
rect 50602 65254 68816 65306
rect 1104 65232 68816 65254
rect 1578 64880 1584 64932
rect 1636 64880 1642 64932
rect 1104 64762 68816 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 34934 64762
rect 34986 64710 34998 64762
rect 35050 64710 35062 64762
rect 35114 64710 35126 64762
rect 35178 64710 35190 64762
rect 35242 64710 65654 64762
rect 65706 64710 65718 64762
rect 65770 64710 65782 64762
rect 65834 64710 65846 64762
rect 65898 64710 65910 64762
rect 65962 64710 68816 64762
rect 1104 64688 68816 64710
rect 1104 64218 68816 64240
rect 1104 64166 19574 64218
rect 19626 64166 19638 64218
rect 19690 64166 19702 64218
rect 19754 64166 19766 64218
rect 19818 64166 19830 64218
rect 19882 64166 50294 64218
rect 50346 64166 50358 64218
rect 50410 64166 50422 64218
rect 50474 64166 50486 64218
rect 50538 64166 50550 64218
rect 50602 64166 68816 64218
rect 1104 64144 68816 64166
rect 1104 63674 68816 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 34934 63674
rect 34986 63622 34998 63674
rect 35050 63622 35062 63674
rect 35114 63622 35126 63674
rect 35178 63622 35190 63674
rect 35242 63622 65654 63674
rect 65706 63622 65718 63674
rect 65770 63622 65782 63674
rect 65834 63622 65846 63674
rect 65898 63622 65910 63674
rect 65962 63622 68816 63674
rect 1104 63600 68816 63622
rect 68462 63316 68468 63368
rect 68520 63316 68526 63368
rect 1104 63130 68816 63152
rect 1104 63078 19574 63130
rect 19626 63078 19638 63130
rect 19690 63078 19702 63130
rect 19754 63078 19766 63130
rect 19818 63078 19830 63130
rect 19882 63078 50294 63130
rect 50346 63078 50358 63130
rect 50410 63078 50422 63130
rect 50474 63078 50486 63130
rect 50538 63078 50550 63130
rect 50602 63078 68816 63130
rect 1104 63056 68816 63078
rect 1104 62586 68816 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 34934 62586
rect 34986 62534 34998 62586
rect 35050 62534 35062 62586
rect 35114 62534 35126 62586
rect 35178 62534 35190 62586
rect 35242 62534 65654 62586
rect 65706 62534 65718 62586
rect 65770 62534 65782 62586
rect 65834 62534 65846 62586
rect 65898 62534 65910 62586
rect 65962 62534 68816 62586
rect 1104 62512 68816 62534
rect 1104 62042 68816 62064
rect 1104 61990 19574 62042
rect 19626 61990 19638 62042
rect 19690 61990 19702 62042
rect 19754 61990 19766 62042
rect 19818 61990 19830 62042
rect 19882 61990 50294 62042
rect 50346 61990 50358 62042
rect 50410 61990 50422 62042
rect 50474 61990 50486 62042
rect 50538 61990 50550 62042
rect 50602 61990 68816 62042
rect 1104 61968 68816 61990
rect 1104 61498 68816 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 65654 61498
rect 65706 61446 65718 61498
rect 65770 61446 65782 61498
rect 65834 61446 65846 61498
rect 65898 61446 65910 61498
rect 65962 61446 68816 61498
rect 1104 61424 68816 61446
rect 1104 60954 68816 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 68816 60954
rect 1104 60880 68816 60902
rect 67821 60707 67879 60713
rect 67821 60673 67833 60707
rect 67867 60704 67879 60707
rect 68186 60704 68192 60716
rect 67867 60676 68192 60704
rect 67867 60673 67879 60676
rect 67821 60667 67879 60673
rect 68186 60664 68192 60676
rect 68244 60664 68250 60716
rect 68370 60528 68376 60580
rect 68428 60528 68434 60580
rect 1104 60410 68816 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 65654 60410
rect 65706 60358 65718 60410
rect 65770 60358 65782 60410
rect 65834 60358 65846 60410
rect 65898 60358 65910 60410
rect 65962 60358 68816 60410
rect 1104 60336 68816 60358
rect 1104 59866 68816 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 68816 59866
rect 1104 59792 68816 59814
rect 1578 59372 1584 59424
rect 1636 59372 1642 59424
rect 1104 59322 68816 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 65654 59322
rect 65706 59270 65718 59322
rect 65770 59270 65782 59322
rect 65834 59270 65846 59322
rect 65898 59270 65910 59322
rect 65962 59270 68816 59322
rect 1104 59248 68816 59270
rect 1104 58778 68816 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 68816 58778
rect 1104 58704 68816 58726
rect 1104 58234 68816 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 65654 58234
rect 65706 58182 65718 58234
rect 65770 58182 65782 58234
rect 65834 58182 65846 58234
rect 65898 58182 65910 58234
rect 65962 58182 68816 58234
rect 1104 58160 68816 58182
rect 68462 57876 68468 57928
rect 68520 57876 68526 57928
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 1578 56788 1584 56840
rect 1636 56788 1642 56840
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 68462 55088 68468 55140
rect 68520 55088 68526 55140
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 68462 52436 68468 52488
rect 68520 52436 68526 52488
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 934 51348 940 51400
rect 992 51388 998 51400
rect 1581 51391 1639 51397
rect 1581 51388 1593 51391
rect 992 51360 1593 51388
rect 992 51348 998 51360
rect 1581 51357 1593 51360
rect 1627 51357 1639 51391
rect 1581 51351 1639 51357
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 68462 49716 68468 49768
rect 68520 49716 68526 49768
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 934 48492 940 48544
rect 992 48532 998 48544
rect 1581 48535 1639 48541
rect 1581 48532 1593 48535
rect 992 48504 1593 48532
rect 992 48492 998 48504
rect 1581 48501 1593 48504
rect 1627 48501 1639 48535
rect 1581 48495 1639 48501
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 68462 46996 68468 47048
rect 68520 46996 68526 47048
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 934 45908 940 45960
rect 992 45948 998 45960
rect 1581 45951 1639 45957
rect 1581 45948 1593 45951
rect 992 45920 1593 45948
rect 992 45908 998 45920
rect 1581 45917 1593 45920
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 68462 44208 68468 44260
rect 68520 44208 68526 44260
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 934 43052 940 43104
rect 992 43092 998 43104
rect 1581 43095 1639 43101
rect 1581 43092 1593 43095
rect 992 43064 1593 43092
rect 992 43052 998 43064
rect 1581 43061 1593 43064
rect 1627 43061 1639 43095
rect 1581 43055 1639 43061
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 68462 41556 68468 41608
rect 68520 41556 68526 41608
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 934 37612 940 37664
rect 992 37652 998 37664
rect 1581 37655 1639 37661
rect 1581 37652 1593 37655
rect 992 37624 1593 37652
rect 992 37612 998 37624
rect 1581 37621 1593 37624
rect 1627 37621 1639 37655
rect 1581 37615 1639 37621
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 68462 36116 68468 36168
rect 68520 36116 68526 36168
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 934 35028 940 35080
rect 992 35068 998 35080
rect 1581 35071 1639 35077
rect 1581 35068 1593 35071
rect 992 35040 1593 35068
rect 992 35028 998 35040
rect 1581 35037 1593 35040
rect 1627 35037 1639 35071
rect 1581 35031 1639 35037
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 68281 33507 68339 33513
rect 68281 33473 68293 33507
rect 68327 33504 68339 33507
rect 68738 33504 68744 33516
rect 68327 33476 68744 33504
rect 68327 33473 68339 33476
rect 68281 33467 68339 33473
rect 68738 33464 68744 33476
rect 68796 33464 68802 33516
rect 68370 33260 68376 33312
rect 68428 33260 68434 33312
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 934 32172 940 32224
rect 992 32212 998 32224
rect 1581 32215 1639 32221
rect 1581 32212 1593 32215
rect 992 32184 1593 32212
rect 992 32172 998 32184
rect 1581 32181 1593 32184
rect 1627 32181 1639 32215
rect 1581 32175 1639 32181
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 68462 30676 68468 30728
rect 68520 30676 68526 30728
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 934 29588 940 29640
rect 992 29628 998 29640
rect 1581 29631 1639 29637
rect 1581 29628 1593 29631
rect 992 29600 1593 29628
rect 992 29588 998 29600
rect 1581 29597 1593 29600
rect 1627 29597 1639 29631
rect 1581 29591 1639 29597
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 68462 27888 68468 27940
rect 68520 27888 68526 27940
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 934 26732 940 26784
rect 992 26772 998 26784
rect 1581 26775 1639 26781
rect 1581 26772 1593 26775
rect 992 26744 1593 26772
rect 992 26732 998 26744
rect 1581 26741 1593 26744
rect 1627 26741 1639 26775
rect 1581 26735 1639 26741
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25245 28779 25279
rect 28721 25239 28779 25245
rect 28736 25208 28764 25239
rect 28902 25236 28908 25288
rect 28960 25236 28966 25288
rect 31202 25236 31208 25288
rect 31260 25236 31266 25288
rect 68462 25236 68468 25288
rect 68520 25236 68526 25288
rect 29546 25208 29552 25220
rect 28736 25180 29552 25208
rect 29546 25168 29552 25180
rect 29604 25168 29610 25220
rect 28810 25100 28816 25152
rect 28868 25100 28874 25152
rect 30926 25100 30932 25152
rect 30984 25140 30990 25152
rect 31757 25143 31815 25149
rect 31757 25140 31769 25143
rect 30984 25112 31769 25140
rect 30984 25100 30990 25112
rect 31757 25109 31769 25112
rect 31803 25109 31815 25143
rect 31757 25103 31815 25109
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 31202 24896 31208 24948
rect 31260 24936 31266 24948
rect 31389 24939 31447 24945
rect 31389 24936 31401 24939
rect 31260 24908 31401 24936
rect 31260 24896 31266 24908
rect 31389 24905 31401 24908
rect 31435 24936 31447 24939
rect 31662 24936 31668 24948
rect 31435 24908 31668 24936
rect 31435 24905 31447 24908
rect 31389 24899 31447 24905
rect 31662 24896 31668 24908
rect 31720 24896 31726 24948
rect 28436 24871 28494 24877
rect 28436 24837 28448 24871
rect 28482 24868 28494 24871
rect 28810 24868 28816 24880
rect 28482 24840 28816 24868
rect 28482 24837 28494 24840
rect 28436 24831 28494 24837
rect 28810 24828 28816 24840
rect 28868 24828 28874 24880
rect 34054 24868 34060 24880
rect 33980 24840 34060 24868
rect 30282 24809 30288 24812
rect 30276 24763 30288 24809
rect 30282 24760 30288 24763
rect 30340 24760 30346 24812
rect 31846 24760 31852 24812
rect 31904 24800 31910 24812
rect 32490 24800 32496 24812
rect 31904 24772 32496 24800
rect 31904 24760 31910 24772
rect 32490 24760 32496 24772
rect 32548 24800 32554 24812
rect 33980 24809 34008 24840
rect 34054 24828 34060 24840
rect 34112 24868 34118 24880
rect 34112 24840 35480 24868
rect 34112 24828 34118 24840
rect 34238 24809 34244 24812
rect 33965 24803 34023 24809
rect 33965 24800 33977 24803
rect 32548 24772 33977 24800
rect 32548 24760 32554 24772
rect 33965 24769 33977 24772
rect 34011 24769 34023 24803
rect 33965 24763 34023 24769
rect 34232 24763 34244 24809
rect 34238 24760 34244 24763
rect 34296 24760 34302 24812
rect 35452 24809 35480 24840
rect 35437 24803 35495 24809
rect 35437 24769 35449 24803
rect 35483 24769 35495 24803
rect 35437 24763 35495 24769
rect 35704 24803 35762 24809
rect 35704 24769 35716 24803
rect 35750 24800 35762 24803
rect 36078 24800 36084 24812
rect 35750 24772 36084 24800
rect 35750 24769 35762 24772
rect 35704 24763 35762 24769
rect 36078 24760 36084 24772
rect 36136 24760 36142 24812
rect 28169 24735 28227 24741
rect 28169 24701 28181 24735
rect 28215 24701 28227 24735
rect 28169 24695 28227 24701
rect 28184 24596 28212 24695
rect 30006 24692 30012 24744
rect 30064 24692 30070 24744
rect 37277 24735 37335 24741
rect 37277 24732 37289 24735
rect 36832 24704 37289 24732
rect 30024 24664 30052 24692
rect 29104 24636 30052 24664
rect 29104 24596 29132 24636
rect 36832 24608 36860 24704
rect 37277 24701 37289 24704
rect 37323 24701 37335 24735
rect 37277 24695 37335 24701
rect 28184 24568 29132 24596
rect 29454 24556 29460 24608
rect 29512 24596 29518 24608
rect 29549 24599 29607 24605
rect 29549 24596 29561 24599
rect 29512 24568 29561 24596
rect 29512 24556 29518 24568
rect 29549 24565 29561 24568
rect 29595 24565 29607 24599
rect 29549 24559 29607 24565
rect 35342 24556 35348 24608
rect 35400 24556 35406 24608
rect 36814 24556 36820 24608
rect 36872 24556 36878 24608
rect 36998 24556 37004 24608
rect 37056 24596 37062 24608
rect 37921 24599 37979 24605
rect 37921 24596 37933 24599
rect 37056 24568 37933 24596
rect 37056 24556 37062 24568
rect 37921 24565 37933 24568
rect 37967 24565 37979 24599
rect 37921 24559 37979 24565
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 28813 24395 28871 24401
rect 28813 24361 28825 24395
rect 28859 24392 28871 24395
rect 28902 24392 28908 24404
rect 28859 24364 28908 24392
rect 28859 24361 28871 24364
rect 28813 24355 28871 24361
rect 28902 24352 28908 24364
rect 28960 24352 28966 24404
rect 29546 24352 29552 24404
rect 29604 24392 29610 24404
rect 30285 24395 30343 24401
rect 30285 24392 30297 24395
rect 29604 24364 30297 24392
rect 29604 24352 29610 24364
rect 30285 24361 30297 24364
rect 30331 24361 30343 24395
rect 31202 24392 31208 24404
rect 30285 24355 30343 24361
rect 30576 24364 31208 24392
rect 30576 24336 30604 24364
rect 31202 24352 31208 24364
rect 31260 24392 31266 24404
rect 31570 24392 31576 24404
rect 31260 24364 31576 24392
rect 31260 24352 31266 24364
rect 31570 24352 31576 24364
rect 31628 24352 31634 24404
rect 33229 24395 33287 24401
rect 33229 24392 33241 24395
rect 31726 24364 33241 24392
rect 30558 24324 30564 24336
rect 29012 24296 30564 24324
rect 934 24148 940 24200
rect 992 24188 998 24200
rect 29012 24197 29040 24296
rect 30558 24284 30564 24296
rect 30616 24284 30622 24336
rect 31726 24324 31754 24364
rect 33229 24361 33241 24364
rect 33275 24361 33287 24395
rect 33229 24355 33287 24361
rect 35342 24352 35348 24404
rect 35400 24352 35406 24404
rect 36998 24352 37004 24404
rect 37056 24352 37062 24404
rect 31220 24296 31754 24324
rect 30653 24259 30711 24265
rect 30653 24256 30665 24259
rect 29564 24228 30665 24256
rect 29564 24200 29592 24228
rect 30653 24225 30665 24228
rect 30699 24225 30711 24259
rect 30653 24219 30711 24225
rect 31018 24216 31024 24268
rect 31076 24256 31082 24268
rect 31220 24265 31248 24296
rect 31205 24259 31263 24265
rect 31205 24256 31217 24259
rect 31076 24228 31217 24256
rect 31076 24216 31082 24228
rect 31205 24225 31217 24228
rect 31251 24225 31263 24259
rect 31205 24219 31263 24225
rect 31846 24216 31852 24268
rect 31904 24216 31910 24268
rect 35360 24265 35388 24352
rect 35526 24284 35532 24336
rect 35584 24324 35590 24336
rect 35989 24327 36047 24333
rect 35989 24324 36001 24327
rect 35584 24296 36001 24324
rect 35584 24284 35590 24296
rect 35989 24293 36001 24296
rect 36035 24293 36047 24327
rect 37016 24324 37044 24352
rect 35989 24287 36047 24293
rect 36096 24296 37044 24324
rect 35345 24259 35403 24265
rect 35345 24225 35357 24259
rect 35391 24256 35403 24259
rect 35894 24256 35900 24268
rect 35391 24228 35900 24256
rect 35391 24225 35403 24228
rect 35345 24219 35403 24225
rect 35894 24216 35900 24228
rect 35952 24216 35958 24268
rect 1581 24191 1639 24197
rect 1581 24188 1593 24191
rect 992 24160 1593 24188
rect 992 24148 998 24160
rect 1581 24157 1593 24160
rect 1627 24157 1639 24191
rect 1581 24151 1639 24157
rect 28997 24191 29055 24197
rect 28997 24157 29009 24191
rect 29043 24157 29055 24191
rect 28997 24151 29055 24157
rect 29089 24191 29147 24197
rect 29089 24157 29101 24191
rect 29135 24188 29147 24191
rect 29454 24188 29460 24200
rect 29135 24160 29460 24188
rect 29135 24157 29147 24160
rect 29089 24151 29147 24157
rect 29454 24148 29460 24160
rect 29512 24148 29518 24200
rect 29546 24148 29552 24200
rect 29604 24148 29610 24200
rect 30469 24191 30527 24197
rect 30469 24157 30481 24191
rect 30515 24157 30527 24191
rect 30469 24151 30527 24157
rect 28813 24123 28871 24129
rect 28813 24089 28825 24123
rect 28859 24120 28871 24123
rect 30193 24123 30251 24129
rect 30193 24120 30205 24123
rect 28859 24092 30205 24120
rect 28859 24089 28871 24092
rect 28813 24083 28871 24089
rect 30193 24089 30205 24092
rect 30239 24089 30251 24123
rect 30484 24120 30512 24151
rect 30558 24148 30564 24200
rect 30616 24148 30622 24200
rect 30745 24191 30803 24197
rect 30745 24157 30757 24191
rect 30791 24188 30803 24191
rect 31386 24188 31392 24200
rect 30791 24160 31392 24188
rect 30791 24157 30803 24160
rect 30745 24151 30803 24157
rect 31386 24148 31392 24160
rect 31444 24188 31450 24200
rect 31444 24182 31892 24188
rect 31956 24182 33824 24188
rect 31444 24160 33824 24182
rect 31444 24148 31450 24160
rect 31864 24154 31984 24160
rect 30484 24092 30604 24120
rect 30193 24083 30251 24089
rect 29914 24012 29920 24064
rect 29972 24052 29978 24064
rect 30576 24052 30604 24092
rect 31294 24080 31300 24132
rect 31352 24120 31358 24132
rect 32094 24123 32152 24129
rect 32094 24120 32106 24123
rect 31352 24092 32106 24120
rect 31352 24080 31358 24092
rect 32094 24089 32106 24092
rect 32140 24089 32152 24123
rect 32094 24083 32152 24089
rect 31478 24052 31484 24064
rect 29972 24024 31484 24052
rect 29972 24012 29978 24024
rect 31478 24012 31484 24024
rect 31536 24012 31542 24064
rect 31754 24012 31760 24064
rect 31812 24012 31818 24064
rect 33796 24052 33824 24160
rect 35912 24120 35940 24216
rect 36096 24197 36124 24296
rect 36262 24216 36268 24268
rect 36320 24256 36326 24268
rect 36357 24259 36415 24265
rect 36357 24256 36369 24259
rect 36320 24228 36369 24256
rect 36320 24216 36326 24228
rect 36357 24225 36369 24228
rect 36403 24225 36415 24259
rect 36357 24219 36415 24225
rect 36081 24191 36139 24197
rect 36081 24157 36093 24191
rect 36127 24157 36139 24191
rect 36081 24151 36139 24157
rect 36173 24191 36231 24197
rect 36173 24157 36185 24191
rect 36219 24188 36231 24191
rect 36538 24188 36544 24200
rect 36219 24160 36544 24188
rect 36219 24157 36231 24160
rect 36173 24151 36231 24157
rect 36538 24148 36544 24160
rect 36596 24148 36602 24200
rect 36722 24148 36728 24200
rect 36780 24148 36786 24200
rect 37369 24191 37427 24197
rect 37369 24157 37381 24191
rect 37415 24188 37427 24191
rect 37415 24160 37872 24188
rect 37415 24157 37427 24160
rect 37369 24151 37427 24157
rect 36446 24120 36452 24132
rect 35912 24092 36452 24120
rect 36446 24080 36452 24092
rect 36504 24080 36510 24132
rect 37636 24123 37694 24129
rect 37636 24089 37648 24123
rect 37682 24120 37694 24123
rect 37734 24120 37740 24132
rect 37682 24092 37740 24120
rect 37682 24089 37694 24092
rect 37636 24083 37694 24089
rect 37734 24080 37740 24092
rect 37792 24080 37798 24132
rect 37844 24064 37872 24160
rect 35894 24052 35900 24064
rect 33796 24024 35900 24052
rect 35894 24012 35900 24024
rect 35952 24012 35958 24064
rect 36354 24012 36360 24064
rect 36412 24012 36418 24064
rect 37277 24055 37335 24061
rect 37277 24021 37289 24055
rect 37323 24052 37335 24055
rect 37550 24052 37556 24064
rect 37323 24024 37556 24052
rect 37323 24021 37335 24024
rect 37277 24015 37335 24021
rect 37550 24012 37556 24024
rect 37608 24012 37614 24064
rect 37826 24012 37832 24064
rect 37884 24012 37890 24064
rect 38286 24012 38292 24064
rect 38344 24052 38350 24064
rect 38749 24055 38807 24061
rect 38749 24052 38761 24055
rect 38344 24024 38761 24052
rect 38344 24012 38350 24024
rect 38749 24021 38761 24024
rect 38795 24021 38807 24055
rect 38749 24015 38807 24021
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 30282 23808 30288 23860
rect 30340 23848 30346 23860
rect 30377 23851 30435 23857
rect 30377 23848 30389 23851
rect 30340 23820 30389 23848
rect 30340 23808 30346 23820
rect 30377 23817 30389 23820
rect 30423 23817 30435 23851
rect 32214 23848 32220 23860
rect 30377 23811 30435 23817
rect 31220 23820 32220 23848
rect 28353 23783 28411 23789
rect 28353 23749 28365 23783
rect 28399 23780 28411 23783
rect 28813 23783 28871 23789
rect 28813 23780 28825 23783
rect 28399 23752 28825 23780
rect 28399 23749 28411 23752
rect 28353 23743 28411 23749
rect 28813 23749 28825 23752
rect 28859 23749 28871 23783
rect 29086 23780 29092 23792
rect 28813 23743 28871 23749
rect 28920 23752 29092 23780
rect 27154 23672 27160 23724
rect 27212 23672 27218 23724
rect 28261 23715 28319 23721
rect 28261 23681 28273 23715
rect 28307 23681 28319 23715
rect 28261 23675 28319 23681
rect 28276 23576 28304 23675
rect 28442 23672 28448 23724
rect 28500 23672 28506 23724
rect 28583 23715 28641 23721
rect 28583 23681 28595 23715
rect 28629 23712 28641 23715
rect 28920 23712 28948 23752
rect 29086 23740 29092 23752
rect 29144 23740 29150 23792
rect 29546 23780 29552 23792
rect 29196 23752 29552 23780
rect 29196 23724 29224 23752
rect 29546 23740 29552 23752
rect 29604 23740 29610 23792
rect 31113 23783 31171 23789
rect 31113 23780 31125 23783
rect 30576 23752 31125 23780
rect 28629 23684 28948 23712
rect 28997 23715 29055 23721
rect 28629 23681 28641 23684
rect 28583 23675 28641 23681
rect 28997 23681 29009 23715
rect 29043 23681 29055 23715
rect 28997 23675 29055 23681
rect 28721 23647 28779 23653
rect 28721 23613 28733 23647
rect 28767 23644 28779 23647
rect 28902 23644 28908 23656
rect 28767 23616 28908 23644
rect 28767 23613 28779 23616
rect 28721 23607 28779 23613
rect 28902 23604 28908 23616
rect 28960 23644 28966 23656
rect 29012 23644 29040 23675
rect 29178 23672 29184 23724
rect 29236 23672 29242 23724
rect 29273 23715 29331 23721
rect 29273 23681 29285 23715
rect 29319 23712 29331 23715
rect 29365 23715 29423 23721
rect 29365 23712 29377 23715
rect 29319 23684 29377 23712
rect 29319 23681 29331 23684
rect 29273 23675 29331 23681
rect 29365 23681 29377 23684
rect 29411 23712 29423 23715
rect 29454 23712 29460 23724
rect 29411 23684 29460 23712
rect 29411 23681 29423 23684
rect 29365 23675 29423 23681
rect 29454 23672 29460 23684
rect 29512 23672 29518 23724
rect 30576 23721 30604 23752
rect 31113 23749 31125 23752
rect 31159 23749 31171 23783
rect 31113 23743 31171 23749
rect 31220 23721 31248 23820
rect 32214 23808 32220 23820
rect 32272 23808 32278 23860
rect 35342 23848 35348 23860
rect 34256 23820 35348 23848
rect 31294 23740 31300 23792
rect 31352 23740 31358 23792
rect 31570 23740 31576 23792
rect 31628 23780 31634 23792
rect 34256 23789 34284 23820
rect 35342 23808 35348 23820
rect 35400 23808 35406 23860
rect 35544 23820 36032 23848
rect 34241 23783 34299 23789
rect 31628 23752 32352 23780
rect 31628 23740 31634 23752
rect 29641 23715 29699 23721
rect 29641 23681 29653 23715
rect 29687 23681 29699 23715
rect 29641 23675 29699 23681
rect 30561 23715 30619 23721
rect 30561 23681 30573 23715
rect 30607 23681 30619 23715
rect 31021 23715 31079 23721
rect 31021 23712 31033 23715
rect 30561 23675 30619 23681
rect 30760 23684 31033 23712
rect 29656 23644 29684 23675
rect 28960 23616 29684 23644
rect 28960 23604 28966 23616
rect 29457 23579 29515 23585
rect 29457 23576 29469 23579
rect 28276 23548 29469 23576
rect 29457 23545 29469 23548
rect 29503 23545 29515 23579
rect 30760 23576 30788 23684
rect 31021 23681 31033 23684
rect 31067 23681 31079 23715
rect 31021 23675 31079 23681
rect 31205 23715 31263 23721
rect 31205 23681 31217 23715
rect 31251 23681 31263 23715
rect 31205 23675 31263 23681
rect 31481 23715 31539 23721
rect 31481 23681 31493 23715
rect 31527 23681 31539 23715
rect 31481 23675 31539 23681
rect 30837 23647 30895 23653
rect 30837 23613 30849 23647
rect 30883 23644 30895 23647
rect 30926 23644 30932 23656
rect 30883 23616 30932 23644
rect 30883 23613 30895 23616
rect 30837 23607 30895 23613
rect 30926 23604 30932 23616
rect 30984 23604 30990 23656
rect 31496 23576 31524 23675
rect 31754 23672 31760 23724
rect 31812 23672 31818 23724
rect 32214 23672 32220 23724
rect 32272 23672 32278 23724
rect 32324 23721 32352 23752
rect 34241 23749 34253 23783
rect 34287 23749 34299 23783
rect 34241 23743 34299 23749
rect 34457 23783 34515 23789
rect 34457 23749 34469 23783
rect 34503 23780 34515 23783
rect 34698 23780 34704 23792
rect 34503 23752 34704 23780
rect 34503 23749 34515 23752
rect 34457 23743 34515 23749
rect 34698 23740 34704 23752
rect 34756 23740 34762 23792
rect 35544 23780 35572 23820
rect 34808 23752 35572 23780
rect 32309 23715 32367 23721
rect 32309 23681 32321 23715
rect 32355 23681 32367 23715
rect 32309 23675 32367 23681
rect 32398 23672 32404 23724
rect 32456 23712 32462 23724
rect 32585 23715 32643 23721
rect 32585 23712 32597 23715
rect 32456 23684 32597 23712
rect 32456 23672 32462 23684
rect 32585 23681 32597 23684
rect 32631 23681 32643 23715
rect 32585 23675 32643 23681
rect 32769 23715 32827 23721
rect 32769 23681 32781 23715
rect 32815 23681 32827 23715
rect 32769 23675 32827 23681
rect 31938 23604 31944 23656
rect 31996 23644 32002 23656
rect 32125 23647 32183 23653
rect 32125 23644 32137 23647
rect 31996 23616 32137 23644
rect 31996 23604 32002 23616
rect 32125 23613 32137 23616
rect 32171 23613 32183 23647
rect 32232 23644 32260 23672
rect 32784 23644 32812 23675
rect 32950 23644 32956 23656
rect 32232 23616 32956 23644
rect 32125 23607 32183 23613
rect 32950 23604 32956 23616
rect 33008 23604 33014 23656
rect 34701 23647 34759 23653
rect 34701 23644 34713 23647
rect 34532 23616 34713 23644
rect 32585 23579 32643 23585
rect 32585 23576 32597 23579
rect 30760 23548 31432 23576
rect 31496 23548 32597 23576
rect 29457 23539 29515 23545
rect 26970 23468 26976 23520
rect 27028 23468 27034 23520
rect 28074 23468 28080 23520
rect 28132 23468 28138 23520
rect 30190 23468 30196 23520
rect 30248 23508 30254 23520
rect 30745 23511 30803 23517
rect 30745 23508 30757 23511
rect 30248 23480 30757 23508
rect 30248 23468 30254 23480
rect 30745 23477 30757 23480
rect 30791 23477 30803 23511
rect 31404 23508 31432 23548
rect 32585 23545 32597 23548
rect 32631 23545 32643 23579
rect 32585 23539 32643 23545
rect 34238 23536 34244 23588
rect 34296 23576 34302 23588
rect 34532 23576 34560 23616
rect 34701 23613 34713 23616
rect 34747 23613 34759 23647
rect 34701 23607 34759 23613
rect 34296 23548 34560 23576
rect 34609 23579 34667 23585
rect 34296 23536 34302 23548
rect 34609 23545 34621 23579
rect 34655 23576 34667 23579
rect 34808 23576 34836 23752
rect 35176 23721 35204 23752
rect 34885 23715 34943 23721
rect 34885 23681 34897 23715
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 35161 23715 35219 23721
rect 35161 23681 35173 23715
rect 35207 23681 35219 23715
rect 35161 23675 35219 23681
rect 35345 23715 35403 23721
rect 35345 23681 35357 23715
rect 35391 23712 35403 23715
rect 35526 23712 35532 23724
rect 35391 23684 35532 23712
rect 35391 23681 35403 23684
rect 35345 23675 35403 23681
rect 34900 23644 34928 23675
rect 35526 23672 35532 23684
rect 35584 23672 35590 23724
rect 35437 23647 35495 23653
rect 35437 23644 35449 23647
rect 34900 23616 35449 23644
rect 35437 23613 35449 23616
rect 35483 23613 35495 23647
rect 35437 23607 35495 23613
rect 35618 23604 35624 23656
rect 35676 23604 35682 23656
rect 35713 23647 35771 23653
rect 35713 23613 35725 23647
rect 35759 23613 35771 23647
rect 35713 23607 35771 23613
rect 34655 23548 34836 23576
rect 34655 23545 34667 23548
rect 34609 23539 34667 23545
rect 35342 23536 35348 23588
rect 35400 23576 35406 23588
rect 35728 23576 35756 23607
rect 35802 23604 35808 23656
rect 35860 23604 35866 23656
rect 35894 23604 35900 23656
rect 35952 23604 35958 23656
rect 36004 23644 36032 23820
rect 36078 23808 36084 23860
rect 36136 23848 36142 23860
rect 36173 23851 36231 23857
rect 36173 23848 36185 23851
rect 36136 23820 36185 23848
rect 36136 23808 36142 23820
rect 36173 23817 36185 23820
rect 36219 23817 36231 23851
rect 36173 23811 36231 23817
rect 36354 23808 36360 23860
rect 36412 23808 36418 23860
rect 36446 23808 36452 23860
rect 36504 23848 36510 23860
rect 36725 23851 36783 23857
rect 36725 23848 36737 23851
rect 36504 23820 36737 23848
rect 36504 23808 36510 23820
rect 36725 23817 36737 23820
rect 36771 23817 36783 23851
rect 36725 23811 36783 23817
rect 38028 23820 38608 23848
rect 36372 23780 36400 23808
rect 36096 23752 36400 23780
rect 36096 23721 36124 23752
rect 36538 23740 36544 23792
rect 36596 23780 36602 23792
rect 38028 23789 38056 23820
rect 38580 23792 38608 23820
rect 36909 23783 36967 23789
rect 36909 23780 36921 23783
rect 36596 23752 36921 23780
rect 36596 23740 36602 23752
rect 36909 23749 36921 23752
rect 36955 23749 36967 23783
rect 36909 23743 36967 23749
rect 38013 23783 38071 23789
rect 38013 23749 38025 23783
rect 38059 23749 38071 23783
rect 38013 23743 38071 23749
rect 38243 23749 38301 23755
rect 38243 23746 38255 23749
rect 36081 23715 36139 23721
rect 36081 23681 36093 23715
rect 36127 23681 36139 23715
rect 36081 23675 36139 23681
rect 36265 23715 36323 23721
rect 36265 23681 36277 23715
rect 36311 23681 36323 23715
rect 36265 23675 36323 23681
rect 36280 23644 36308 23675
rect 36814 23672 36820 23724
rect 36872 23672 36878 23724
rect 37182 23672 37188 23724
rect 37240 23712 37246 23724
rect 38228 23715 38255 23746
rect 38289 23715 38301 23749
rect 38562 23740 38568 23792
rect 38620 23740 38626 23792
rect 38228 23712 38301 23715
rect 37240 23709 38301 23712
rect 38832 23715 38890 23721
rect 37240 23684 38256 23709
rect 37240 23672 37246 23684
rect 38832 23681 38844 23715
rect 38878 23712 38890 23715
rect 39298 23712 39304 23724
rect 38878 23684 39304 23712
rect 38878 23681 38890 23684
rect 38832 23675 38890 23681
rect 39298 23672 39304 23684
rect 39356 23672 39362 23724
rect 45554 23672 45560 23724
rect 45612 23712 45618 23724
rect 46661 23715 46719 23721
rect 46661 23712 46673 23715
rect 45612 23684 46673 23712
rect 45612 23672 45618 23684
rect 46661 23681 46673 23684
rect 46707 23712 46719 23715
rect 46842 23712 46848 23724
rect 46707 23684 46848 23712
rect 46707 23681 46719 23684
rect 46661 23675 46719 23681
rect 46842 23672 46848 23684
rect 46900 23672 46906 23724
rect 36004 23616 36308 23644
rect 36541 23647 36599 23653
rect 36541 23613 36553 23647
rect 36587 23644 36599 23647
rect 37369 23647 37427 23653
rect 37369 23644 37381 23647
rect 36587 23616 37381 23644
rect 36587 23613 36599 23616
rect 36541 23607 36599 23613
rect 37369 23613 37381 23616
rect 37415 23613 37427 23647
rect 37369 23607 37427 23613
rect 36814 23576 36820 23588
rect 35400 23548 36820 23576
rect 35400 23536 35406 23548
rect 36814 23536 36820 23548
rect 36872 23536 36878 23588
rect 37384 23576 37412 23607
rect 37826 23604 37832 23656
rect 37884 23644 37890 23656
rect 38565 23647 38623 23653
rect 38565 23644 38577 23647
rect 37884 23616 38577 23644
rect 37884 23604 37890 23616
rect 38565 23613 38577 23616
rect 38611 23613 38623 23647
rect 38565 23607 38623 23613
rect 46017 23647 46075 23653
rect 46017 23613 46029 23647
rect 46063 23644 46075 23647
rect 47026 23644 47032 23656
rect 46063 23616 47032 23644
rect 46063 23613 46075 23616
rect 46017 23607 46075 23613
rect 47026 23604 47032 23616
rect 47084 23604 47090 23656
rect 38286 23576 38292 23588
rect 37384 23548 38292 23576
rect 31665 23511 31723 23517
rect 31665 23508 31677 23511
rect 31404 23480 31677 23508
rect 30745 23471 30803 23477
rect 31665 23477 31677 23480
rect 31711 23508 31723 23511
rect 32493 23511 32551 23517
rect 32493 23508 32505 23511
rect 31711 23480 32505 23508
rect 31711 23477 31723 23480
rect 31665 23471 31723 23477
rect 32493 23477 32505 23480
rect 32539 23477 32551 23511
rect 32493 23471 32551 23477
rect 34425 23511 34483 23517
rect 34425 23477 34437 23511
rect 34471 23508 34483 23511
rect 35434 23508 35440 23520
rect 34471 23480 35440 23508
rect 34471 23477 34483 23480
rect 34425 23471 34483 23477
rect 35434 23468 35440 23480
rect 35492 23468 35498 23520
rect 37093 23511 37151 23517
rect 37093 23477 37105 23511
rect 37139 23508 37151 23511
rect 37366 23508 37372 23520
rect 37139 23480 37372 23508
rect 37139 23477 37151 23480
rect 37093 23471 37151 23477
rect 37366 23468 37372 23480
rect 37424 23468 37430 23520
rect 37458 23468 37464 23520
rect 37516 23508 37522 23520
rect 38212 23517 38240 23548
rect 38286 23536 38292 23548
rect 38344 23536 38350 23588
rect 37921 23511 37979 23517
rect 37921 23508 37933 23511
rect 37516 23480 37933 23508
rect 37516 23468 37522 23480
rect 37921 23477 37933 23480
rect 37967 23477 37979 23511
rect 37921 23471 37979 23477
rect 38197 23511 38255 23517
rect 38197 23477 38209 23511
rect 38243 23477 38255 23511
rect 38197 23471 38255 23477
rect 38378 23468 38384 23520
rect 38436 23468 38442 23520
rect 38562 23468 38568 23520
rect 38620 23508 38626 23520
rect 39945 23511 40003 23517
rect 39945 23508 39957 23511
rect 38620 23480 39957 23508
rect 38620 23468 38626 23480
rect 39945 23477 39957 23480
rect 39991 23477 40003 23511
rect 39945 23471 40003 23477
rect 46106 23468 46112 23520
rect 46164 23508 46170 23520
rect 46569 23511 46627 23517
rect 46569 23508 46581 23511
rect 46164 23480 46581 23508
rect 46164 23468 46170 23480
rect 46569 23477 46581 23480
rect 46615 23477 46627 23511
rect 46569 23471 46627 23477
rect 46753 23511 46811 23517
rect 46753 23477 46765 23511
rect 46799 23508 46811 23511
rect 46934 23508 46940 23520
rect 46799 23480 46940 23508
rect 46799 23477 46811 23480
rect 46753 23471 46811 23477
rect 46934 23468 46940 23480
rect 46992 23468 46998 23520
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 28442 23264 28448 23316
rect 28500 23304 28506 23316
rect 29089 23307 29147 23313
rect 29089 23304 29101 23307
rect 28500 23276 29101 23304
rect 28500 23264 28506 23276
rect 29089 23273 29101 23276
rect 29135 23304 29147 23307
rect 30190 23304 30196 23316
rect 29135 23276 30196 23304
rect 29135 23273 29147 23276
rect 29089 23267 29147 23273
rect 30190 23264 30196 23276
rect 30248 23264 30254 23316
rect 31018 23264 31024 23316
rect 31076 23264 31082 23316
rect 32674 23304 32680 23316
rect 32048 23276 32680 23304
rect 32048 23245 32076 23276
rect 32674 23264 32680 23276
rect 32732 23264 32738 23316
rect 33042 23264 33048 23316
rect 33100 23304 33106 23316
rect 34514 23304 34520 23316
rect 33100 23276 34520 23304
rect 33100 23264 33106 23276
rect 34514 23264 34520 23276
rect 34572 23264 34578 23316
rect 34698 23264 34704 23316
rect 34756 23304 34762 23316
rect 35069 23307 35127 23313
rect 35069 23304 35081 23307
rect 34756 23276 35081 23304
rect 34756 23264 34762 23276
rect 35069 23273 35081 23276
rect 35115 23304 35127 23307
rect 35342 23304 35348 23316
rect 35115 23276 35348 23304
rect 35115 23273 35127 23276
rect 35069 23267 35127 23273
rect 35342 23264 35348 23276
rect 35400 23264 35406 23316
rect 36449 23307 36507 23313
rect 36449 23304 36461 23307
rect 35636 23276 36461 23304
rect 35636 23248 35664 23276
rect 36449 23273 36461 23276
rect 36495 23304 36507 23307
rect 36538 23304 36544 23316
rect 36495 23276 36544 23304
rect 36495 23273 36507 23276
rect 36449 23267 36507 23273
rect 36538 23264 36544 23276
rect 36596 23264 36602 23316
rect 36722 23264 36728 23316
rect 36780 23304 36786 23316
rect 37001 23307 37059 23313
rect 37001 23304 37013 23307
rect 36780 23276 37013 23304
rect 36780 23264 36786 23276
rect 37001 23273 37013 23276
rect 37047 23273 37059 23307
rect 37001 23267 37059 23273
rect 37090 23264 37096 23316
rect 37148 23304 37154 23316
rect 37277 23307 37335 23313
rect 37277 23304 37289 23307
rect 37148 23276 37289 23304
rect 37148 23264 37154 23276
rect 37277 23273 37289 23276
rect 37323 23273 37335 23307
rect 37277 23267 37335 23273
rect 37734 23264 37740 23316
rect 37792 23264 37798 23316
rect 38304 23276 38700 23304
rect 27985 23239 28043 23245
rect 27985 23205 27997 23239
rect 28031 23205 28043 23239
rect 31205 23239 31263 23245
rect 31205 23236 31217 23239
rect 27985 23199 28043 23205
rect 28736 23208 31217 23236
rect 26602 23060 26608 23112
rect 26660 23060 26666 23112
rect 28000 23100 28028 23199
rect 28736 23177 28764 23208
rect 31205 23205 31217 23208
rect 31251 23205 31263 23239
rect 31205 23199 31263 23205
rect 32033 23239 32091 23245
rect 32033 23205 32045 23239
rect 32079 23205 32091 23239
rect 35618 23236 35624 23248
rect 32033 23199 32091 23205
rect 34348 23208 35624 23236
rect 28721 23171 28779 23177
rect 28721 23137 28733 23171
rect 28767 23137 28779 23171
rect 28721 23131 28779 23137
rect 28813 23171 28871 23177
rect 28813 23137 28825 23171
rect 28859 23168 28871 23171
rect 29178 23168 29184 23180
rect 28859 23140 29184 23168
rect 28859 23137 28871 23140
rect 28813 23131 28871 23137
rect 29178 23128 29184 23140
rect 29236 23128 29242 23180
rect 29454 23128 29460 23180
rect 29512 23168 29518 23180
rect 29914 23168 29920 23180
rect 29512 23140 29920 23168
rect 29512 23128 29518 23140
rect 28902 23102 28908 23112
rect 28736 23100 28908 23102
rect 28000 23074 28908 23100
rect 28000 23072 28764 23074
rect 28902 23060 28908 23074
rect 28960 23060 28966 23112
rect 29086 23060 29092 23112
rect 29144 23060 29150 23112
rect 29564 23109 29592 23140
rect 29914 23128 29920 23140
rect 29972 23128 29978 23180
rect 31110 23168 31116 23180
rect 30944 23140 31116 23168
rect 30944 23109 30972 23140
rect 31110 23128 31116 23140
rect 31168 23168 31174 23180
rect 31168 23140 31616 23168
rect 31168 23128 31174 23140
rect 29273 23103 29331 23109
rect 29273 23069 29285 23103
rect 29319 23069 29331 23103
rect 29273 23063 29331 23069
rect 29549 23103 29607 23109
rect 29549 23069 29561 23103
rect 29595 23069 29607 23103
rect 29549 23063 29607 23069
rect 29641 23103 29699 23109
rect 29641 23069 29653 23103
rect 29687 23100 29699 23103
rect 29825 23103 29883 23109
rect 29825 23100 29837 23103
rect 29687 23072 29837 23100
rect 29687 23069 29699 23072
rect 29641 23063 29699 23069
rect 29825 23069 29837 23072
rect 29871 23069 29883 23103
rect 30193 23103 30251 23109
rect 30193 23100 30205 23103
rect 29825 23063 29883 23069
rect 29932 23072 30205 23100
rect 26872 23035 26930 23041
rect 26872 23001 26884 23035
rect 26918 23032 26930 23035
rect 26970 23032 26976 23044
rect 26918 23004 26976 23032
rect 26918 23001 26930 23004
rect 26872 22995 26930 23001
rect 26970 22992 26976 23004
rect 27028 22992 27034 23044
rect 29288 23032 29316 23063
rect 28966 23004 29316 23032
rect 28534 22924 28540 22976
rect 28592 22964 28598 22976
rect 28966 22964 28994 23004
rect 28592 22936 28994 22964
rect 28592 22924 28598 22936
rect 29270 22924 29276 22976
rect 29328 22964 29334 22976
rect 29932 22964 29960 23072
rect 30193 23069 30205 23072
rect 30239 23069 30251 23103
rect 30193 23063 30251 23069
rect 30929 23103 30987 23109
rect 30929 23069 30941 23103
rect 30975 23069 30987 23103
rect 30929 23063 30987 23069
rect 31021 23103 31079 23109
rect 31021 23069 31033 23103
rect 31067 23100 31079 23103
rect 31481 23103 31539 23109
rect 31481 23100 31493 23103
rect 31067 23072 31493 23100
rect 31067 23069 31079 23072
rect 31021 23063 31079 23069
rect 31481 23069 31493 23072
rect 31527 23069 31539 23103
rect 31481 23063 31539 23069
rect 31588 23094 31616 23140
rect 31846 23128 31852 23180
rect 31904 23128 31910 23180
rect 32401 23171 32459 23177
rect 32401 23137 32413 23171
rect 32447 23138 32459 23171
rect 32447 23137 32536 23138
rect 32401 23131 32536 23137
rect 32416 23112 32536 23131
rect 31662 23094 31668 23112
rect 31588 23066 31668 23094
rect 30009 23035 30067 23041
rect 30009 23001 30021 23035
rect 30055 23001 30067 23035
rect 30009 22995 30067 23001
rect 30101 23035 30159 23041
rect 30101 23001 30113 23035
rect 30147 23032 30159 23035
rect 30561 23035 30619 23041
rect 30561 23032 30573 23035
rect 30147 23004 30573 23032
rect 30147 23001 30159 23004
rect 30101 22995 30159 23001
rect 30561 23001 30573 23004
rect 30607 23032 30619 23035
rect 31294 23032 31300 23044
rect 30607 23004 31300 23032
rect 30607 23001 30619 23004
rect 30561 22995 30619 23001
rect 29328 22936 29960 22964
rect 30024 22964 30052 22995
rect 31294 22992 31300 23004
rect 31352 22992 31358 23044
rect 31496 23032 31524 23063
rect 31662 23060 31668 23066
rect 31720 23060 31726 23112
rect 32306 23060 32312 23112
rect 32364 23060 32370 23112
rect 32416 23110 32496 23112
rect 32490 23060 32496 23110
rect 32548 23060 32554 23112
rect 34348 23109 34376 23208
rect 35618 23196 35624 23208
rect 35676 23196 35682 23248
rect 36096 23208 37228 23236
rect 36096 23177 36124 23208
rect 37200 23180 37228 23208
rect 37550 23196 37556 23248
rect 37608 23236 37614 23248
rect 38304 23245 38332 23276
rect 37829 23239 37887 23245
rect 37829 23236 37841 23239
rect 37608 23208 37841 23236
rect 37608 23196 37614 23208
rect 37829 23205 37841 23208
rect 37875 23205 37887 23239
rect 38289 23239 38347 23245
rect 38289 23236 38301 23239
rect 37829 23199 37887 23205
rect 37936 23208 38301 23236
rect 34425 23171 34483 23177
rect 34425 23137 34437 23171
rect 34471 23168 34483 23171
rect 35161 23171 35219 23177
rect 34471 23140 34928 23168
rect 34471 23137 34483 23140
rect 34425 23131 34483 23137
rect 34333 23103 34391 23109
rect 34333 23069 34345 23103
rect 34379 23069 34391 23103
rect 34333 23063 34391 23069
rect 34514 23060 34520 23112
rect 34572 23060 34578 23112
rect 34900 23109 34928 23140
rect 35161 23137 35173 23171
rect 35207 23168 35219 23171
rect 35989 23171 36047 23177
rect 35989 23168 36001 23171
rect 35207 23140 36001 23168
rect 35207 23137 35219 23140
rect 35161 23131 35219 23137
rect 35989 23137 36001 23140
rect 36035 23137 36047 23171
rect 35989 23131 36047 23137
rect 36081 23171 36139 23177
rect 36081 23137 36093 23171
rect 36127 23137 36139 23171
rect 36081 23131 36139 23137
rect 34885 23103 34943 23109
rect 34885 23069 34897 23103
rect 34931 23069 34943 23103
rect 34885 23063 34943 23069
rect 35434 23060 35440 23112
rect 35492 23100 35498 23112
rect 36096 23100 36124 23131
rect 36446 23128 36452 23180
rect 36504 23168 36510 23180
rect 36817 23171 36875 23177
rect 36817 23168 36829 23171
rect 36504 23140 36829 23168
rect 36504 23128 36510 23140
rect 36817 23137 36829 23140
rect 36863 23137 36875 23171
rect 36817 23131 36875 23137
rect 35492 23072 36124 23100
rect 36265 23097 36323 23103
rect 35492 23060 35498 23072
rect 36265 23063 36277 23097
rect 36311 23063 36323 23097
rect 36265 23057 36323 23063
rect 36538 23060 36544 23112
rect 36596 23100 36602 23112
rect 36633 23103 36691 23109
rect 36633 23100 36645 23103
rect 36596 23072 36645 23100
rect 36596 23060 36602 23072
rect 36633 23069 36645 23072
rect 36679 23069 36691 23103
rect 36633 23063 36691 23069
rect 31496 23004 31754 23032
rect 30190 22964 30196 22976
rect 30024 22936 30196 22964
rect 29328 22924 29334 22936
rect 30190 22924 30196 22936
rect 30248 22924 30254 22976
rect 30374 22924 30380 22976
rect 30432 22924 30438 22976
rect 31018 22924 31024 22976
rect 31076 22964 31082 22976
rect 31478 22964 31484 22976
rect 31076 22936 31484 22964
rect 31076 22924 31082 22936
rect 31478 22924 31484 22936
rect 31536 22964 31542 22976
rect 31573 22967 31631 22973
rect 31573 22964 31585 22967
rect 31536 22936 31585 22964
rect 31536 22924 31542 22936
rect 31573 22933 31585 22936
rect 31619 22933 31631 22967
rect 31726 22964 31754 23004
rect 32030 22992 32036 23044
rect 32088 22992 32094 23044
rect 32122 22992 32128 23044
rect 32180 23032 32186 23044
rect 32674 23041 32680 23044
rect 32217 23035 32275 23041
rect 32217 23032 32229 23035
rect 32180 23004 32229 23032
rect 32180 22992 32186 23004
rect 32217 23001 32229 23004
rect 32263 23001 32275 23035
rect 32217 22995 32275 23001
rect 32668 22995 32680 23041
rect 32732 23032 32738 23044
rect 32732 23004 32768 23032
rect 32674 22992 32680 22995
rect 32732 22992 32738 23004
rect 32490 22964 32496 22976
rect 31726 22936 32496 22964
rect 31573 22927 31631 22933
rect 32490 22924 32496 22936
rect 32548 22964 32554 22976
rect 33781 22967 33839 22973
rect 33781 22964 33793 22967
rect 32548 22936 33793 22964
rect 32548 22924 32554 22936
rect 33781 22933 33793 22936
rect 33827 22933 33839 22967
rect 33781 22927 33839 22933
rect 34701 22967 34759 22973
rect 34701 22933 34713 22967
rect 34747 22964 34759 22967
rect 34790 22964 34796 22976
rect 34747 22936 34796 22964
rect 34747 22933 34759 22936
rect 34701 22927 34759 22933
rect 34790 22924 34796 22936
rect 34848 22924 34854 22976
rect 35342 22924 35348 22976
rect 35400 22964 35406 22976
rect 36280 22964 36308 23057
rect 36832 23032 36860 23131
rect 37182 23128 37188 23180
rect 37240 23128 37246 23180
rect 37366 23128 37372 23180
rect 37424 23168 37430 23180
rect 37936 23168 37964 23208
rect 38289 23205 38301 23208
rect 38335 23205 38347 23239
rect 38289 23199 38347 23205
rect 38378 23196 38384 23248
rect 38436 23196 38442 23248
rect 38396 23168 38424 23196
rect 37424 23140 37964 23168
rect 38028 23140 38424 23168
rect 38473 23171 38531 23177
rect 37424 23128 37430 23140
rect 37001 23103 37059 23109
rect 37001 23069 37013 23103
rect 37047 23100 37059 23103
rect 37458 23100 37464 23112
rect 37047 23072 37464 23100
rect 37047 23069 37059 23072
rect 37001 23063 37059 23069
rect 37458 23060 37464 23072
rect 37516 23060 37522 23112
rect 37752 23109 37780 23140
rect 37737 23103 37795 23109
rect 37737 23069 37749 23103
rect 37783 23069 37795 23103
rect 38028 23100 38056 23140
rect 38473 23137 38485 23171
rect 38519 23137 38531 23171
rect 38473 23131 38531 23137
rect 37737 23063 37795 23069
rect 37844 23072 38056 23100
rect 38197 23103 38255 23109
rect 37093 23035 37151 23041
rect 37093 23032 37105 23035
rect 36832 23004 37105 23032
rect 37093 23001 37105 23004
rect 37139 23001 37151 23035
rect 37093 22995 37151 23001
rect 37309 23035 37367 23041
rect 37309 23001 37321 23035
rect 37355 23032 37367 23035
rect 37844 23032 37872 23072
rect 38197 23069 38209 23103
rect 38243 23069 38255 23103
rect 38488 23100 38516 23131
rect 38562 23128 38568 23180
rect 38620 23128 38626 23180
rect 38197 23063 38255 23069
rect 38304 23072 38516 23100
rect 38672 23100 38700 23276
rect 39298 23264 39304 23316
rect 39356 23264 39362 23316
rect 46860 23276 49188 23304
rect 46860 23248 46888 23276
rect 46842 23196 46848 23248
rect 46900 23196 46906 23248
rect 45557 23171 45615 23177
rect 45557 23137 45569 23171
rect 45603 23168 45615 23171
rect 47673 23171 47731 23177
rect 47673 23168 47685 23171
rect 45603 23140 47685 23168
rect 45603 23137 45615 23140
rect 45557 23131 45615 23137
rect 47673 23137 47685 23140
rect 47719 23168 47731 23171
rect 48038 23168 48044 23180
rect 47719 23140 48044 23168
rect 47719 23137 47731 23140
rect 47673 23131 47731 23137
rect 48038 23128 48044 23140
rect 48096 23128 48102 23180
rect 39577 23103 39635 23109
rect 39577 23100 39589 23103
rect 38672 23072 39589 23100
rect 37355 23004 37872 23032
rect 37355 23001 37367 23004
rect 37309 22995 37367 23001
rect 38010 22992 38016 23044
rect 38068 22992 38074 23044
rect 35400 22936 36308 22964
rect 36725 22967 36783 22973
rect 35400 22924 35406 22936
rect 36725 22933 36737 22967
rect 36771 22964 36783 22967
rect 36814 22964 36820 22976
rect 36771 22936 36820 22964
rect 36771 22933 36783 22936
rect 36725 22927 36783 22933
rect 36814 22924 36820 22936
rect 36872 22924 36878 22976
rect 37461 22967 37519 22973
rect 37461 22933 37473 22967
rect 37507 22964 37519 22967
rect 37734 22964 37740 22976
rect 37507 22936 37740 22964
rect 37507 22933 37519 22936
rect 37461 22927 37519 22933
rect 37734 22924 37740 22936
rect 37792 22924 37798 22976
rect 38212 22964 38240 23063
rect 38304 23044 38332 23072
rect 39577 23069 39589 23072
rect 39623 23069 39635 23103
rect 45005 23103 45063 23109
rect 45005 23100 45017 23103
rect 39577 23063 39635 23069
rect 44468 23072 45017 23100
rect 38286 22992 38292 23044
rect 38344 22992 38350 23044
rect 38473 23035 38531 23041
rect 38473 23001 38485 23035
rect 38519 23032 38531 23035
rect 39301 23035 39359 23041
rect 39301 23032 39313 23035
rect 38519 23004 39313 23032
rect 38519 23001 38531 23004
rect 38473 22995 38531 23001
rect 39301 23001 39313 23004
rect 39347 23001 39359 23035
rect 39301 22995 39359 23001
rect 44468 22976 44496 23072
rect 45005 23069 45017 23072
rect 45051 23100 45063 23103
rect 45462 23100 45468 23112
rect 45051 23072 45468 23100
rect 45051 23069 45063 23072
rect 45005 23063 45063 23069
rect 45462 23060 45468 23072
rect 45520 23060 45526 23112
rect 46934 23060 46940 23112
rect 46992 23060 46998 23112
rect 49160 23100 49188 23276
rect 49510 23100 49516 23112
rect 49160 23072 49516 23100
rect 49510 23060 49516 23072
rect 49568 23060 49574 23112
rect 45833 23035 45891 23041
rect 45833 23001 45845 23035
rect 45879 23032 45891 23035
rect 46106 23032 46112 23044
rect 45879 23004 46112 23032
rect 45879 23001 45891 23004
rect 45833 22995 45891 23001
rect 46106 22992 46112 23004
rect 46164 22992 46170 23044
rect 47946 22992 47952 23044
rect 48004 22992 48010 23044
rect 49605 23035 49663 23041
rect 49605 23032 49617 23035
rect 49174 23004 49617 23032
rect 49605 23001 49617 23004
rect 49651 23001 49663 23035
rect 49605 22995 49663 23001
rect 39209 22967 39267 22973
rect 39209 22964 39221 22967
rect 38212 22936 39221 22964
rect 39209 22933 39221 22936
rect 39255 22964 39267 22967
rect 39485 22967 39543 22973
rect 39485 22964 39497 22967
rect 39255 22936 39497 22964
rect 39255 22933 39267 22936
rect 39209 22927 39267 22933
rect 39485 22933 39497 22936
rect 39531 22933 39543 22967
rect 39485 22927 39543 22933
rect 44450 22924 44456 22976
rect 44508 22924 44514 22976
rect 45094 22924 45100 22976
rect 45152 22924 45158 22976
rect 47305 22967 47363 22973
rect 47305 22933 47317 22967
rect 47351 22964 47363 22967
rect 47578 22964 47584 22976
rect 47351 22936 47584 22964
rect 47351 22933 47363 22936
rect 47305 22927 47363 22933
rect 47578 22924 47584 22936
rect 47636 22924 47642 22976
rect 49418 22924 49424 22976
rect 49476 22924 49482 22976
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 27154 22720 27160 22772
rect 27212 22760 27218 22772
rect 27341 22763 27399 22769
rect 27341 22760 27353 22763
rect 27212 22732 27353 22760
rect 27212 22720 27218 22732
rect 27341 22729 27353 22732
rect 27387 22729 27399 22763
rect 27341 22723 27399 22729
rect 28074 22720 28080 22772
rect 28132 22720 28138 22772
rect 30282 22720 30288 22772
rect 30340 22760 30346 22772
rect 31202 22760 31208 22772
rect 30340 22732 31208 22760
rect 30340 22720 30346 22732
rect 31202 22720 31208 22732
rect 31260 22760 31266 22772
rect 31681 22763 31739 22769
rect 31681 22760 31693 22763
rect 31260 22732 31693 22760
rect 31260 22720 31266 22732
rect 31681 22729 31693 22732
rect 31727 22729 31739 22763
rect 31681 22723 31739 22729
rect 32122 22720 32128 22772
rect 32180 22760 32186 22772
rect 32953 22763 33011 22769
rect 32953 22760 32965 22763
rect 32180 22732 32965 22760
rect 32180 22720 32186 22732
rect 32953 22729 32965 22732
rect 32999 22729 33011 22763
rect 32953 22723 33011 22729
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22624 27215 22627
rect 28092 22624 28120 22720
rect 31478 22692 31484 22704
rect 31036 22664 31484 22692
rect 27203 22596 28120 22624
rect 30285 22627 30343 22633
rect 27203 22593 27215 22596
rect 27157 22587 27215 22593
rect 30285 22593 30297 22627
rect 30331 22624 30343 22627
rect 30834 22624 30840 22636
rect 30331 22596 30840 22624
rect 30331 22593 30343 22596
rect 30285 22587 30343 22593
rect 30834 22584 30840 22596
rect 30892 22584 30898 22636
rect 31036 22633 31064 22664
rect 31478 22652 31484 22664
rect 31536 22652 31542 22704
rect 32490 22652 32496 22704
rect 32548 22652 32554 22704
rect 31021 22627 31079 22633
rect 31021 22593 31033 22627
rect 31067 22593 31079 22627
rect 31021 22587 31079 22593
rect 31113 22627 31171 22633
rect 31113 22593 31125 22627
rect 31159 22624 31171 22627
rect 32401 22627 32459 22633
rect 32401 22624 32413 22627
rect 31159 22596 32413 22624
rect 31159 22593 31171 22596
rect 31113 22587 31171 22593
rect 32401 22593 32413 22596
rect 32447 22624 32459 22627
rect 32508 22624 32536 22652
rect 32447 22596 32536 22624
rect 32968 22624 32996 22723
rect 34790 22720 34796 22772
rect 34848 22720 34854 22772
rect 35434 22720 35440 22772
rect 35492 22720 35498 22772
rect 35618 22720 35624 22772
rect 35676 22760 35682 22772
rect 36262 22760 36268 22772
rect 35676 22732 36268 22760
rect 35676 22720 35682 22732
rect 36262 22720 36268 22732
rect 36320 22760 36326 22772
rect 38286 22760 38292 22772
rect 36320 22732 38292 22760
rect 36320 22720 36326 22732
rect 38286 22720 38292 22732
rect 38344 22720 38350 22772
rect 45002 22720 45008 22772
rect 45060 22760 45066 22772
rect 46017 22763 46075 22769
rect 46017 22760 46029 22763
rect 45060 22732 46029 22760
rect 45060 22720 45066 22732
rect 46017 22729 46029 22732
rect 46063 22729 46075 22763
rect 46017 22723 46075 22729
rect 46385 22763 46443 22769
rect 46385 22729 46397 22763
rect 46431 22760 46443 22763
rect 47118 22760 47124 22772
rect 46431 22732 47124 22760
rect 46431 22729 46443 22732
rect 46385 22723 46443 22729
rect 47118 22720 47124 22732
rect 47176 22720 47182 22772
rect 33045 22627 33103 22633
rect 33045 22624 33057 22627
rect 32968 22596 33057 22624
rect 32447 22593 32459 22596
rect 32401 22587 32459 22593
rect 33045 22593 33057 22596
rect 33091 22593 33103 22627
rect 33045 22587 33103 22593
rect 34054 22584 34060 22636
rect 34112 22584 34118 22636
rect 34324 22627 34382 22633
rect 34324 22593 34336 22627
rect 34370 22624 34382 22627
rect 34808 22624 34836 22720
rect 37366 22652 37372 22704
rect 37424 22692 37430 22704
rect 38010 22692 38016 22704
rect 37424 22664 38016 22692
rect 37424 22652 37430 22664
rect 38010 22652 38016 22664
rect 38068 22692 38074 22704
rect 38841 22695 38899 22701
rect 38841 22692 38853 22695
rect 38068 22664 38853 22692
rect 38068 22652 38074 22664
rect 38841 22661 38853 22664
rect 38887 22692 38899 22695
rect 44082 22692 44088 22704
rect 38887 22664 44088 22692
rect 38887 22661 38899 22664
rect 38841 22655 38899 22661
rect 44082 22652 44088 22664
rect 44140 22652 44146 22704
rect 45094 22652 45100 22704
rect 45152 22652 45158 22704
rect 46477 22695 46535 22701
rect 46477 22661 46489 22695
rect 46523 22692 46535 22695
rect 47302 22692 47308 22704
rect 46523 22664 47308 22692
rect 46523 22661 46535 22664
rect 46477 22655 46535 22661
rect 47302 22652 47308 22664
rect 47360 22652 47366 22704
rect 34370 22596 34836 22624
rect 38473 22627 38531 22633
rect 34370 22593 34382 22596
rect 34324 22587 34382 22593
rect 38473 22593 38485 22627
rect 38519 22624 38531 22627
rect 38565 22627 38623 22633
rect 38565 22624 38577 22627
rect 38519 22596 38577 22624
rect 38519 22593 38531 22596
rect 38473 22587 38531 22593
rect 38565 22593 38577 22596
rect 38611 22593 38623 22627
rect 46566 22624 46572 22636
rect 38565 22587 38623 22593
rect 45848 22596 46572 22624
rect 26694 22516 26700 22568
rect 26752 22556 26758 22568
rect 26973 22559 27031 22565
rect 26973 22556 26985 22559
rect 26752 22528 26985 22556
rect 26752 22516 26758 22528
rect 26973 22525 26985 22528
rect 27019 22525 27031 22559
rect 26973 22519 27031 22525
rect 30929 22559 30987 22565
rect 30929 22525 30941 22559
rect 30975 22525 30987 22559
rect 30929 22519 30987 22525
rect 31205 22559 31263 22565
rect 31205 22525 31217 22559
rect 31251 22556 31263 22559
rect 31294 22556 31300 22568
rect 31251 22528 31300 22556
rect 31251 22525 31263 22528
rect 31205 22519 31263 22525
rect 30944 22488 30972 22519
rect 31294 22516 31300 22528
rect 31352 22556 31358 22568
rect 31570 22556 31576 22568
rect 31352 22528 31576 22556
rect 31352 22516 31358 22528
rect 31570 22516 31576 22528
rect 31628 22516 31634 22568
rect 31662 22516 31668 22568
rect 31720 22516 31726 22568
rect 32030 22516 32036 22568
rect 32088 22516 32094 22568
rect 33318 22516 33324 22568
rect 33376 22516 33382 22568
rect 37458 22516 37464 22568
rect 37516 22556 37522 22568
rect 37829 22559 37887 22565
rect 37829 22556 37841 22559
rect 37516 22528 37841 22556
rect 37516 22516 37522 22528
rect 37829 22525 37841 22528
rect 37875 22525 37887 22559
rect 37829 22519 37887 22525
rect 43622 22516 43628 22568
rect 43680 22556 43686 22568
rect 44085 22559 44143 22565
rect 44085 22556 44097 22559
rect 43680 22528 44097 22556
rect 43680 22516 43686 22528
rect 44085 22525 44097 22528
rect 44131 22525 44143 22559
rect 44085 22519 44143 22525
rect 44358 22516 44364 22568
rect 44416 22516 44422 22568
rect 31680 22488 31708 22516
rect 30944 22460 31708 22488
rect 32048 22488 32076 22516
rect 33229 22491 33287 22497
rect 33229 22488 33241 22491
rect 32048 22460 33241 22488
rect 30101 22423 30159 22429
rect 30101 22389 30113 22423
rect 30147 22420 30159 22423
rect 30466 22420 30472 22432
rect 30147 22392 30472 22420
rect 30147 22389 30159 22392
rect 30101 22383 30159 22389
rect 30466 22380 30472 22392
rect 30524 22380 30530 22432
rect 30742 22380 30748 22432
rect 30800 22380 30806 22432
rect 31680 22429 31708 22460
rect 33229 22457 33241 22460
rect 33275 22457 33287 22491
rect 33229 22451 33287 22457
rect 38657 22491 38715 22497
rect 38657 22457 38669 22491
rect 38703 22488 38715 22491
rect 39022 22488 39028 22500
rect 38703 22460 39028 22488
rect 38703 22457 38715 22460
rect 38657 22451 38715 22457
rect 39022 22448 39028 22460
rect 39080 22448 39086 22500
rect 45848 22497 45876 22596
rect 46566 22584 46572 22596
rect 46624 22624 46630 22636
rect 46624 22596 46704 22624
rect 46624 22584 46630 22596
rect 46676 22565 46704 22596
rect 46842 22584 46848 22636
rect 46900 22584 46906 22636
rect 47029 22627 47087 22633
rect 47029 22593 47041 22627
rect 47075 22593 47087 22627
rect 47029 22587 47087 22593
rect 46661 22559 46719 22565
rect 46661 22525 46673 22559
rect 46707 22525 46719 22559
rect 47044 22556 47072 22587
rect 48866 22584 48872 22636
rect 48924 22624 48930 22636
rect 49418 22624 49424 22636
rect 48924 22596 49424 22624
rect 48924 22584 48930 22596
rect 49418 22584 49424 22596
rect 49476 22584 49482 22636
rect 47578 22556 47584 22568
rect 47044 22528 47584 22556
rect 46661 22519 46719 22525
rect 47578 22516 47584 22528
rect 47636 22516 47642 22568
rect 45833 22491 45891 22497
rect 45833 22457 45845 22491
rect 45879 22457 45891 22491
rect 45833 22451 45891 22457
rect 68462 22448 68468 22500
rect 68520 22448 68526 22500
rect 31665 22423 31723 22429
rect 31665 22389 31677 22423
rect 31711 22389 31723 22423
rect 31665 22383 31723 22389
rect 31849 22423 31907 22429
rect 31849 22389 31861 22423
rect 31895 22420 31907 22423
rect 32398 22420 32404 22432
rect 31895 22392 32404 22420
rect 31895 22389 31907 22392
rect 31849 22383 31907 22389
rect 32398 22380 32404 22392
rect 32456 22420 32462 22432
rect 33137 22423 33195 22429
rect 33137 22420 33149 22423
rect 32456 22392 33149 22420
rect 32456 22380 32462 22392
rect 33137 22389 33149 22392
rect 33183 22389 33195 22423
rect 33137 22383 33195 22389
rect 38746 22380 38752 22432
rect 38804 22380 38810 22432
rect 46658 22380 46664 22432
rect 46716 22420 46722 22432
rect 46845 22423 46903 22429
rect 46845 22420 46857 22423
rect 46716 22392 46857 22420
rect 46716 22380 46722 22392
rect 46845 22389 46857 22392
rect 46891 22389 46903 22423
rect 46845 22383 46903 22389
rect 47394 22380 47400 22432
rect 47452 22420 47458 22432
rect 48225 22423 48283 22429
rect 48225 22420 48237 22423
rect 47452 22392 48237 22420
rect 47452 22380 47458 22392
rect 48225 22389 48237 22392
rect 48271 22389 48283 22423
rect 48225 22383 48283 22389
rect 48314 22380 48320 22432
rect 48372 22420 48378 22432
rect 49421 22423 49479 22429
rect 49421 22420 49433 22423
rect 48372 22392 49433 22420
rect 48372 22380 48378 22392
rect 49421 22389 49433 22392
rect 49467 22389 49479 22423
rect 49421 22383 49479 22389
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 28905 22219 28963 22225
rect 28905 22185 28917 22219
rect 28951 22185 28963 22219
rect 28905 22179 28963 22185
rect 28920 22094 28948 22179
rect 29086 22176 29092 22228
rect 29144 22216 29150 22228
rect 29181 22219 29239 22225
rect 29181 22216 29193 22219
rect 29144 22188 29193 22216
rect 29144 22176 29150 22188
rect 29181 22185 29193 22188
rect 29227 22185 29239 22219
rect 29181 22179 29239 22185
rect 31570 22176 31576 22228
rect 31628 22176 31634 22228
rect 37458 22176 37464 22228
rect 37516 22176 37522 22228
rect 44358 22176 44364 22228
rect 44416 22216 44422 22228
rect 44637 22219 44695 22225
rect 44637 22216 44649 22219
rect 44416 22188 44649 22216
rect 44416 22176 44422 22188
rect 44637 22185 44649 22188
rect 44683 22185 44695 22219
rect 44637 22179 44695 22185
rect 47302 22176 47308 22228
rect 47360 22176 47366 22228
rect 47857 22219 47915 22225
rect 47857 22185 47869 22219
rect 47903 22216 47915 22219
rect 47946 22216 47952 22228
rect 47903 22188 47952 22216
rect 47903 22185 47915 22188
rect 47857 22179 47915 22185
rect 47946 22176 47952 22188
rect 48004 22176 48010 22228
rect 48130 22176 48136 22228
rect 48188 22216 48194 22228
rect 48593 22219 48651 22225
rect 48188 22188 48544 22216
rect 48188 22176 48194 22188
rect 29825 22151 29883 22157
rect 29825 22117 29837 22151
rect 29871 22117 29883 22151
rect 29825 22111 29883 22117
rect 28920 22080 28994 22094
rect 29086 22080 29092 22092
rect 28920 22066 29092 22080
rect 28966 22052 29092 22066
rect 29086 22040 29092 22052
rect 29144 22080 29150 22092
rect 29549 22083 29607 22089
rect 29549 22080 29561 22083
rect 29144 22052 29561 22080
rect 29144 22040 29150 22052
rect 29549 22049 29561 22052
rect 29595 22049 29607 22083
rect 29549 22043 29607 22049
rect 27341 22015 27399 22021
rect 27341 21981 27353 22015
rect 27387 22012 27399 22015
rect 28074 22012 28080 22024
rect 27387 21984 28080 22012
rect 27387 21981 27399 21984
rect 27341 21975 27399 21981
rect 28074 21972 28080 21984
rect 28132 21972 28138 22024
rect 28721 22015 28779 22021
rect 28721 21981 28733 22015
rect 28767 22012 28779 22015
rect 29840 22012 29868 22111
rect 33226 22108 33232 22160
rect 33284 22148 33290 22160
rect 33284 22120 34008 22148
rect 33284 22108 33290 22120
rect 33980 22080 34008 22120
rect 34054 22108 34060 22160
rect 34112 22148 34118 22160
rect 34698 22148 34704 22160
rect 34112 22120 34704 22148
rect 34112 22108 34118 22120
rect 34698 22108 34704 22120
rect 34756 22148 34762 22160
rect 46385 22151 46443 22157
rect 34756 22120 35940 22148
rect 34756 22108 34762 22120
rect 35069 22083 35127 22089
rect 35069 22080 35081 22083
rect 33980 22052 35081 22080
rect 35069 22049 35081 22052
rect 35115 22080 35127 22083
rect 35618 22080 35624 22092
rect 35115 22052 35624 22080
rect 35115 22049 35127 22052
rect 35069 22043 35127 22049
rect 35618 22040 35624 22052
rect 35676 22040 35682 22092
rect 35912 22089 35940 22120
rect 46385 22117 46397 22151
rect 46431 22148 46443 22151
rect 46750 22148 46756 22160
rect 46431 22120 46756 22148
rect 46431 22117 46443 22120
rect 46385 22111 46443 22117
rect 46750 22108 46756 22120
rect 46808 22108 46814 22160
rect 47320 22148 47348 22176
rect 48314 22148 48320 22160
rect 47320 22120 48320 22148
rect 48314 22108 48320 22120
rect 48372 22108 48378 22160
rect 48516 22148 48544 22188
rect 48593 22185 48605 22219
rect 48639 22216 48651 22219
rect 48639 22188 49004 22216
rect 48639 22185 48651 22188
rect 48593 22179 48651 22185
rect 48777 22151 48835 22157
rect 48777 22148 48789 22151
rect 48516 22120 48789 22148
rect 48777 22117 48789 22120
rect 48823 22117 48835 22151
rect 48777 22111 48835 22117
rect 48976 22092 49004 22188
rect 35897 22083 35955 22089
rect 35897 22049 35909 22083
rect 35943 22049 35955 22083
rect 35897 22043 35955 22049
rect 37826 22040 37832 22092
rect 37884 22040 37890 22092
rect 47394 22080 47400 22092
rect 46216 22052 46612 22080
rect 28767 21984 29868 22012
rect 28767 21981 28779 21984
rect 28721 21975 28779 21981
rect 28828 21888 28856 21984
rect 30006 21972 30012 22024
rect 30064 22012 30070 22024
rect 30466 22021 30472 22024
rect 30193 22015 30251 22021
rect 30193 22012 30205 22015
rect 30064 21984 30205 22012
rect 30064 21972 30070 21984
rect 30193 21981 30205 21984
rect 30239 21981 30251 22015
rect 30193 21975 30251 21981
rect 30460 21975 30472 22021
rect 30466 21972 30472 21975
rect 30524 21972 30530 22024
rect 35250 21972 35256 22024
rect 35308 21972 35314 22024
rect 35437 22015 35495 22021
rect 35437 21981 35449 22015
rect 35483 22012 35495 22015
rect 35713 22015 35771 22021
rect 35713 22012 35725 22015
rect 35483 21984 35725 22012
rect 35483 21981 35495 21984
rect 35437 21975 35495 21981
rect 35713 21981 35725 21984
rect 35759 21981 35771 22015
rect 37734 22012 37740 22024
rect 35713 21975 35771 21981
rect 36556 21984 37740 22012
rect 30098 21904 30104 21956
rect 30156 21904 30162 21956
rect 36142 21947 36200 21953
rect 36142 21944 36154 21947
rect 35544 21916 36154 21944
rect 27614 21836 27620 21888
rect 27672 21876 27678 21888
rect 27893 21879 27951 21885
rect 27893 21876 27905 21879
rect 27672 21848 27905 21876
rect 27672 21836 27678 21848
rect 27893 21845 27905 21848
rect 27939 21845 27951 21879
rect 27893 21839 27951 21845
rect 28810 21836 28816 21888
rect 28868 21836 28874 21888
rect 30009 21879 30067 21885
rect 30009 21845 30021 21879
rect 30055 21876 30067 21879
rect 30116 21876 30144 21904
rect 35544 21885 35572 21916
rect 36142 21913 36154 21916
rect 36188 21913 36200 21947
rect 36142 21907 36200 21913
rect 36556 21888 36584 21984
rect 37734 21972 37740 21984
rect 37792 21972 37798 22024
rect 38096 22015 38154 22021
rect 38096 21981 38108 22015
rect 38142 22012 38154 22015
rect 38654 22012 38660 22024
rect 38142 21984 38660 22012
rect 38142 21981 38154 21984
rect 38096 21975 38154 21981
rect 38654 21972 38660 21984
rect 38712 21972 38718 22024
rect 44818 21972 44824 22024
rect 44876 21972 44882 22024
rect 45738 21972 45744 22024
rect 45796 21972 45802 22024
rect 37458 21904 37464 21956
rect 37516 21904 37522 21956
rect 46216 21888 46244 22052
rect 46477 22015 46535 22021
rect 46477 22012 46489 22015
rect 46400 21984 46489 22012
rect 30055 21848 30144 21876
rect 35529 21879 35587 21885
rect 30055 21845 30067 21848
rect 30009 21839 30067 21845
rect 35529 21845 35541 21879
rect 35575 21845 35587 21879
rect 35529 21839 35587 21845
rect 36538 21836 36544 21888
rect 36596 21836 36602 21888
rect 37274 21836 37280 21888
rect 37332 21876 37338 21888
rect 37645 21879 37703 21885
rect 37645 21876 37657 21879
rect 37332 21848 37657 21876
rect 37332 21836 37338 21848
rect 37645 21845 37657 21848
rect 37691 21845 37703 21879
rect 37645 21839 37703 21845
rect 39206 21836 39212 21888
rect 39264 21836 39270 21888
rect 46198 21836 46204 21888
rect 46256 21836 46262 21888
rect 46400 21876 46428 21984
rect 46477 21981 46489 21984
rect 46523 21981 46535 22015
rect 46477 21975 46535 21981
rect 46584 21944 46612 22052
rect 46768 22052 47400 22080
rect 46658 21972 46664 22024
rect 46716 21972 46722 22024
rect 46768 22021 46796 22052
rect 47394 22040 47400 22052
rect 47452 22040 47458 22092
rect 48866 22040 48872 22092
rect 48924 22040 48930 22092
rect 48958 22040 48964 22092
rect 49016 22040 49022 22092
rect 46753 22015 46811 22021
rect 46753 21981 46765 22015
rect 46799 21981 46811 22015
rect 46753 21975 46811 21981
rect 46845 22015 46903 22021
rect 46845 21981 46857 22015
rect 46891 21981 46903 22015
rect 46845 21975 46903 21981
rect 46860 21944 46888 21975
rect 46934 21972 46940 22024
rect 46992 22012 46998 22024
rect 46992 21984 47440 22012
rect 46992 21972 46998 21984
rect 47302 21944 47308 21956
rect 46584 21916 46888 21944
rect 46952 21916 47308 21944
rect 46952 21876 46980 21916
rect 47302 21904 47308 21916
rect 47360 21904 47366 21956
rect 47412 21944 47440 21984
rect 47486 21972 47492 22024
rect 47544 21972 47550 22024
rect 47670 21972 47676 22024
rect 47728 21972 47734 22024
rect 47765 22015 47823 22021
rect 47765 21981 47777 22015
rect 47811 22012 47823 22015
rect 48041 22015 48099 22021
rect 47811 21984 47900 22012
rect 47811 21981 47823 21984
rect 47765 21975 47823 21981
rect 47872 21944 47900 21984
rect 48041 21981 48053 22015
rect 48087 21981 48099 22015
rect 48041 21975 48099 21981
rect 47412 21916 47900 21944
rect 48056 21944 48084 21975
rect 48222 21972 48228 22024
rect 48280 21972 48286 22024
rect 48314 21972 48320 22024
rect 48372 21972 48378 22024
rect 48976 22012 49004 22040
rect 49053 22015 49111 22021
rect 49053 22012 49065 22015
rect 48976 21984 49065 22012
rect 49053 21981 49065 21984
rect 49099 21981 49111 22015
rect 49053 21975 49111 21981
rect 49602 21972 49608 22024
rect 49660 21972 49666 22024
rect 49694 21972 49700 22024
rect 49752 21972 49758 22024
rect 48130 21944 48136 21956
rect 48056 21916 48136 21944
rect 47872 21888 47900 21916
rect 48130 21904 48136 21916
rect 48188 21904 48194 21956
rect 48406 21904 48412 21956
rect 48464 21944 48470 21956
rect 49712 21944 49740 21972
rect 48464 21916 49740 21944
rect 48464 21904 48470 21916
rect 46400 21848 46980 21876
rect 47026 21836 47032 21888
rect 47084 21836 47090 21888
rect 47854 21836 47860 21888
rect 47912 21836 47918 21888
rect 48590 21836 48596 21888
rect 48648 21885 48654 21888
rect 48648 21879 48667 21885
rect 48655 21845 48667 21879
rect 48648 21839 48667 21845
rect 48648 21836 48654 21839
rect 49234 21836 49240 21888
rect 49292 21836 49298 21888
rect 49697 21879 49755 21885
rect 49697 21845 49709 21879
rect 49743 21876 49755 21879
rect 49786 21876 49792 21888
rect 49743 21848 49792 21876
rect 49743 21845 49755 21848
rect 49697 21839 49755 21845
rect 49786 21836 49792 21848
rect 49844 21836 49850 21888
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 29086 21632 29092 21684
rect 29144 21632 29150 21684
rect 30742 21632 30748 21684
rect 30800 21672 30806 21684
rect 30853 21675 30911 21681
rect 30853 21672 30865 21675
rect 30800 21644 30865 21672
rect 30800 21632 30806 21644
rect 30853 21641 30865 21644
rect 30899 21641 30911 21675
rect 30853 21635 30911 21641
rect 31018 21632 31024 21684
rect 31076 21632 31082 21684
rect 34054 21632 34060 21684
rect 34112 21632 34118 21684
rect 35250 21632 35256 21684
rect 35308 21632 35314 21684
rect 35342 21632 35348 21684
rect 35400 21672 35406 21684
rect 35529 21675 35587 21681
rect 35529 21672 35541 21675
rect 35400 21644 35541 21672
rect 35400 21632 35406 21644
rect 35529 21641 35541 21644
rect 35575 21641 35587 21675
rect 35529 21635 35587 21641
rect 35897 21675 35955 21681
rect 35897 21641 35909 21675
rect 35943 21672 35955 21675
rect 35943 21644 37044 21672
rect 35943 21641 35955 21644
rect 35897 21635 35955 21641
rect 26602 21604 26608 21616
rect 25424 21576 26608 21604
rect 934 21496 940 21548
rect 992 21536 998 21548
rect 1489 21539 1547 21545
rect 1489 21536 1501 21539
rect 992 21508 1501 21536
rect 992 21496 998 21508
rect 1489 21505 1501 21508
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 24946 21428 24952 21480
rect 25004 21468 25010 21480
rect 25424 21477 25452 21576
rect 26602 21564 26608 21576
rect 26660 21604 26666 21616
rect 28902 21604 28908 21616
rect 26660 21576 27384 21604
rect 26660 21564 26666 21576
rect 25676 21539 25734 21545
rect 25676 21505 25688 21539
rect 25722 21536 25734 21539
rect 26973 21539 27031 21545
rect 26973 21536 26985 21539
rect 25722 21508 26985 21536
rect 25722 21505 25734 21508
rect 25676 21499 25734 21505
rect 26973 21505 26985 21508
rect 27019 21505 27031 21539
rect 26973 21499 27031 21505
rect 27154 21496 27160 21548
rect 27212 21496 27218 21548
rect 25409 21471 25467 21477
rect 25409 21468 25421 21471
rect 25004 21440 25421 21468
rect 25004 21428 25010 21440
rect 25409 21437 25421 21440
rect 25455 21437 25467 21471
rect 27356 21468 27384 21576
rect 27816 21576 28908 21604
rect 27430 21496 27436 21548
rect 27488 21496 27494 21548
rect 27614 21496 27620 21548
rect 27672 21496 27678 21548
rect 27709 21471 27767 21477
rect 27709 21468 27721 21471
rect 27356 21440 27721 21468
rect 25409 21431 25467 21437
rect 27709 21437 27721 21440
rect 27755 21468 27767 21471
rect 27816 21468 27844 21576
rect 28902 21564 28908 21576
rect 28960 21604 28966 21616
rect 30006 21604 30012 21616
rect 28960 21576 30012 21604
rect 28960 21564 28966 21576
rect 30006 21564 30012 21576
rect 30064 21564 30070 21616
rect 30650 21564 30656 21616
rect 30708 21564 30714 21616
rect 34072 21604 34100 21632
rect 32324 21576 34100 21604
rect 35268 21604 35296 21632
rect 36357 21607 36415 21613
rect 36357 21604 36369 21607
rect 35268 21576 36369 21604
rect 27976 21539 28034 21545
rect 27976 21505 27988 21539
rect 28022 21536 28034 21539
rect 28718 21536 28724 21548
rect 28022 21508 28724 21536
rect 28022 21505 28034 21508
rect 27976 21499 28034 21505
rect 28718 21496 28724 21508
rect 28776 21496 28782 21548
rect 29086 21496 29092 21548
rect 29144 21536 29150 21548
rect 29457 21539 29515 21545
rect 29457 21536 29469 21539
rect 29144 21508 29469 21536
rect 29144 21496 29150 21508
rect 29457 21505 29469 21508
rect 29503 21505 29515 21539
rect 29457 21499 29515 21505
rect 31754 21496 31760 21548
rect 31812 21536 31818 21548
rect 32324 21545 32352 21576
rect 36357 21573 36369 21576
rect 36403 21573 36415 21607
rect 36357 21567 36415 21573
rect 36464 21576 36676 21604
rect 32582 21545 32588 21548
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 31812 21508 32321 21536
rect 31812 21496 31818 21508
rect 32309 21505 32321 21508
rect 32355 21505 32367 21539
rect 32309 21499 32367 21505
rect 32576 21499 32588 21545
rect 32582 21496 32588 21499
rect 32640 21496 32646 21548
rect 33502 21496 33508 21548
rect 33560 21536 33566 21548
rect 34517 21539 34575 21545
rect 34517 21536 34529 21539
rect 33560 21508 34529 21536
rect 33560 21496 33566 21508
rect 34517 21505 34529 21508
rect 34563 21505 34575 21539
rect 34517 21499 34575 21505
rect 33781 21471 33839 21477
rect 33781 21468 33793 21471
rect 27755 21440 27844 21468
rect 33704 21440 33793 21468
rect 27755 21437 27767 21440
rect 27709 21431 27767 21437
rect 33704 21412 33732 21440
rect 33781 21437 33793 21440
rect 33827 21437 33839 21471
rect 33781 21431 33839 21437
rect 35989 21471 36047 21477
rect 35989 21437 36001 21471
rect 36035 21437 36047 21471
rect 35989 21431 36047 21437
rect 36173 21471 36231 21477
rect 36173 21437 36185 21471
rect 36219 21468 36231 21471
rect 36464 21468 36492 21576
rect 36648 21548 36676 21576
rect 36538 21496 36544 21548
rect 36596 21496 36602 21548
rect 36630 21496 36636 21548
rect 36688 21496 36694 21548
rect 36725 21539 36783 21545
rect 36725 21505 36737 21539
rect 36771 21505 36783 21539
rect 36725 21499 36783 21505
rect 36863 21539 36921 21545
rect 36863 21505 36875 21539
rect 36909 21505 36921 21539
rect 36863 21499 36921 21505
rect 36740 21468 36768 21499
rect 36219 21440 36492 21468
rect 36648 21440 36768 21468
rect 36878 21468 36906 21499
rect 37016 21477 37044 21644
rect 37458 21632 37464 21684
rect 37516 21672 37522 21684
rect 38473 21675 38531 21681
rect 38473 21672 38485 21675
rect 37516 21644 38485 21672
rect 37516 21632 37522 21644
rect 38473 21641 38485 21644
rect 38519 21641 38531 21675
rect 39206 21672 39212 21684
rect 38473 21635 38531 21641
rect 38580 21644 39212 21672
rect 38286 21604 38292 21616
rect 37936 21576 38292 21604
rect 37936 21545 37964 21576
rect 38286 21564 38292 21576
rect 38344 21604 38350 21616
rect 38580 21613 38608 21644
rect 39206 21632 39212 21644
rect 39264 21632 39270 21684
rect 46109 21675 46167 21681
rect 46109 21672 46121 21675
rect 43916 21644 46121 21672
rect 43916 21613 43944 21644
rect 46109 21641 46121 21644
rect 46155 21641 46167 21675
rect 46109 21635 46167 21641
rect 46216 21644 46704 21672
rect 46216 21616 46244 21644
rect 38565 21607 38623 21613
rect 38565 21604 38577 21607
rect 38344 21576 38577 21604
rect 38344 21564 38350 21576
rect 38565 21573 38577 21576
rect 38611 21573 38623 21607
rect 38765 21607 38823 21613
rect 38765 21604 38777 21607
rect 38565 21567 38623 21573
rect 38672 21576 38777 21604
rect 37921 21539 37979 21545
rect 37921 21505 37933 21539
rect 37967 21505 37979 21539
rect 37921 21499 37979 21505
rect 37001 21471 37059 21477
rect 36878 21440 36952 21468
rect 36219 21437 36231 21440
rect 36173 21431 36231 21437
rect 33686 21360 33692 21412
rect 33744 21360 33750 21412
rect 36004 21400 36032 21431
rect 36648 21400 36676 21440
rect 36004 21372 36676 21400
rect 36096 21344 36124 21372
rect 36924 21344 36952 21440
rect 37001 21437 37013 21471
rect 37047 21437 37059 21471
rect 37001 21431 37059 21437
rect 1762 21292 1768 21344
rect 1820 21292 1826 21344
rect 26789 21335 26847 21341
rect 26789 21301 26801 21335
rect 26835 21332 26847 21335
rect 26878 21332 26884 21344
rect 26835 21304 26884 21332
rect 26835 21301 26847 21304
rect 26789 21295 26847 21301
rect 26878 21292 26884 21304
rect 26936 21332 26942 21344
rect 28074 21332 28080 21344
rect 26936 21304 28080 21332
rect 26936 21292 26942 21304
rect 28074 21292 28080 21304
rect 28132 21292 28138 21344
rect 30098 21292 30104 21344
rect 30156 21292 30162 21344
rect 30374 21292 30380 21344
rect 30432 21332 30438 21344
rect 30837 21335 30895 21341
rect 30837 21332 30849 21335
rect 30432 21304 30849 21332
rect 30432 21292 30438 21304
rect 30837 21301 30849 21304
rect 30883 21301 30895 21335
rect 30837 21295 30895 21301
rect 33410 21292 33416 21344
rect 33468 21332 33474 21344
rect 34425 21335 34483 21341
rect 34425 21332 34437 21335
rect 33468 21304 34437 21332
rect 33468 21292 33474 21304
rect 34425 21301 34437 21304
rect 34471 21301 34483 21335
rect 34425 21295 34483 21301
rect 34790 21292 34796 21344
rect 34848 21332 34854 21344
rect 35161 21335 35219 21341
rect 35161 21332 35173 21335
rect 34848 21304 35173 21332
rect 34848 21292 34854 21304
rect 35161 21301 35173 21304
rect 35207 21301 35219 21335
rect 35161 21295 35219 21301
rect 36078 21292 36084 21344
rect 36136 21292 36142 21344
rect 36906 21292 36912 21344
rect 36964 21292 36970 21344
rect 37016 21332 37044 21431
rect 37734 21428 37740 21480
rect 37792 21468 37798 21480
rect 38672 21468 38700 21576
rect 38765 21573 38777 21576
rect 38811 21573 38823 21607
rect 38765 21567 38823 21573
rect 43901 21607 43959 21613
rect 43901 21573 43913 21607
rect 43947 21573 43959 21607
rect 43901 21567 43959 21573
rect 44542 21564 44548 21616
rect 44600 21564 44606 21616
rect 45738 21604 45744 21616
rect 45388 21576 45744 21604
rect 42426 21496 42432 21548
rect 42484 21536 42490 21548
rect 42702 21536 42708 21548
rect 42484 21508 42708 21536
rect 42484 21496 42490 21508
rect 42702 21496 42708 21508
rect 42760 21496 42766 21548
rect 42794 21496 42800 21548
rect 42852 21536 42858 21548
rect 43622 21536 43628 21548
rect 42852 21508 43628 21536
rect 42852 21496 42858 21508
rect 43622 21496 43628 21508
rect 43680 21496 43686 21548
rect 45388 21477 45416 21576
rect 45738 21564 45744 21576
rect 45796 21564 45802 21616
rect 46198 21564 46204 21616
rect 46256 21564 46262 21616
rect 46474 21564 46480 21616
rect 46532 21564 46538 21616
rect 46566 21564 46572 21616
rect 46624 21564 46630 21616
rect 46290 21496 46296 21548
rect 46348 21496 46354 21548
rect 46382 21496 46388 21548
rect 46440 21496 46446 21548
rect 46676 21545 46704 21644
rect 46750 21632 46756 21684
rect 46808 21632 46814 21684
rect 46934 21632 46940 21684
rect 46992 21632 46998 21684
rect 47026 21632 47032 21684
rect 47084 21632 47090 21684
rect 47136 21644 47440 21672
rect 46768 21604 46796 21632
rect 46768 21576 46888 21604
rect 46860 21545 46888 21576
rect 46952 21545 46980 21632
rect 46676 21539 46745 21545
rect 46676 21508 46699 21539
rect 46687 21505 46699 21508
rect 46733 21505 46745 21539
rect 46687 21499 46745 21505
rect 46845 21539 46903 21545
rect 46845 21505 46857 21539
rect 46891 21505 46903 21539
rect 46845 21499 46903 21505
rect 46937 21539 46995 21545
rect 46937 21505 46949 21539
rect 46983 21505 46995 21539
rect 46937 21499 46995 21505
rect 47026 21496 47032 21548
rect 47084 21536 47090 21548
rect 47136 21545 47164 21644
rect 47302 21604 47308 21616
rect 47228 21576 47308 21604
rect 47228 21545 47256 21576
rect 47302 21564 47308 21576
rect 47360 21564 47366 21616
rect 47412 21545 47440 21644
rect 47854 21632 47860 21684
rect 47912 21672 47918 21684
rect 48590 21672 48596 21684
rect 47912 21644 48596 21672
rect 47912 21632 47918 21644
rect 48590 21632 48596 21644
rect 48648 21632 48654 21684
rect 49234 21632 49240 21684
rect 49292 21632 49298 21684
rect 49252 21604 49280 21632
rect 47964 21576 49280 21604
rect 47121 21539 47179 21545
rect 47121 21536 47133 21539
rect 47084 21508 47133 21536
rect 47084 21496 47090 21508
rect 47121 21505 47133 21508
rect 47167 21505 47179 21539
rect 47121 21499 47179 21505
rect 47213 21539 47271 21545
rect 47213 21505 47225 21539
rect 47259 21505 47271 21539
rect 47213 21499 47271 21505
rect 47397 21539 47455 21545
rect 47397 21505 47409 21539
rect 47443 21505 47455 21539
rect 47397 21499 47455 21505
rect 47762 21496 47768 21548
rect 47820 21536 47826 21548
rect 47964 21536 47992 21576
rect 49786 21564 49792 21616
rect 49844 21564 49850 21616
rect 47820 21508 47992 21536
rect 48777 21539 48835 21545
rect 47820 21496 47826 21508
rect 48777 21505 48789 21539
rect 48823 21536 48835 21539
rect 48958 21536 48964 21548
rect 48823 21508 48964 21536
rect 48823 21505 48835 21508
rect 48777 21499 48835 21505
rect 48958 21496 48964 21508
rect 49016 21496 49022 21548
rect 51537 21539 51595 21545
rect 51537 21536 51549 21539
rect 50724 21508 51549 21536
rect 37792 21440 38700 21468
rect 45373 21471 45431 21477
rect 37792 21428 37798 21440
rect 45373 21437 45385 21471
rect 45419 21437 45431 21471
rect 45373 21431 45431 21437
rect 45557 21471 45615 21477
rect 45557 21437 45569 21471
rect 45603 21468 45615 21471
rect 46201 21471 46259 21477
rect 46201 21468 46213 21471
rect 45603 21440 46213 21468
rect 45603 21437 45615 21440
rect 45557 21431 45615 21437
rect 46201 21437 46213 21440
rect 46247 21437 46259 21471
rect 46201 21431 46259 21437
rect 46308 21400 46336 21496
rect 46474 21428 46480 21480
rect 46532 21468 46538 21480
rect 47305 21471 47363 21477
rect 47305 21468 47317 21471
rect 46532 21440 47317 21468
rect 46532 21428 46538 21440
rect 47305 21437 47317 21440
rect 47351 21437 47363 21471
rect 47305 21431 47363 21437
rect 47780 21400 47808 21496
rect 48222 21428 48228 21480
rect 48280 21468 48286 21480
rect 49053 21471 49111 21477
rect 49053 21468 49065 21471
rect 48280 21440 49065 21468
rect 48280 21428 48286 21440
rect 49053 21437 49065 21440
rect 49099 21437 49111 21471
rect 49053 21431 49111 21437
rect 46308 21372 47808 21400
rect 37274 21332 37280 21344
rect 37016 21304 37280 21332
rect 37274 21292 37280 21304
rect 37332 21332 37338 21344
rect 38749 21335 38807 21341
rect 38749 21332 38761 21335
rect 37332 21304 38761 21332
rect 37332 21292 37338 21304
rect 38749 21301 38761 21304
rect 38795 21301 38807 21335
rect 38749 21295 38807 21301
rect 38933 21335 38991 21341
rect 38933 21301 38945 21335
rect 38979 21332 38991 21335
rect 39022 21332 39028 21344
rect 38979 21304 39028 21332
rect 38979 21301 38991 21304
rect 38933 21295 38991 21301
rect 39022 21292 39028 21304
rect 39080 21292 39086 21344
rect 42518 21292 42524 21344
rect 42576 21292 42582 21344
rect 46382 21292 46388 21344
rect 46440 21332 46446 21344
rect 47486 21332 47492 21344
rect 46440 21304 47492 21332
rect 46440 21292 46446 21304
rect 47486 21292 47492 21304
rect 47544 21292 47550 21344
rect 48866 21292 48872 21344
rect 48924 21292 48930 21344
rect 49068 21332 49096 21431
rect 49326 21428 49332 21480
rect 49384 21428 49390 21480
rect 50724 21344 50752 21508
rect 51537 21505 51549 21508
rect 51583 21505 51595 21539
rect 51537 21499 51595 21505
rect 50893 21471 50951 21477
rect 50893 21437 50905 21471
rect 50939 21437 50951 21471
rect 50893 21431 50951 21437
rect 50062 21332 50068 21344
rect 49068 21304 50068 21332
rect 50062 21292 50068 21304
rect 50120 21292 50126 21344
rect 50706 21292 50712 21344
rect 50764 21292 50770 21344
rect 50798 21292 50804 21344
rect 50856 21332 50862 21344
rect 50908 21332 50936 21431
rect 50856 21304 50936 21332
rect 50856 21292 50862 21304
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 26605 21131 26663 21137
rect 26605 21097 26617 21131
rect 26651 21128 26663 21131
rect 27154 21128 27160 21140
rect 26651 21100 27160 21128
rect 26651 21097 26663 21100
rect 26605 21091 26663 21097
rect 27154 21088 27160 21100
rect 27212 21088 27218 21140
rect 28718 21088 28724 21140
rect 28776 21128 28782 21140
rect 29549 21131 29607 21137
rect 29549 21128 29561 21131
rect 28776 21100 29561 21128
rect 28776 21088 28782 21100
rect 29549 21097 29561 21100
rect 29595 21097 29607 21131
rect 29549 21091 29607 21097
rect 30098 21088 30104 21140
rect 30156 21088 30162 21140
rect 33410 21088 33416 21140
rect 33468 21088 33474 21140
rect 33686 21088 33692 21140
rect 33744 21088 33750 21140
rect 36906 21088 36912 21140
rect 36964 21088 36970 21140
rect 40034 21128 40040 21140
rect 39408 21100 40040 21128
rect 28534 21020 28540 21072
rect 28592 21060 28598 21072
rect 28592 21032 29868 21060
rect 28592 21020 28598 21032
rect 25501 20995 25559 21001
rect 25501 20961 25513 20995
rect 25547 20992 25559 20995
rect 25685 20995 25743 21001
rect 25685 20992 25697 20995
rect 25547 20964 25697 20992
rect 25547 20961 25559 20964
rect 25501 20955 25559 20961
rect 25685 20961 25697 20964
rect 25731 20961 25743 20995
rect 27430 20992 27436 21004
rect 25685 20955 25743 20961
rect 26804 20964 27436 20992
rect 26804 20936 26832 20964
rect 27430 20952 27436 20964
rect 27488 20952 27494 21004
rect 25409 20927 25467 20933
rect 25409 20893 25421 20927
rect 25455 20893 25467 20927
rect 25409 20887 25467 20893
rect 25593 20927 25651 20933
rect 25593 20893 25605 20927
rect 25639 20924 25651 20927
rect 26786 20924 26792 20936
rect 25639 20896 26792 20924
rect 25639 20893 25651 20896
rect 25593 20887 25651 20893
rect 25424 20856 25452 20887
rect 26786 20884 26792 20896
rect 26844 20884 26850 20936
rect 26878 20884 26884 20936
rect 26936 20884 26942 20936
rect 27065 20927 27123 20933
rect 27065 20893 27077 20927
rect 27111 20893 27123 20927
rect 27065 20887 27123 20893
rect 26510 20856 26516 20868
rect 25424 20828 26516 20856
rect 26510 20816 26516 20828
rect 26568 20816 26574 20868
rect 25774 20748 25780 20800
rect 25832 20788 25838 20800
rect 26329 20791 26387 20797
rect 26329 20788 26341 20791
rect 25832 20760 26341 20788
rect 25832 20748 25838 20760
rect 26329 20757 26341 20760
rect 26375 20757 26387 20791
rect 27080 20788 27108 20887
rect 27154 20884 27160 20936
rect 27212 20884 27218 20936
rect 27798 20924 27804 20936
rect 27264 20896 27804 20924
rect 27264 20788 27292 20896
rect 27798 20884 27804 20896
rect 27856 20924 27862 20936
rect 28810 20924 28816 20936
rect 27856 20896 28816 20924
rect 27856 20884 27862 20896
rect 28810 20884 28816 20896
rect 28868 20924 28874 20936
rect 29840 20933 29868 21032
rect 30116 20933 30144 21088
rect 32950 20952 32956 21004
rect 33008 20992 33014 21004
rect 33505 20995 33563 21001
rect 33505 20992 33517 20995
rect 33008 20964 33517 20992
rect 33008 20952 33014 20964
rect 33505 20961 33517 20964
rect 33551 20961 33563 20995
rect 33704 20992 33732 21088
rect 38565 21063 38623 21069
rect 38565 21060 38577 21063
rect 36832 21032 38577 21060
rect 33704 20964 34008 20992
rect 33505 20955 33563 20961
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 28868 20896 29745 20924
rect 28868 20884 28874 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 29825 20927 29883 20933
rect 29825 20893 29837 20927
rect 29871 20893 29883 20927
rect 29825 20887 29883 20893
rect 30009 20927 30067 20933
rect 30009 20893 30021 20927
rect 30055 20893 30067 20927
rect 30009 20887 30067 20893
rect 30101 20927 30159 20933
rect 30101 20893 30113 20927
rect 30147 20893 30159 20927
rect 30101 20887 30159 20893
rect 31665 20927 31723 20933
rect 31665 20893 31677 20927
rect 31711 20924 31723 20927
rect 31754 20924 31760 20936
rect 31711 20896 31760 20924
rect 31711 20893 31723 20896
rect 31665 20887 31723 20893
rect 29362 20816 29368 20868
rect 29420 20856 29426 20868
rect 30024 20856 30052 20887
rect 31754 20884 31760 20896
rect 31812 20884 31818 20936
rect 33226 20924 33232 20936
rect 32048 20896 33232 20924
rect 29420 20828 30052 20856
rect 31932 20859 31990 20865
rect 29420 20816 29426 20828
rect 31932 20825 31944 20859
rect 31978 20856 31990 20859
rect 32048 20856 32076 20896
rect 33226 20884 33232 20896
rect 33284 20884 33290 20936
rect 33594 20884 33600 20936
rect 33652 20884 33658 20936
rect 33980 20933 34008 20964
rect 34698 20952 34704 21004
rect 34756 20952 34762 21004
rect 33873 20927 33931 20933
rect 33873 20893 33885 20927
rect 33919 20893 33931 20927
rect 33873 20887 33931 20893
rect 33965 20927 34023 20933
rect 33965 20893 33977 20927
rect 34011 20893 34023 20927
rect 33965 20887 34023 20893
rect 33888 20856 33916 20887
rect 34790 20884 34796 20936
rect 34848 20924 34854 20936
rect 36832 20933 36860 21032
rect 38565 21029 38577 21032
rect 38611 21029 38623 21063
rect 38565 21023 38623 21029
rect 38654 21020 38660 21072
rect 38712 21060 38718 21072
rect 38749 21063 38807 21069
rect 38749 21060 38761 21063
rect 38712 21032 38761 21060
rect 38712 21020 38718 21032
rect 38749 21029 38761 21032
rect 38795 21029 38807 21063
rect 38749 21023 38807 21029
rect 34957 20927 35015 20933
rect 34957 20924 34969 20927
rect 34848 20896 34969 20924
rect 34848 20884 34854 20896
rect 34957 20893 34969 20896
rect 35003 20893 35015 20927
rect 34957 20887 35015 20893
rect 36817 20927 36875 20933
rect 36817 20893 36829 20927
rect 36863 20893 36875 20927
rect 36817 20887 36875 20893
rect 37001 20927 37059 20933
rect 37001 20893 37013 20927
rect 37047 20893 37059 20927
rect 37001 20887 37059 20893
rect 31978 20828 32076 20856
rect 33060 20828 33916 20856
rect 31978 20825 31990 20828
rect 31932 20819 31990 20825
rect 27080 20760 27292 20788
rect 26329 20751 26387 20757
rect 32214 20748 32220 20800
rect 32272 20788 32278 20800
rect 33060 20797 33088 20828
rect 36262 20816 36268 20868
rect 36320 20856 36326 20868
rect 36538 20856 36544 20868
rect 36320 20828 36544 20856
rect 36320 20816 36326 20828
rect 36538 20816 36544 20828
rect 36596 20856 36602 20868
rect 37016 20856 37044 20887
rect 38286 20884 38292 20936
rect 38344 20884 38350 20936
rect 39022 20884 39028 20936
rect 39080 20884 39086 20936
rect 39408 20933 39436 21100
rect 40034 21088 40040 21100
rect 40092 21088 40098 21140
rect 42518 21088 42524 21140
rect 42576 21088 42582 21140
rect 44542 21088 44548 21140
rect 44600 21088 44606 21140
rect 45738 21088 45744 21140
rect 45796 21088 45802 21140
rect 46198 21088 46204 21140
rect 46256 21088 46262 21140
rect 46385 21131 46443 21137
rect 46385 21097 46397 21131
rect 46431 21097 46443 21131
rect 46385 21091 46443 21097
rect 39577 21063 39635 21069
rect 39577 21029 39589 21063
rect 39623 21060 39635 21063
rect 39758 21060 39764 21072
rect 39623 21032 39764 21060
rect 39623 21029 39635 21032
rect 39577 21023 39635 21029
rect 39758 21020 39764 21032
rect 39816 21020 39822 21072
rect 39853 20995 39911 21001
rect 39592 20964 39804 20992
rect 39393 20927 39451 20933
rect 39393 20893 39405 20927
rect 39439 20893 39451 20927
rect 39393 20887 39451 20893
rect 36596 20828 37044 20856
rect 36596 20816 36602 20828
rect 38010 20816 38016 20868
rect 38068 20816 38074 20868
rect 38197 20859 38255 20865
rect 38197 20825 38209 20859
rect 38243 20856 38255 20859
rect 38243 20828 38700 20856
rect 38243 20825 38255 20828
rect 38197 20819 38255 20825
rect 33045 20791 33103 20797
rect 33045 20788 33057 20791
rect 32272 20760 33057 20788
rect 32272 20748 32278 20760
rect 33045 20757 33057 20760
rect 33091 20757 33103 20791
rect 33045 20751 33103 20757
rect 33137 20791 33195 20797
rect 33137 20757 33149 20791
rect 33183 20788 33195 20791
rect 33318 20788 33324 20800
rect 33183 20760 33324 20788
rect 33183 20757 33195 20760
rect 33137 20751 33195 20757
rect 33318 20748 33324 20760
rect 33376 20748 33382 20800
rect 33778 20748 33784 20800
rect 33836 20748 33842 20800
rect 34054 20748 34060 20800
rect 34112 20748 34118 20800
rect 36078 20748 36084 20800
rect 36136 20748 36142 20800
rect 37918 20748 37924 20800
rect 37976 20788 37982 20800
rect 38212 20788 38240 20819
rect 37976 20760 38240 20788
rect 37976 20748 37982 20760
rect 38286 20748 38292 20800
rect 38344 20788 38350 20800
rect 38381 20791 38439 20797
rect 38381 20788 38393 20791
rect 38344 20760 38393 20788
rect 38344 20748 38350 20760
rect 38381 20757 38393 20760
rect 38427 20757 38439 20791
rect 38672 20788 38700 20828
rect 38746 20816 38752 20868
rect 38804 20816 38810 20868
rect 38930 20788 38936 20800
rect 38672 20760 38936 20788
rect 38381 20751 38439 20757
rect 38930 20748 38936 20760
rect 38988 20748 38994 20800
rect 39040 20788 39068 20884
rect 39209 20859 39267 20865
rect 39209 20825 39221 20859
rect 39255 20856 39267 20859
rect 39592 20856 39620 20964
rect 39666 20884 39672 20936
rect 39724 20884 39730 20936
rect 39255 20828 39620 20856
rect 39776 20856 39804 20964
rect 39853 20961 39865 20995
rect 39899 20961 39911 20995
rect 42536 20992 42564 21088
rect 45756 21060 45784 21088
rect 46400 21060 46428 21091
rect 46566 21088 46572 21140
rect 46624 21128 46630 21140
rect 47213 21131 47271 21137
rect 47213 21128 47225 21131
rect 46624 21100 47225 21128
rect 46624 21088 46630 21100
rect 47213 21097 47225 21100
rect 47259 21097 47271 21131
rect 47213 21091 47271 21097
rect 45756 21032 46428 21060
rect 47228 21060 47256 21091
rect 47302 21088 47308 21140
rect 47360 21128 47366 21140
rect 47397 21131 47455 21137
rect 47397 21128 47409 21131
rect 47360 21100 47409 21128
rect 47360 21088 47366 21100
rect 47397 21097 47409 21100
rect 47443 21097 47455 21131
rect 47397 21091 47455 21097
rect 47673 21131 47731 21137
rect 47673 21097 47685 21131
rect 47719 21128 47731 21131
rect 47719 21100 47808 21128
rect 47719 21097 47731 21100
rect 47673 21091 47731 21097
rect 47228 21032 47716 21060
rect 46290 20992 46296 21004
rect 42536 20964 43852 20992
rect 39853 20955 39911 20961
rect 39868 20924 39896 20955
rect 41322 20924 41328 20936
rect 39868 20896 41328 20924
rect 40098 20859 40156 20865
rect 40098 20856 40110 20859
rect 39776 20828 40110 20856
rect 39255 20825 39267 20828
rect 39209 20819 39267 20825
rect 40098 20825 40110 20828
rect 40144 20825 40156 20859
rect 40098 20819 40156 20825
rect 40328 20800 40356 20896
rect 41322 20884 41328 20896
rect 41380 20884 41386 20936
rect 42334 20884 42340 20936
rect 42392 20924 42398 20936
rect 43824 20933 43852 20964
rect 44008 20964 45324 20992
rect 44008 20933 44036 20964
rect 45296 20936 45324 20964
rect 46032 20964 46296 20992
rect 42797 20927 42855 20933
rect 42797 20924 42809 20927
rect 42392 20896 42809 20924
rect 42392 20884 42398 20896
rect 42797 20893 42809 20896
rect 42843 20893 42855 20927
rect 42797 20887 42855 20893
rect 43441 20927 43499 20933
rect 43441 20893 43453 20927
rect 43487 20924 43499 20927
rect 43717 20927 43775 20933
rect 43717 20924 43729 20927
rect 43487 20896 43729 20924
rect 43487 20893 43499 20896
rect 43441 20887 43499 20893
rect 43717 20893 43729 20896
rect 43763 20893 43775 20927
rect 43717 20887 43775 20893
rect 43809 20927 43867 20933
rect 43809 20893 43821 20927
rect 43855 20893 43867 20927
rect 43809 20887 43867 20893
rect 43993 20927 44051 20933
rect 43993 20893 44005 20927
rect 44039 20893 44051 20927
rect 43993 20887 44051 20893
rect 44082 20884 44088 20936
rect 44140 20884 44146 20936
rect 44450 20924 44456 20936
rect 44192 20896 44456 20924
rect 41592 20859 41650 20865
rect 41592 20825 41604 20859
rect 41638 20856 41650 20859
rect 43533 20859 43591 20865
rect 43533 20856 43545 20859
rect 41638 20828 43545 20856
rect 41638 20825 41650 20828
rect 41592 20819 41650 20825
rect 43533 20825 43545 20828
rect 43579 20825 43591 20859
rect 43533 20819 43591 20825
rect 44192 20800 44220 20896
rect 44450 20884 44456 20896
rect 44508 20884 44514 20936
rect 45278 20884 45284 20936
rect 45336 20884 45342 20936
rect 46032 20933 46060 20964
rect 46290 20952 46296 20964
rect 46348 20952 46354 21004
rect 46017 20927 46075 20933
rect 46017 20893 46029 20927
rect 46063 20893 46075 20927
rect 46017 20887 46075 20893
rect 45833 20859 45891 20865
rect 45833 20825 45845 20859
rect 45879 20856 45891 20859
rect 46198 20856 46204 20868
rect 45879 20828 46204 20856
rect 45879 20825 45891 20828
rect 45833 20819 45891 20825
rect 46198 20816 46204 20828
rect 46256 20816 46262 20868
rect 46293 20859 46351 20865
rect 46293 20825 46305 20859
rect 46339 20825 46351 20859
rect 46400 20856 46428 21032
rect 47578 20992 47584 21004
rect 46768 20964 47584 20992
rect 46658 20884 46664 20936
rect 46716 20884 46722 20936
rect 46768 20933 46796 20964
rect 47578 20952 47584 20964
rect 47636 20952 47642 21004
rect 46753 20927 46811 20933
rect 46753 20893 46765 20927
rect 46799 20893 46811 20927
rect 46753 20887 46811 20893
rect 47489 20927 47547 20933
rect 47489 20893 47501 20927
rect 47535 20924 47547 20927
rect 47688 20924 47716 21032
rect 47535 20896 47716 20924
rect 47535 20893 47547 20896
rect 47489 20887 47547 20893
rect 47029 20859 47087 20865
rect 47029 20856 47041 20859
rect 46400 20828 47041 20856
rect 46293 20819 46351 20825
rect 47029 20825 47041 20828
rect 47075 20856 47087 20859
rect 47780 20856 47808 21100
rect 48314 21088 48320 21140
rect 48372 21128 48378 21140
rect 48774 21128 48780 21140
rect 48372 21100 48780 21128
rect 48372 21088 48378 21100
rect 48774 21088 48780 21100
rect 48832 21088 48838 21140
rect 48958 21088 48964 21140
rect 49016 21128 49022 21140
rect 49145 21131 49203 21137
rect 49145 21128 49157 21131
rect 49016 21100 49157 21128
rect 49016 21088 49022 21100
rect 49145 21097 49157 21100
rect 49191 21097 49203 21131
rect 49145 21091 49203 21097
rect 49237 21131 49295 21137
rect 49237 21097 49249 21131
rect 49283 21128 49295 21131
rect 49326 21128 49332 21140
rect 49283 21100 49332 21128
rect 49283 21097 49295 21100
rect 49237 21091 49295 21097
rect 49326 21088 49332 21100
rect 49384 21088 49390 21140
rect 50798 21060 50804 21072
rect 48608 21032 50804 21060
rect 48608 20868 48636 21032
rect 50798 21020 50804 21032
rect 50856 21020 50862 21072
rect 48866 20952 48872 21004
rect 48924 20992 48930 21004
rect 48924 20964 49556 20992
rect 48924 20952 48930 20964
rect 49528 20933 49556 20964
rect 49694 20952 49700 21004
rect 49752 20952 49758 21004
rect 49881 20995 49939 21001
rect 49881 20961 49893 20995
rect 49927 20992 49939 20995
rect 50706 20992 50712 21004
rect 49927 20964 50712 20992
rect 49927 20961 49939 20964
rect 49881 20955 49939 20961
rect 50706 20952 50712 20964
rect 50764 20952 50770 21004
rect 49421 20927 49479 20933
rect 49421 20926 49433 20927
rect 49344 20898 49433 20926
rect 47075 20828 47808 20856
rect 47075 20825 47087 20828
rect 47029 20819 47087 20825
rect 39574 20788 39580 20800
rect 39040 20760 39580 20788
rect 39574 20748 39580 20760
rect 39632 20748 39638 20800
rect 40310 20748 40316 20800
rect 40368 20748 40374 20800
rect 40402 20748 40408 20800
rect 40460 20788 40466 20800
rect 41233 20791 41291 20797
rect 41233 20788 41245 20791
rect 40460 20760 41245 20788
rect 40460 20748 40466 20760
rect 41233 20757 41245 20760
rect 41279 20757 41291 20791
rect 41233 20751 41291 20757
rect 42334 20748 42340 20800
rect 42392 20788 42398 20800
rect 42705 20791 42763 20797
rect 42705 20788 42717 20791
rect 42392 20760 42717 20788
rect 42392 20748 42398 20760
rect 42705 20757 42717 20760
rect 42751 20757 42763 20791
rect 42705 20751 42763 20757
rect 44174 20748 44180 20800
rect 44232 20748 44238 20800
rect 46308 20788 46336 20819
rect 48590 20816 48596 20868
rect 48648 20816 48654 20868
rect 46566 20788 46572 20800
rect 46308 20760 46572 20788
rect 46566 20748 46572 20760
rect 46624 20748 46630 20800
rect 46934 20748 46940 20800
rect 46992 20748 46998 20800
rect 47239 20791 47297 20797
rect 47239 20757 47251 20791
rect 47285 20788 47297 20791
rect 47762 20788 47768 20800
rect 47285 20760 47768 20788
rect 47285 20757 47297 20760
rect 47239 20751 47297 20757
rect 47762 20748 47768 20760
rect 47820 20748 47826 20800
rect 47854 20748 47860 20800
rect 47912 20748 47918 20800
rect 48498 20748 48504 20800
rect 48556 20788 48562 20800
rect 48777 20791 48835 20797
rect 48777 20788 48789 20791
rect 48556 20760 48789 20788
rect 48556 20748 48562 20760
rect 48777 20757 48789 20760
rect 48823 20757 48835 20791
rect 48777 20751 48835 20757
rect 48866 20748 48872 20800
rect 48924 20748 48930 20800
rect 48961 20791 49019 20797
rect 48961 20757 48973 20791
rect 49007 20788 49019 20791
rect 49142 20788 49148 20800
rect 49007 20760 49148 20788
rect 49007 20757 49019 20760
rect 48961 20751 49019 20757
rect 49142 20748 49148 20760
rect 49200 20748 49206 20800
rect 49344 20788 49372 20898
rect 49421 20893 49433 20898
rect 49467 20893 49479 20927
rect 49421 20887 49479 20893
rect 49513 20927 49571 20933
rect 49513 20893 49525 20927
rect 49559 20893 49571 20927
rect 49513 20887 49571 20893
rect 49605 20927 49663 20933
rect 49605 20893 49617 20927
rect 49651 20924 49663 20927
rect 49712 20924 49740 20952
rect 50341 20927 50399 20933
rect 50341 20924 50353 20927
rect 49651 20896 49740 20924
rect 49896 20896 50353 20924
rect 49651 20893 49663 20896
rect 49605 20887 49663 20893
rect 49896 20868 49924 20896
rect 50341 20893 50353 20896
rect 50387 20893 50399 20927
rect 50341 20887 50399 20893
rect 50430 20884 50436 20936
rect 50488 20884 50494 20936
rect 50525 20927 50583 20933
rect 50525 20893 50537 20927
rect 50571 20893 50583 20927
rect 50525 20887 50583 20893
rect 50617 20927 50675 20933
rect 50617 20893 50629 20927
rect 50663 20924 50675 20927
rect 50816 20924 50844 21020
rect 50663 20896 50844 20924
rect 50663 20893 50675 20896
rect 50617 20887 50675 20893
rect 49786 20865 49792 20868
rect 49743 20859 49792 20865
rect 49743 20825 49755 20859
rect 49789 20825 49792 20859
rect 49743 20819 49792 20825
rect 49786 20816 49792 20819
rect 49844 20816 49850 20868
rect 49878 20816 49884 20868
rect 49936 20816 49942 20868
rect 49970 20816 49976 20868
rect 50028 20856 50034 20868
rect 50540 20856 50568 20887
rect 50028 20828 50568 20856
rect 50028 20816 50034 20828
rect 50157 20791 50215 20797
rect 50157 20788 50169 20791
rect 49344 20760 50169 20788
rect 50157 20757 50169 20760
rect 50203 20757 50215 20791
rect 50157 20751 50215 20757
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 26786 20544 26792 20596
rect 26844 20544 26850 20596
rect 28074 20544 28080 20596
rect 28132 20544 28138 20596
rect 28261 20587 28319 20593
rect 28261 20553 28273 20587
rect 28307 20584 28319 20587
rect 32769 20587 32827 20593
rect 28307 20556 28764 20584
rect 28307 20553 28319 20556
rect 28261 20547 28319 20553
rect 25216 20519 25274 20525
rect 25216 20485 25228 20519
rect 25262 20516 25274 20519
rect 25774 20516 25780 20528
rect 25262 20488 25780 20516
rect 25262 20485 25274 20488
rect 25216 20479 25274 20485
rect 25774 20476 25780 20488
rect 25832 20476 25838 20528
rect 28736 20460 28764 20556
rect 32769 20553 32781 20587
rect 32815 20584 32827 20587
rect 33061 20587 33119 20593
rect 33061 20584 33073 20587
rect 32815 20556 33073 20584
rect 32815 20553 32827 20556
rect 32769 20547 32827 20553
rect 33061 20553 33073 20556
rect 33107 20553 33119 20587
rect 33061 20547 33119 20553
rect 33226 20544 33232 20596
rect 33284 20584 33290 20596
rect 33965 20587 34023 20593
rect 33965 20584 33977 20587
rect 33284 20556 33977 20584
rect 33284 20544 33290 20556
rect 33965 20553 33977 20556
rect 34011 20553 34023 20587
rect 33965 20547 34023 20553
rect 38746 20544 38752 20596
rect 38804 20584 38810 20596
rect 39485 20587 39543 20593
rect 39485 20584 39497 20587
rect 38804 20556 39497 20584
rect 38804 20544 38810 20556
rect 39485 20553 39497 20556
rect 39531 20553 39543 20587
rect 39485 20547 39543 20553
rect 39850 20544 39856 20596
rect 39908 20584 39914 20596
rect 40221 20587 40279 20593
rect 40221 20584 40233 20587
rect 39908 20556 40233 20584
rect 39908 20544 39914 20556
rect 40221 20553 40233 20556
rect 40267 20584 40279 20587
rect 40497 20587 40555 20593
rect 40497 20584 40509 20587
rect 40267 20556 40509 20584
rect 40267 20553 40279 20556
rect 40221 20547 40279 20553
rect 40497 20553 40509 20556
rect 40543 20553 40555 20587
rect 40497 20547 40555 20553
rect 40957 20587 41015 20593
rect 40957 20553 40969 20587
rect 41003 20553 41015 20587
rect 40957 20547 41015 20553
rect 41141 20587 41199 20593
rect 41141 20553 41153 20587
rect 41187 20584 41199 20587
rect 42334 20584 42340 20596
rect 41187 20556 42340 20584
rect 41187 20553 41199 20556
rect 41141 20547 41199 20553
rect 32030 20476 32036 20528
rect 32088 20516 32094 20528
rect 32861 20519 32919 20525
rect 32861 20516 32873 20519
rect 32088 20488 32873 20516
rect 32088 20476 32094 20488
rect 32861 20485 32873 20488
rect 32907 20485 32919 20519
rect 32861 20479 32919 20485
rect 34698 20476 34704 20528
rect 34756 20516 34762 20528
rect 34793 20519 34851 20525
rect 34793 20516 34805 20519
rect 34756 20488 34805 20516
rect 34756 20476 34762 20488
rect 34793 20485 34805 20488
rect 34839 20485 34851 20519
rect 37645 20519 37703 20525
rect 34793 20479 34851 20485
rect 36096 20488 36492 20516
rect 36096 20460 36124 20488
rect 24946 20408 24952 20460
rect 25004 20408 25010 20460
rect 26602 20408 26608 20460
rect 26660 20408 26666 20460
rect 28534 20408 28540 20460
rect 28592 20408 28598 20460
rect 28718 20408 28724 20460
rect 28776 20408 28782 20460
rect 28813 20451 28871 20457
rect 28813 20417 28825 20451
rect 28859 20448 28871 20451
rect 28902 20448 28908 20460
rect 28859 20420 28908 20448
rect 28859 20417 28871 20420
rect 28813 20411 28871 20417
rect 28902 20408 28908 20420
rect 28960 20408 28966 20460
rect 29086 20457 29092 20460
rect 29080 20411 29092 20457
rect 29086 20408 29092 20411
rect 29144 20408 29150 20460
rect 30558 20457 30564 20460
rect 30552 20411 30564 20457
rect 30558 20408 30564 20411
rect 30616 20408 30622 20460
rect 32214 20408 32220 20460
rect 32272 20408 32278 20460
rect 33318 20408 33324 20460
rect 33376 20408 33382 20460
rect 34057 20451 34115 20457
rect 34057 20417 34069 20451
rect 34103 20448 34115 20451
rect 34514 20448 34520 20460
rect 34103 20420 34520 20448
rect 34103 20417 34115 20420
rect 34057 20411 34115 20417
rect 34514 20408 34520 20420
rect 34572 20408 34578 20460
rect 35161 20451 35219 20457
rect 35161 20417 35173 20451
rect 35207 20448 35219 20451
rect 36078 20448 36084 20460
rect 35207 20420 36084 20448
rect 35207 20417 35219 20420
rect 35161 20411 35219 20417
rect 36078 20408 36084 20420
rect 36136 20408 36142 20460
rect 36262 20408 36268 20460
rect 36320 20408 36326 20460
rect 36464 20457 36492 20488
rect 37645 20485 37657 20519
rect 37691 20485 37703 20519
rect 37645 20479 37703 20485
rect 37861 20519 37919 20525
rect 37861 20485 37873 20519
rect 37907 20516 37919 20519
rect 37907 20488 38884 20516
rect 37907 20485 37919 20488
rect 37861 20479 37919 20485
rect 36449 20451 36507 20457
rect 36449 20417 36461 20451
rect 36495 20417 36507 20451
rect 36449 20411 36507 20417
rect 26421 20383 26479 20389
rect 26421 20349 26433 20383
rect 26467 20380 26479 20383
rect 27065 20383 27123 20389
rect 27065 20380 27077 20383
rect 26467 20352 27077 20380
rect 26467 20349 26479 20352
rect 26421 20343 26479 20349
rect 27065 20349 27077 20352
rect 27111 20349 27123 20383
rect 27065 20343 27123 20349
rect 26329 20315 26387 20321
rect 26329 20281 26341 20315
rect 26375 20312 26387 20315
rect 26436 20312 26464 20343
rect 26375 20284 26464 20312
rect 27080 20312 27108 20343
rect 27154 20340 27160 20392
rect 27212 20380 27218 20392
rect 27614 20380 27620 20392
rect 27212 20352 27620 20380
rect 27212 20340 27218 20352
rect 27614 20340 27620 20352
rect 27672 20340 27678 20392
rect 30006 20340 30012 20392
rect 30064 20380 30070 20392
rect 30285 20383 30343 20389
rect 30285 20380 30297 20383
rect 30064 20352 30297 20380
rect 30064 20340 30070 20352
rect 30285 20349 30297 20352
rect 30331 20349 30343 20383
rect 37660 20380 37688 20479
rect 38197 20451 38255 20457
rect 38197 20417 38209 20451
rect 38243 20448 38255 20451
rect 38654 20448 38660 20460
rect 38243 20420 38660 20448
rect 38243 20417 38255 20420
rect 38197 20411 38255 20417
rect 38654 20408 38660 20420
rect 38712 20408 38718 20460
rect 38856 20448 38884 20488
rect 38930 20476 38936 20528
rect 38988 20516 38994 20528
rect 40402 20516 40408 20528
rect 38988 20488 40408 20516
rect 38988 20476 38994 20488
rect 39684 20457 39712 20488
rect 40402 20476 40408 20488
rect 40460 20476 40466 20528
rect 40972 20516 41000 20547
rect 42334 20544 42340 20556
rect 42392 20544 42398 20596
rect 42702 20544 42708 20596
rect 42760 20544 42766 20596
rect 45278 20544 45284 20596
rect 45336 20544 45342 20596
rect 46750 20544 46756 20596
rect 46808 20584 46814 20596
rect 47397 20587 47455 20593
rect 47397 20584 47409 20587
rect 46808 20556 47409 20584
rect 46808 20544 46814 20556
rect 47397 20553 47409 20556
rect 47443 20553 47455 20587
rect 47397 20547 47455 20553
rect 48317 20587 48375 20593
rect 48317 20553 48329 20587
rect 48363 20553 48375 20587
rect 49142 20584 49148 20596
rect 48317 20547 48375 20553
rect 48884 20556 49148 20584
rect 40696 20488 41000 20516
rect 39669 20451 39727 20457
rect 38856 20420 38976 20448
rect 38010 20380 38016 20392
rect 37660 20352 38016 20380
rect 30285 20343 30343 20349
rect 38010 20340 38016 20352
rect 38068 20380 38074 20392
rect 38841 20383 38899 20389
rect 38841 20380 38853 20383
rect 38068 20352 38853 20380
rect 38068 20340 38074 20352
rect 38841 20349 38853 20352
rect 38887 20349 38899 20383
rect 38948 20380 38976 20420
rect 39669 20417 39681 20451
rect 39715 20417 39727 20451
rect 39669 20411 39727 20417
rect 39758 20408 39764 20460
rect 39816 20448 39822 20460
rect 40313 20451 40371 20457
rect 39816 20420 40172 20448
rect 39816 20408 39822 20420
rect 39776 20380 39804 20408
rect 38948 20352 39804 20380
rect 38841 20343 38899 20349
rect 27709 20315 27767 20321
rect 27709 20312 27721 20315
rect 27080 20284 27721 20312
rect 26375 20281 26387 20284
rect 26329 20275 26387 20281
rect 27709 20281 27721 20284
rect 27755 20281 27767 20315
rect 27709 20275 27767 20281
rect 30024 20284 30328 20312
rect 30024 20256 30052 20284
rect 27614 20204 27620 20256
rect 27672 20204 27678 20256
rect 28074 20204 28080 20256
rect 28132 20204 28138 20256
rect 28629 20247 28687 20253
rect 28629 20213 28641 20247
rect 28675 20244 28687 20247
rect 29730 20244 29736 20256
rect 28675 20216 29736 20244
rect 28675 20213 28687 20216
rect 28629 20207 28687 20213
rect 29730 20204 29736 20216
rect 29788 20204 29794 20256
rect 30006 20204 30012 20256
rect 30064 20204 30070 20256
rect 30190 20204 30196 20256
rect 30248 20204 30254 20256
rect 30300 20244 30328 20284
rect 31220 20284 33548 20312
rect 30650 20244 30656 20256
rect 30300 20216 30656 20244
rect 30650 20204 30656 20216
rect 30708 20244 30714 20256
rect 31220 20244 31248 20284
rect 30708 20216 31248 20244
rect 30708 20204 30714 20216
rect 31662 20204 31668 20256
rect 31720 20204 31726 20256
rect 33060 20253 33088 20284
rect 33045 20247 33103 20253
rect 33045 20213 33057 20247
rect 33091 20213 33103 20247
rect 33045 20207 33103 20213
rect 33229 20247 33287 20253
rect 33229 20213 33241 20247
rect 33275 20244 33287 20247
rect 33318 20244 33324 20256
rect 33275 20216 33324 20244
rect 33275 20213 33287 20216
rect 33229 20207 33287 20213
rect 33318 20204 33324 20216
rect 33376 20204 33382 20256
rect 33520 20244 33548 20284
rect 33594 20272 33600 20324
rect 33652 20312 33658 20324
rect 35713 20315 35771 20321
rect 35713 20312 35725 20315
rect 33652 20284 35725 20312
rect 33652 20272 33658 20284
rect 35713 20281 35725 20284
rect 35759 20281 35771 20315
rect 35713 20275 35771 20281
rect 37366 20272 37372 20324
rect 37424 20312 37430 20324
rect 38749 20315 38807 20321
rect 38749 20312 38761 20315
rect 37424 20284 38761 20312
rect 37424 20272 37430 20284
rect 38749 20281 38761 20284
rect 38795 20281 38807 20315
rect 38749 20275 38807 20281
rect 38856 20256 38884 20343
rect 40034 20340 40040 20392
rect 40092 20340 40098 20392
rect 40144 20380 40172 20420
rect 40313 20417 40325 20451
rect 40359 20448 40371 20451
rect 40494 20448 40500 20460
rect 40359 20420 40500 20448
rect 40359 20417 40371 20420
rect 40313 20411 40371 20417
rect 40494 20408 40500 20420
rect 40552 20408 40558 20460
rect 40696 20457 40724 20488
rect 41322 20476 41328 20528
rect 41380 20516 41386 20528
rect 42720 20516 42748 20544
rect 41380 20488 42748 20516
rect 41380 20476 41386 20488
rect 40589 20451 40647 20457
rect 40589 20417 40601 20451
rect 40635 20417 40647 20451
rect 40589 20411 40647 20417
rect 40681 20451 40739 20457
rect 40681 20417 40693 20451
rect 40727 20417 40739 20451
rect 40681 20411 40739 20417
rect 40604 20380 40632 20411
rect 40862 20408 40868 20460
rect 40920 20408 40926 20460
rect 41138 20451 41196 20457
rect 41138 20417 41150 20451
rect 41184 20448 41196 20451
rect 42426 20448 42432 20460
rect 41184 20420 42432 20448
rect 41184 20417 41196 20420
rect 41138 20411 41196 20417
rect 42426 20408 42432 20420
rect 42484 20408 42490 20460
rect 42536 20457 42564 20488
rect 43530 20476 43536 20528
rect 43588 20476 43594 20528
rect 47302 20516 47308 20528
rect 47136 20488 47308 20516
rect 42521 20451 42579 20457
rect 42521 20417 42533 20451
rect 42567 20417 42579 20451
rect 42521 20411 42579 20417
rect 45097 20451 45155 20457
rect 45097 20417 45109 20451
rect 45143 20448 45155 20451
rect 46106 20448 46112 20460
rect 45143 20420 46112 20448
rect 45143 20417 45155 20420
rect 45097 20411 45155 20417
rect 46106 20408 46112 20420
rect 46164 20408 46170 20460
rect 46474 20408 46480 20460
rect 46532 20448 46538 20460
rect 47136 20457 47164 20488
rect 47302 20476 47308 20488
rect 47360 20516 47366 20528
rect 48332 20516 48360 20547
rect 48884 20516 48912 20556
rect 49142 20544 49148 20556
rect 49200 20544 49206 20596
rect 49970 20544 49976 20596
rect 50028 20584 50034 20596
rect 50028 20556 50384 20584
rect 50028 20544 50034 20556
rect 50154 20516 50160 20528
rect 47360 20488 48912 20516
rect 48976 20488 50160 20516
rect 47360 20476 47366 20488
rect 46753 20451 46811 20457
rect 46753 20448 46765 20451
rect 46532 20420 46765 20448
rect 46532 20408 46538 20420
rect 46753 20417 46765 20420
rect 46799 20417 46811 20451
rect 46753 20411 46811 20417
rect 47121 20451 47179 20457
rect 47121 20417 47133 20451
rect 47167 20417 47179 20451
rect 47121 20411 47179 20417
rect 47213 20451 47271 20457
rect 47213 20417 47225 20451
rect 47259 20448 47271 20451
rect 47762 20448 47768 20460
rect 47259 20420 47768 20448
rect 47259 20417 47271 20420
rect 47213 20411 47271 20417
rect 47762 20408 47768 20420
rect 47820 20408 47826 20460
rect 48041 20451 48099 20457
rect 48041 20417 48053 20451
rect 48087 20448 48099 20451
rect 48314 20448 48320 20460
rect 48087 20420 48320 20448
rect 48087 20417 48099 20420
rect 48041 20411 48099 20417
rect 48314 20408 48320 20420
rect 48372 20408 48378 20460
rect 48409 20451 48467 20457
rect 48409 20417 48421 20451
rect 48455 20417 48467 20451
rect 48409 20411 48467 20417
rect 48685 20451 48743 20457
rect 48685 20417 48697 20451
rect 48731 20417 48743 20451
rect 48976 20448 49004 20488
rect 50154 20476 50160 20488
rect 50212 20516 50218 20528
rect 50249 20519 50307 20525
rect 50249 20516 50261 20519
rect 50212 20488 50261 20516
rect 50212 20476 50218 20488
rect 50249 20485 50261 20488
rect 50295 20485 50307 20519
rect 50249 20479 50307 20485
rect 50356 20479 50384 20556
rect 50341 20473 50399 20479
rect 48685 20411 48743 20417
rect 48792 20420 49004 20448
rect 40144 20352 40632 20380
rect 41598 20340 41604 20392
rect 41656 20340 41662 20392
rect 42794 20340 42800 20392
rect 42852 20340 42858 20392
rect 44361 20383 44419 20389
rect 44361 20380 44373 20383
rect 44284 20352 44373 20380
rect 40052 20312 40080 20340
rect 40313 20315 40371 20321
rect 40313 20312 40325 20315
rect 40052 20284 40325 20312
rect 40313 20281 40325 20284
rect 40359 20281 40371 20315
rect 40313 20275 40371 20281
rect 44284 20256 44312 20352
rect 44361 20349 44373 20352
rect 44407 20349 44419 20383
rect 44361 20343 44419 20349
rect 47673 20315 47731 20321
rect 47673 20312 47685 20315
rect 47044 20284 47685 20312
rect 47044 20256 47072 20284
rect 47673 20281 47685 20284
rect 47719 20281 47731 20315
rect 47854 20312 47860 20324
rect 47673 20275 47731 20281
rect 47780 20284 47860 20312
rect 33870 20244 33876 20256
rect 33520 20216 33876 20244
rect 33870 20204 33876 20216
rect 33928 20204 33934 20256
rect 36262 20204 36268 20256
rect 36320 20244 36326 20256
rect 36357 20247 36415 20253
rect 36357 20244 36369 20247
rect 36320 20216 36369 20244
rect 36320 20204 36326 20216
rect 36357 20213 36369 20216
rect 36403 20213 36415 20247
rect 36357 20207 36415 20213
rect 37829 20247 37887 20253
rect 37829 20213 37841 20247
rect 37875 20244 37887 20247
rect 37918 20244 37924 20256
rect 37875 20216 37924 20244
rect 37875 20213 37887 20216
rect 37829 20207 37887 20213
rect 37918 20204 37924 20216
rect 37976 20204 37982 20256
rect 38013 20247 38071 20253
rect 38013 20213 38025 20247
rect 38059 20244 38071 20247
rect 38654 20244 38660 20256
rect 38059 20216 38660 20244
rect 38059 20213 38071 20216
rect 38013 20207 38071 20213
rect 38654 20204 38660 20216
rect 38712 20204 38718 20256
rect 38838 20204 38844 20256
rect 38896 20204 38902 20256
rect 40678 20204 40684 20256
rect 40736 20204 40742 20256
rect 41506 20204 41512 20256
rect 41564 20204 41570 20256
rect 44266 20204 44272 20256
rect 44324 20204 44330 20256
rect 44450 20204 44456 20256
rect 44508 20244 44514 20256
rect 45005 20247 45063 20253
rect 45005 20244 45017 20247
rect 44508 20216 45017 20244
rect 44508 20204 44514 20216
rect 45005 20213 45017 20216
rect 45051 20213 45063 20247
rect 45005 20207 45063 20213
rect 46934 20204 46940 20256
rect 46992 20204 46998 20256
rect 47026 20204 47032 20256
rect 47084 20204 47090 20256
rect 47486 20204 47492 20256
rect 47544 20244 47550 20256
rect 47780 20244 47808 20284
rect 47854 20272 47860 20284
rect 47912 20312 47918 20324
rect 48133 20315 48191 20321
rect 48133 20312 48145 20315
rect 47912 20284 48145 20312
rect 47912 20272 47918 20284
rect 48133 20281 48145 20284
rect 48179 20281 48191 20315
rect 48424 20312 48452 20411
rect 48498 20340 48504 20392
rect 48556 20380 48562 20392
rect 48700 20380 48728 20411
rect 48792 20392 48820 20420
rect 49142 20408 49148 20460
rect 49200 20448 49206 20460
rect 49878 20448 49884 20460
rect 49200 20420 49884 20448
rect 49200 20408 49206 20420
rect 49878 20408 49884 20420
rect 49936 20448 49942 20460
rect 50065 20451 50123 20457
rect 50065 20448 50077 20451
rect 49936 20420 50077 20448
rect 49936 20408 49942 20420
rect 50065 20417 50077 20420
rect 50111 20417 50123 20451
rect 50341 20439 50353 20473
rect 50387 20439 50399 20473
rect 50341 20433 50399 20439
rect 50065 20411 50123 20417
rect 48556 20352 48728 20380
rect 48556 20340 48562 20352
rect 48774 20340 48780 20392
rect 48832 20340 48838 20392
rect 50080 20380 50108 20411
rect 50798 20408 50804 20460
rect 50856 20408 50862 20460
rect 50816 20380 50844 20408
rect 50080 20352 50844 20380
rect 49053 20315 49111 20321
rect 49053 20312 49065 20315
rect 48424 20284 49065 20312
rect 48133 20275 48191 20281
rect 49053 20281 49065 20284
rect 49099 20281 49111 20315
rect 49053 20275 49111 20281
rect 47544 20216 47808 20244
rect 47544 20204 47550 20216
rect 47946 20204 47952 20256
rect 48004 20244 48010 20256
rect 48590 20244 48596 20256
rect 48004 20216 48596 20244
rect 48004 20204 48010 20216
rect 48590 20204 48596 20216
rect 48648 20204 48654 20256
rect 49602 20204 49608 20256
rect 49660 20244 49666 20256
rect 50157 20247 50215 20253
rect 50157 20244 50169 20247
rect 49660 20216 50169 20244
rect 49660 20204 49666 20216
rect 50157 20213 50169 20216
rect 50203 20213 50215 20247
rect 50157 20207 50215 20213
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 26510 20000 26516 20052
rect 26568 20000 26574 20052
rect 27614 20000 27620 20052
rect 27672 20000 27678 20052
rect 27798 20000 27804 20052
rect 27856 20000 27862 20052
rect 29733 20043 29791 20049
rect 29733 20009 29745 20043
rect 29779 20040 29791 20043
rect 30006 20040 30012 20052
rect 29779 20012 30012 20040
rect 29779 20009 29791 20012
rect 29733 20003 29791 20009
rect 30006 20000 30012 20012
rect 30064 20000 30070 20052
rect 30558 20000 30564 20052
rect 30616 20040 30622 20052
rect 30653 20043 30711 20049
rect 30653 20040 30665 20043
rect 30616 20012 30665 20040
rect 30616 20000 30622 20012
rect 30653 20009 30665 20012
rect 30699 20009 30711 20043
rect 32030 20040 32036 20052
rect 30653 20003 30711 20009
rect 31128 20012 32036 20040
rect 27632 19972 27660 20000
rect 26436 19944 27660 19972
rect 27816 19972 27844 20000
rect 31021 19975 31079 19981
rect 31021 19972 31033 19975
rect 27816 19944 31033 19972
rect 26436 19904 26464 19944
rect 31021 19941 31033 19944
rect 31067 19941 31079 19975
rect 31021 19935 31079 19941
rect 26344 19876 26464 19904
rect 26605 19907 26663 19913
rect 26344 19845 26372 19876
rect 26605 19873 26617 19907
rect 26651 19904 26663 19907
rect 26694 19904 26700 19916
rect 26651 19876 26700 19904
rect 26651 19873 26663 19876
rect 26605 19867 26663 19873
rect 26694 19864 26700 19876
rect 26752 19864 26758 19916
rect 27341 19907 27399 19913
rect 27341 19873 27353 19907
rect 27387 19904 27399 19907
rect 27893 19907 27951 19913
rect 27893 19904 27905 19907
rect 27387 19876 27905 19904
rect 27387 19873 27399 19876
rect 27341 19867 27399 19873
rect 27893 19873 27905 19876
rect 27939 19904 27951 19907
rect 28626 19904 28632 19916
rect 27939 19876 28632 19904
rect 27939 19873 27951 19876
rect 27893 19867 27951 19873
rect 28626 19864 28632 19876
rect 28684 19864 28690 19916
rect 28902 19864 28908 19916
rect 28960 19904 28966 19916
rect 31128 19913 31156 20012
rect 32030 20000 32036 20012
rect 32088 20000 32094 20052
rect 32582 20000 32588 20052
rect 32640 20000 32646 20052
rect 32953 20043 33011 20049
rect 32953 20009 32965 20043
rect 32999 20040 33011 20043
rect 32999 20012 34468 20040
rect 32999 20009 33011 20012
rect 32953 20003 33011 20009
rect 31662 19932 31668 19984
rect 31720 19932 31726 19984
rect 33318 19972 33324 19984
rect 32784 19944 33324 19972
rect 29181 19907 29239 19913
rect 29181 19904 29193 19907
rect 28960 19876 29193 19904
rect 28960 19864 28966 19876
rect 29181 19873 29193 19876
rect 29227 19873 29239 19907
rect 29181 19867 29239 19873
rect 31113 19907 31171 19913
rect 31113 19873 31125 19907
rect 31159 19873 31171 19907
rect 31113 19867 31171 19873
rect 31481 19907 31539 19913
rect 31481 19873 31493 19907
rect 31527 19904 31539 19907
rect 31680 19904 31708 19932
rect 31527 19876 32352 19904
rect 31527 19873 31539 19876
rect 31481 19867 31539 19873
rect 26329 19839 26387 19845
rect 26329 19805 26341 19839
rect 26375 19805 26387 19839
rect 26329 19799 26387 19805
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19805 26479 19839
rect 26421 19799 26479 19805
rect 26436 19768 26464 19799
rect 27154 19796 27160 19848
rect 27212 19796 27218 19848
rect 27246 19796 27252 19848
rect 27304 19796 27310 19848
rect 27433 19839 27491 19845
rect 27433 19805 27445 19839
rect 27479 19836 27491 19839
rect 27522 19836 27528 19848
rect 27479 19808 27528 19836
rect 27479 19805 27491 19808
rect 27433 19799 27491 19805
rect 27522 19796 27528 19808
rect 27580 19796 27586 19848
rect 27614 19796 27620 19848
rect 27672 19796 27678 19848
rect 28077 19839 28135 19845
rect 28077 19805 28089 19839
rect 28123 19836 28135 19839
rect 28718 19836 28724 19848
rect 28123 19808 28724 19836
rect 28123 19805 28135 19808
rect 28077 19799 28135 19805
rect 28718 19796 28724 19808
rect 28776 19796 28782 19848
rect 29638 19836 29644 19848
rect 29564 19808 29644 19836
rect 26602 19768 26608 19780
rect 26436 19740 26608 19768
rect 26602 19728 26608 19740
rect 26660 19768 26666 19780
rect 27632 19768 27660 19796
rect 26660 19740 27660 19768
rect 26660 19728 26666 19740
rect 28442 19728 28448 19780
rect 28500 19728 28506 19780
rect 28626 19728 28632 19780
rect 28684 19768 28690 19780
rect 29564 19777 29592 19808
rect 29638 19796 29644 19808
rect 29696 19836 29702 19848
rect 30190 19836 30196 19848
rect 29696 19808 30196 19836
rect 29696 19796 29702 19808
rect 30190 19796 30196 19808
rect 30248 19796 30254 19848
rect 30837 19839 30895 19845
rect 30837 19805 30849 19839
rect 30883 19836 30895 19839
rect 31128 19836 31248 19838
rect 32214 19836 32220 19848
rect 30883 19830 31340 19836
rect 31496 19830 32220 19836
rect 30883 19810 32220 19830
rect 30883 19808 31156 19810
rect 31220 19808 32220 19810
rect 30883 19805 30895 19808
rect 30837 19799 30895 19805
rect 31312 19802 31524 19808
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 32324 19845 32352 19876
rect 32784 19845 32812 19944
rect 33318 19932 33324 19944
rect 33376 19932 33382 19984
rect 33413 19975 33471 19981
rect 33413 19941 33425 19975
rect 33459 19972 33471 19975
rect 33502 19972 33508 19984
rect 33459 19944 33508 19972
rect 33459 19941 33471 19944
rect 33413 19935 33471 19941
rect 33502 19932 33508 19944
rect 33560 19932 33566 19984
rect 33686 19932 33692 19984
rect 33744 19972 33750 19984
rect 34241 19975 34299 19981
rect 34241 19972 34253 19975
rect 33744 19944 34253 19972
rect 33744 19932 33750 19944
rect 34241 19941 34253 19944
rect 34287 19941 34299 19975
rect 34241 19935 34299 19941
rect 33229 19907 33287 19913
rect 33229 19873 33241 19907
rect 33275 19904 33287 19907
rect 33781 19907 33839 19913
rect 33781 19904 33793 19907
rect 33275 19876 33793 19904
rect 33275 19873 33287 19876
rect 33229 19867 33287 19873
rect 33781 19873 33793 19876
rect 33827 19873 33839 19907
rect 33781 19867 33839 19873
rect 33888 19876 34376 19904
rect 32309 19839 32367 19845
rect 32309 19805 32321 19839
rect 32355 19805 32367 19839
rect 32309 19799 32367 19805
rect 32769 19839 32827 19845
rect 32769 19805 32781 19839
rect 32815 19805 32827 19839
rect 32769 19799 32827 19805
rect 32861 19839 32919 19845
rect 32861 19805 32873 19839
rect 32907 19836 32919 19839
rect 33134 19836 33140 19848
rect 32907 19808 33140 19836
rect 32907 19805 32919 19808
rect 32861 19799 32919 19805
rect 33134 19796 33140 19808
rect 33192 19796 33198 19848
rect 33321 19839 33379 19845
rect 33321 19805 33333 19839
rect 33367 19836 33379 19839
rect 33502 19836 33508 19848
rect 33367 19808 33508 19836
rect 33367 19805 33379 19808
rect 33321 19799 33379 19805
rect 33502 19796 33508 19808
rect 33560 19796 33566 19848
rect 33594 19796 33600 19848
rect 33652 19796 33658 19848
rect 33686 19796 33692 19848
rect 33744 19836 33750 19848
rect 33888 19845 33916 19876
rect 34348 19848 34376 19876
rect 33873 19839 33931 19845
rect 33873 19836 33885 19839
rect 33744 19808 33885 19836
rect 33744 19796 33750 19808
rect 33873 19805 33885 19808
rect 33919 19805 33931 19839
rect 33873 19799 33931 19805
rect 33962 19796 33968 19848
rect 34020 19836 34026 19848
rect 34241 19839 34299 19845
rect 34241 19836 34253 19839
rect 34020 19808 34253 19836
rect 34020 19796 34026 19808
rect 34241 19805 34253 19808
rect 34287 19805 34299 19839
rect 34241 19799 34299 19805
rect 34330 19796 34336 19848
rect 34388 19796 34394 19848
rect 34440 19845 34468 20012
rect 37366 20000 37372 20052
rect 37424 20000 37430 20052
rect 37826 20040 37832 20052
rect 37476 20012 37832 20040
rect 34698 19864 34704 19916
rect 34756 19904 34762 19916
rect 35621 19907 35679 19913
rect 35621 19904 35633 19907
rect 34756 19876 35633 19904
rect 34756 19864 34762 19876
rect 35621 19873 35633 19876
rect 35667 19873 35679 19907
rect 37384 19904 37412 20000
rect 37476 19913 37504 20012
rect 37826 20000 37832 20012
rect 37884 20040 37890 20052
rect 40218 20040 40224 20052
rect 37884 20012 40224 20040
rect 37884 20000 37890 20012
rect 38654 19932 38660 19984
rect 38712 19932 38718 19984
rect 38838 19932 38844 19984
rect 38896 19932 38902 19984
rect 35621 19867 35679 19873
rect 37108 19876 37412 19904
rect 37461 19907 37519 19913
rect 34425 19839 34483 19845
rect 34425 19805 34437 19839
rect 34471 19805 34483 19839
rect 34425 19799 34483 19805
rect 34606 19796 34612 19848
rect 34664 19836 34670 19848
rect 37108 19845 37136 19876
rect 37461 19873 37473 19907
rect 37507 19873 37519 19907
rect 37461 19867 37519 19873
rect 34977 19839 35035 19845
rect 34977 19836 34989 19839
rect 34664 19808 34989 19836
rect 34664 19796 34670 19808
rect 34977 19805 34989 19808
rect 35023 19805 35035 19839
rect 34977 19799 35035 19805
rect 37093 19839 37151 19845
rect 37093 19805 37105 19839
rect 37139 19805 37151 19839
rect 37093 19799 37151 19805
rect 37182 19796 37188 19848
rect 37240 19836 37246 19848
rect 38672 19836 38700 19932
rect 39868 19913 39896 20012
rect 40218 20000 40224 20012
rect 40276 20000 40282 20052
rect 41417 20043 41475 20049
rect 41417 20009 41429 20043
rect 41463 20040 41475 20043
rect 41506 20040 41512 20052
rect 41463 20012 41512 20040
rect 41463 20009 41475 20012
rect 41417 20003 41475 20009
rect 41506 20000 41512 20012
rect 41564 20000 41570 20052
rect 42429 20043 42487 20049
rect 42429 20009 42441 20043
rect 42475 20040 42487 20043
rect 42794 20040 42800 20052
rect 42475 20012 42800 20040
rect 42475 20009 42487 20012
rect 42429 20003 42487 20009
rect 42794 20000 42800 20012
rect 42852 20000 42858 20052
rect 43530 20000 43536 20052
rect 43588 20000 43594 20052
rect 46658 20000 46664 20052
rect 46716 20040 46722 20052
rect 48498 20040 48504 20052
rect 46716 20012 48504 20040
rect 46716 20000 46722 20012
rect 40862 19932 40868 19984
rect 40920 19972 40926 19984
rect 40920 19944 41414 19972
rect 40920 19932 40926 19944
rect 39853 19907 39911 19913
rect 39853 19873 39865 19907
rect 39899 19873 39911 19907
rect 41386 19904 41414 19944
rect 43438 19932 43444 19984
rect 43496 19972 43502 19984
rect 44729 19975 44787 19981
rect 44729 19972 44741 19975
rect 43496 19944 44741 19972
rect 43496 19932 43502 19944
rect 44729 19941 44741 19944
rect 44775 19941 44787 19975
rect 44729 19935 44787 19941
rect 46753 19975 46811 19981
rect 46753 19941 46765 19975
rect 46799 19972 46811 19975
rect 47486 19972 47492 19984
rect 46799 19944 47492 19972
rect 46799 19941 46811 19944
rect 46753 19935 46811 19941
rect 47486 19932 47492 19944
rect 47544 19932 47550 19984
rect 44174 19904 44180 19916
rect 41386 19876 44180 19904
rect 39853 19867 39911 19873
rect 39209 19839 39267 19845
rect 39209 19836 39221 19839
rect 37240 19808 37872 19836
rect 38672 19808 39221 19836
rect 37240 19796 37246 19808
rect 29549 19771 29607 19777
rect 29549 19768 29561 19771
rect 28684 19740 29561 19768
rect 28684 19728 28690 19740
rect 29549 19737 29561 19740
rect 29595 19737 29607 19771
rect 34514 19768 34520 19780
rect 29549 19731 29607 19737
rect 29656 19740 34520 19768
rect 26970 19660 26976 19712
rect 27028 19660 27034 19712
rect 27430 19660 27436 19712
rect 27488 19700 27494 19712
rect 27798 19700 27804 19712
rect 27488 19672 27804 19700
rect 27488 19660 27494 19672
rect 27798 19660 27804 19672
rect 27856 19700 27862 19712
rect 28261 19703 28319 19709
rect 28261 19700 28273 19703
rect 27856 19672 28273 19700
rect 27856 19660 27862 19672
rect 28261 19669 28273 19672
rect 28307 19669 28319 19703
rect 28460 19700 28488 19728
rect 29656 19700 29684 19740
rect 34514 19728 34520 19740
rect 34572 19728 34578 19780
rect 35888 19771 35946 19777
rect 35888 19737 35900 19771
rect 35934 19768 35946 19771
rect 36630 19768 36636 19780
rect 35934 19740 36636 19768
rect 35934 19737 35946 19740
rect 35888 19731 35946 19737
rect 36630 19728 36636 19740
rect 36688 19728 36694 19780
rect 37274 19728 37280 19780
rect 37332 19768 37338 19780
rect 37369 19771 37427 19777
rect 37369 19768 37381 19771
rect 37332 19740 37381 19768
rect 37332 19728 37338 19740
rect 37369 19737 37381 19740
rect 37415 19737 37427 19771
rect 37706 19771 37764 19777
rect 37706 19768 37718 19771
rect 37369 19731 37427 19737
rect 37476 19740 37718 19768
rect 28460 19672 29684 19700
rect 28261 19663 28319 19669
rect 29730 19660 29736 19712
rect 29788 19709 29794 19712
rect 29788 19703 29807 19709
rect 29795 19669 29807 19703
rect 29788 19663 29807 19669
rect 29788 19660 29794 19663
rect 29914 19660 29920 19712
rect 29972 19660 29978 19712
rect 32401 19703 32459 19709
rect 32401 19669 32413 19703
rect 32447 19700 32459 19703
rect 33778 19700 33784 19712
rect 32447 19672 33784 19700
rect 32447 19669 32459 19672
rect 32401 19663 32459 19669
rect 33778 19660 33784 19672
rect 33836 19660 33842 19712
rect 34790 19660 34796 19712
rect 34848 19660 34854 19712
rect 36722 19660 36728 19712
rect 36780 19700 36786 19712
rect 36998 19700 37004 19712
rect 36780 19672 37004 19700
rect 36780 19660 36786 19672
rect 36998 19660 37004 19672
rect 37056 19660 37062 19712
rect 37093 19703 37151 19709
rect 37093 19669 37105 19703
rect 37139 19700 37151 19703
rect 37476 19700 37504 19740
rect 37706 19737 37718 19740
rect 37752 19737 37764 19771
rect 37844 19768 37872 19808
rect 39209 19805 39221 19808
rect 39255 19805 39267 19839
rect 39209 19799 39267 19805
rect 40120 19839 40178 19845
rect 40120 19805 40132 19839
rect 40166 19836 40178 19839
rect 40678 19836 40684 19848
rect 40166 19808 40684 19836
rect 40166 19805 40178 19808
rect 40120 19799 40178 19805
rect 40678 19796 40684 19808
rect 40736 19796 40742 19848
rect 41325 19839 41383 19845
rect 41325 19836 41337 19839
rect 41248 19808 41337 19836
rect 38378 19768 38384 19780
rect 37844 19740 38384 19768
rect 37706 19731 37764 19737
rect 38378 19728 38384 19740
rect 38436 19768 38442 19780
rect 39393 19771 39451 19777
rect 39393 19768 39405 19771
rect 38436 19740 39405 19768
rect 38436 19728 38442 19740
rect 39393 19737 39405 19740
rect 39439 19737 39451 19771
rect 39393 19731 39451 19737
rect 37139 19672 37504 19700
rect 37139 19669 37151 19672
rect 37093 19663 37151 19669
rect 40310 19660 40316 19712
rect 40368 19700 40374 19712
rect 41248 19709 41276 19808
rect 41325 19805 41337 19808
rect 41371 19805 41383 19839
rect 41325 19799 41383 19805
rect 42610 19796 42616 19848
rect 42668 19796 42674 19848
rect 43456 19845 43484 19876
rect 44174 19864 44180 19876
rect 44232 19864 44238 19916
rect 46014 19864 46020 19916
rect 46072 19904 46078 19916
rect 46477 19907 46535 19913
rect 46477 19904 46489 19907
rect 46072 19876 46489 19904
rect 46072 19864 46078 19876
rect 46477 19873 46489 19876
rect 46523 19873 46535 19907
rect 46477 19867 46535 19873
rect 46845 19907 46903 19913
rect 46845 19873 46857 19907
rect 46891 19904 46903 19907
rect 47581 19907 47639 19913
rect 47581 19904 47593 19907
rect 46891 19876 47593 19904
rect 46891 19873 46903 19876
rect 46845 19867 46903 19873
rect 47581 19873 47593 19876
rect 47627 19873 47639 19907
rect 47581 19867 47639 19873
rect 43441 19839 43499 19845
rect 43441 19805 43453 19839
rect 43487 19805 43499 19839
rect 44545 19839 44603 19845
rect 44545 19836 44557 19839
rect 43441 19799 43499 19805
rect 44284 19808 44557 19836
rect 41233 19703 41291 19709
rect 41233 19700 41245 19703
rect 40368 19672 41245 19700
rect 40368 19660 40374 19672
rect 41233 19669 41245 19672
rect 41279 19669 41291 19703
rect 44284 19700 44312 19808
rect 44545 19805 44557 19808
rect 44591 19805 44603 19839
rect 44545 19799 44603 19805
rect 44818 19796 44824 19848
rect 44876 19796 44882 19848
rect 45005 19839 45063 19845
rect 45005 19805 45017 19839
rect 45051 19836 45063 19839
rect 45051 19808 46612 19836
rect 45051 19805 45063 19808
rect 45005 19799 45063 19805
rect 44361 19771 44419 19777
rect 44361 19737 44373 19771
rect 44407 19768 44419 19771
rect 45250 19771 45308 19777
rect 45250 19768 45262 19771
rect 44407 19740 45262 19768
rect 44407 19737 44419 19740
rect 44361 19731 44419 19737
rect 45250 19737 45262 19740
rect 45296 19737 45308 19771
rect 45250 19731 45308 19737
rect 46474 19728 46480 19780
rect 46532 19728 46538 19780
rect 46584 19768 46612 19808
rect 46658 19796 46664 19848
rect 46716 19796 46722 19848
rect 46937 19839 46995 19845
rect 46937 19805 46949 19839
rect 46983 19836 46995 19839
rect 47026 19836 47032 19848
rect 46983 19808 47032 19836
rect 46983 19805 46995 19808
rect 46937 19799 46995 19805
rect 47026 19796 47032 19808
rect 47084 19796 47090 19848
rect 47118 19796 47124 19848
rect 47176 19796 47182 19848
rect 47688 19845 47716 20012
rect 48498 20000 48504 20012
rect 48556 20040 48562 20052
rect 49970 20040 49976 20052
rect 48556 20012 49976 20040
rect 48556 20000 48562 20012
rect 49970 20000 49976 20012
rect 50028 20040 50034 20052
rect 50522 20040 50528 20052
rect 50028 20012 50528 20040
rect 50028 20000 50034 20012
rect 50522 20000 50528 20012
rect 50580 20000 50586 20052
rect 48225 19975 48283 19981
rect 48225 19941 48237 19975
rect 48271 19972 48283 19975
rect 48314 19972 48320 19984
rect 48271 19944 48320 19972
rect 48271 19941 48283 19944
rect 48225 19935 48283 19941
rect 48314 19932 48320 19944
rect 48372 19932 48378 19984
rect 47857 19907 47915 19913
rect 47857 19873 47869 19907
rect 47903 19904 47915 19907
rect 47946 19904 47952 19916
rect 47903 19876 47952 19904
rect 47903 19873 47915 19876
rect 47857 19867 47915 19873
rect 47946 19864 47952 19876
rect 48004 19864 48010 19916
rect 49329 19907 49387 19913
rect 49329 19873 49341 19907
rect 49375 19904 49387 19907
rect 50433 19907 50491 19913
rect 50433 19904 50445 19907
rect 49375 19876 50445 19904
rect 49375 19873 49387 19876
rect 49329 19867 49387 19873
rect 50433 19873 50445 19876
rect 50479 19873 50491 19907
rect 50433 19867 50491 19873
rect 50522 19864 50528 19916
rect 50580 19904 50586 19916
rect 52181 19907 52239 19913
rect 52181 19904 52193 19907
rect 50580 19876 52193 19904
rect 50580 19864 50586 19876
rect 52181 19873 52193 19876
rect 52227 19873 52239 19907
rect 52181 19867 52239 19873
rect 47489 19839 47547 19845
rect 47489 19805 47501 19839
rect 47535 19805 47547 19839
rect 47489 19799 47547 19805
rect 47673 19839 47731 19845
rect 47673 19805 47685 19839
rect 47719 19805 47731 19839
rect 47673 19799 47731 19805
rect 49513 19839 49571 19845
rect 49513 19805 49525 19839
rect 49559 19805 49571 19839
rect 49513 19799 49571 19805
rect 47394 19768 47400 19780
rect 46584 19740 47400 19768
rect 47394 19728 47400 19740
rect 47452 19728 47458 19780
rect 45462 19700 45468 19712
rect 44284 19672 45468 19700
rect 41233 19663 41291 19669
rect 45462 19660 45468 19672
rect 45520 19660 45526 19712
rect 46382 19660 46388 19712
rect 46440 19660 46446 19712
rect 46492 19700 46520 19728
rect 47504 19700 47532 19799
rect 48317 19703 48375 19709
rect 48317 19700 48329 19703
rect 46492 19672 48329 19700
rect 48317 19669 48329 19672
rect 48363 19669 48375 19703
rect 49528 19700 49556 19799
rect 49602 19796 49608 19848
rect 49660 19796 49666 19848
rect 49970 19796 49976 19848
rect 50028 19796 50034 19848
rect 50062 19796 50068 19848
rect 50120 19836 50126 19848
rect 50157 19839 50215 19845
rect 50157 19836 50169 19839
rect 50120 19808 50169 19836
rect 50120 19796 50126 19808
rect 50157 19805 50169 19808
rect 50203 19805 50215 19839
rect 50157 19799 50215 19805
rect 68462 19796 68468 19848
rect 68520 19796 68526 19848
rect 49694 19728 49700 19780
rect 49752 19728 49758 19780
rect 49786 19728 49792 19780
rect 49844 19777 49850 19780
rect 49844 19771 49893 19777
rect 49844 19737 49847 19771
rect 49881 19768 49893 19771
rect 49881 19740 50660 19768
rect 49881 19737 49893 19740
rect 49844 19731 49893 19737
rect 49844 19728 49850 19731
rect 50632 19712 50660 19740
rect 51074 19728 51080 19780
rect 51132 19728 51138 19780
rect 50154 19700 50160 19712
rect 49528 19672 50160 19700
rect 48317 19663 48375 19669
rect 50154 19660 50160 19672
rect 50212 19660 50218 19712
rect 50614 19660 50620 19712
rect 50672 19660 50678 19712
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 26970 19456 26976 19508
rect 27028 19456 27034 19508
rect 27617 19499 27675 19505
rect 27617 19496 27629 19499
rect 27080 19468 27629 19496
rect 26988 19369 27016 19456
rect 26145 19363 26203 19369
rect 26145 19329 26157 19363
rect 26191 19360 26203 19363
rect 26973 19363 27031 19369
rect 26191 19332 26924 19360
rect 26191 19329 26203 19332
rect 26145 19323 26203 19329
rect 26896 19292 26924 19332
rect 26973 19329 26985 19363
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 27080 19292 27108 19468
rect 27617 19465 27629 19468
rect 27663 19465 27675 19499
rect 27617 19459 27675 19465
rect 27706 19456 27712 19508
rect 27764 19456 27770 19508
rect 28997 19499 29055 19505
rect 28997 19465 29009 19499
rect 29043 19496 29055 19499
rect 29086 19496 29092 19508
rect 29043 19468 29092 19496
rect 29043 19465 29055 19468
rect 28997 19459 29055 19465
rect 29086 19456 29092 19468
rect 29144 19456 29150 19508
rect 32950 19496 32956 19508
rect 31864 19468 32956 19496
rect 27724 19428 27752 19456
rect 31864 19440 31892 19468
rect 32950 19456 32956 19468
rect 33008 19456 33014 19508
rect 33502 19456 33508 19508
rect 33560 19496 33566 19508
rect 33781 19499 33839 19505
rect 33781 19496 33793 19499
rect 33560 19468 33793 19496
rect 33560 19456 33566 19468
rect 33781 19465 33793 19468
rect 33827 19496 33839 19499
rect 34054 19496 34060 19508
rect 33827 19468 34060 19496
rect 33827 19465 33839 19468
rect 33781 19459 33839 19465
rect 34054 19456 34060 19468
rect 34112 19456 34118 19508
rect 34790 19456 34796 19508
rect 34848 19456 34854 19508
rect 35621 19499 35679 19505
rect 35621 19465 35633 19499
rect 35667 19465 35679 19499
rect 35621 19459 35679 19465
rect 27724 19400 31524 19428
rect 27249 19363 27307 19369
rect 27249 19329 27261 19363
rect 27295 19329 27307 19363
rect 27249 19323 27307 19329
rect 26896 19264 27108 19292
rect 27264 19224 27292 19323
rect 27338 19320 27344 19372
rect 27396 19320 27402 19372
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19360 27491 19363
rect 27724 19360 27752 19400
rect 31496 19372 31524 19400
rect 31846 19388 31852 19440
rect 31904 19388 31910 19440
rect 32214 19388 32220 19440
rect 32272 19428 32278 19440
rect 33594 19428 33600 19440
rect 32272 19400 33600 19428
rect 32272 19388 32278 19400
rect 33594 19388 33600 19400
rect 33652 19388 33658 19440
rect 33962 19428 33968 19440
rect 33704 19400 33968 19428
rect 33704 19372 33732 19400
rect 33962 19388 33968 19400
rect 34020 19388 34026 19440
rect 34508 19431 34566 19437
rect 34072 19400 34376 19428
rect 34072 19372 34100 19400
rect 27479 19332 27752 19360
rect 27479 19329 27491 19332
rect 27433 19323 27491 19329
rect 27798 19320 27804 19372
rect 27856 19360 27862 19372
rect 27893 19363 27951 19369
rect 27893 19360 27905 19363
rect 27856 19332 27905 19360
rect 27856 19320 27862 19332
rect 27893 19329 27905 19332
rect 27939 19329 27951 19363
rect 27893 19323 27951 19329
rect 27985 19363 28043 19369
rect 27985 19329 27997 19363
rect 28031 19329 28043 19363
rect 27985 19323 28043 19329
rect 28077 19363 28135 19369
rect 28077 19329 28089 19363
rect 28123 19329 28135 19363
rect 28077 19323 28135 19329
rect 28537 19363 28595 19369
rect 28537 19329 28549 19363
rect 28583 19360 28595 19363
rect 28626 19360 28632 19372
rect 28583 19332 28632 19360
rect 28583 19329 28595 19332
rect 28537 19323 28595 19329
rect 27356 19292 27384 19320
rect 28000 19292 28028 19323
rect 27356 19264 28028 19292
rect 28092 19292 28120 19323
rect 28626 19320 28632 19332
rect 28684 19320 28690 19372
rect 28718 19320 28724 19372
rect 28776 19320 28782 19372
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19360 29239 19363
rect 29914 19360 29920 19372
rect 29227 19332 29920 19360
rect 29227 19329 29239 19332
rect 29181 19323 29239 19329
rect 29914 19320 29920 19332
rect 29972 19320 29978 19372
rect 31478 19320 31484 19372
rect 31536 19320 31542 19372
rect 31570 19320 31576 19372
rect 31628 19320 31634 19372
rect 31754 19320 31760 19372
rect 31812 19360 31818 19372
rect 32125 19363 32183 19369
rect 32125 19360 32137 19363
rect 31812 19332 32137 19360
rect 31812 19320 31818 19332
rect 32125 19329 32137 19332
rect 32171 19329 32183 19363
rect 32381 19363 32439 19369
rect 32381 19360 32393 19363
rect 32125 19323 32183 19329
rect 32232 19332 32393 19360
rect 28813 19295 28871 19301
rect 28813 19292 28825 19295
rect 28092 19264 28825 19292
rect 28813 19261 28825 19264
rect 28859 19292 28871 19295
rect 28902 19292 28908 19304
rect 28859 19264 28908 19292
rect 28859 19261 28871 19264
rect 28813 19255 28871 19261
rect 28902 19252 28908 19264
rect 28960 19252 28966 19304
rect 32232 19292 32260 19332
rect 32381 19329 32393 19332
rect 32427 19329 32439 19363
rect 32381 19323 32439 19329
rect 33686 19320 33692 19372
rect 33744 19320 33750 19372
rect 33873 19363 33931 19369
rect 33873 19329 33885 19363
rect 33919 19360 33931 19363
rect 34054 19360 34060 19372
rect 33919 19332 34060 19360
rect 33919 19329 33931 19332
rect 33873 19323 33931 19329
rect 34054 19320 34060 19332
rect 34112 19320 34118 19372
rect 34241 19363 34299 19369
rect 34241 19329 34253 19363
rect 34287 19329 34299 19363
rect 34348 19360 34376 19400
rect 34508 19397 34520 19431
rect 34554 19428 34566 19431
rect 34808 19428 34836 19456
rect 34554 19400 34836 19428
rect 34554 19397 34566 19400
rect 34508 19391 34566 19397
rect 35636 19360 35664 19459
rect 36630 19456 36636 19508
rect 36688 19456 36694 19508
rect 40494 19456 40500 19508
rect 40552 19496 40558 19508
rect 40552 19468 42196 19496
rect 40552 19456 40558 19468
rect 40512 19428 40540 19456
rect 34348 19332 35664 19360
rect 37660 19400 40540 19428
rect 34241 19323 34299 19329
rect 31588 19264 31800 19292
rect 27614 19224 27620 19236
rect 27264 19196 27620 19224
rect 27614 19184 27620 19196
rect 27672 19184 27678 19236
rect 27709 19227 27767 19233
rect 27709 19193 27721 19227
rect 27755 19224 27767 19227
rect 28626 19224 28632 19236
rect 27755 19196 28632 19224
rect 27755 19193 27767 19196
rect 27709 19187 27767 19193
rect 28626 19184 28632 19196
rect 28684 19184 28690 19236
rect 31588 19233 31616 19264
rect 31573 19227 31631 19233
rect 31573 19193 31585 19227
rect 31619 19193 31631 19227
rect 31573 19187 31631 19193
rect 31665 19227 31723 19233
rect 31665 19193 31677 19227
rect 31711 19193 31723 19227
rect 31772 19224 31800 19264
rect 31956 19264 32260 19292
rect 31956 19224 31984 19264
rect 31772 19196 31984 19224
rect 31665 19187 31723 19193
rect 26234 19116 26240 19168
rect 26292 19116 26298 19168
rect 27430 19116 27436 19168
rect 27488 19116 27494 19168
rect 27632 19156 27660 19184
rect 28261 19159 28319 19165
rect 28261 19156 28273 19159
rect 27632 19128 28273 19156
rect 28261 19125 28273 19128
rect 28307 19125 28319 19159
rect 28261 19119 28319 19125
rect 28350 19116 28356 19168
rect 28408 19116 28414 19168
rect 31680 19156 31708 19187
rect 33318 19184 33324 19236
rect 33376 19224 33382 19236
rect 33505 19227 33563 19233
rect 33505 19224 33517 19227
rect 33376 19196 33517 19224
rect 33376 19184 33382 19196
rect 33505 19193 33517 19196
rect 33551 19224 33563 19227
rect 33597 19227 33655 19233
rect 33597 19224 33609 19227
rect 33551 19196 33609 19224
rect 33551 19193 33563 19196
rect 33505 19187 33563 19193
rect 33597 19193 33609 19196
rect 33643 19193 33655 19227
rect 33597 19187 33655 19193
rect 32858 19156 32864 19168
rect 31680 19128 32864 19156
rect 32858 19116 32864 19128
rect 32916 19116 32922 19168
rect 34146 19116 34152 19168
rect 34204 19116 34210 19168
rect 34256 19156 34284 19323
rect 36078 19252 36084 19304
rect 36136 19252 36142 19304
rect 36906 19252 36912 19304
rect 36964 19292 36970 19304
rect 37277 19295 37335 19301
rect 37277 19292 37289 19295
rect 36964 19264 37289 19292
rect 36964 19252 36970 19264
rect 37277 19261 37289 19264
rect 37323 19261 37335 19295
rect 37277 19255 37335 19261
rect 37458 19252 37464 19304
rect 37516 19292 37522 19304
rect 37660 19292 37688 19400
rect 41230 19388 41236 19440
rect 41288 19428 41294 19440
rect 42061 19431 42119 19437
rect 42061 19428 42073 19431
rect 41288 19400 42073 19428
rect 41288 19388 41294 19400
rect 42061 19397 42073 19400
rect 42107 19397 42119 19431
rect 42168 19428 42196 19468
rect 42610 19456 42616 19508
rect 42668 19496 42674 19508
rect 42981 19499 43039 19505
rect 42981 19496 42993 19499
rect 42668 19468 42993 19496
rect 42668 19456 42674 19468
rect 42981 19465 42993 19468
rect 43027 19465 43039 19499
rect 42981 19459 43039 19465
rect 44450 19456 44456 19508
rect 44508 19456 44514 19508
rect 44818 19456 44824 19508
rect 44876 19496 44882 19508
rect 46017 19499 46075 19505
rect 46017 19496 46029 19499
rect 44876 19468 46029 19496
rect 44876 19456 44882 19468
rect 46017 19465 46029 19468
rect 46063 19465 46075 19499
rect 46017 19459 46075 19465
rect 46658 19456 46664 19508
rect 46716 19496 46722 19508
rect 46753 19499 46811 19505
rect 46753 19496 46765 19499
rect 46716 19468 46765 19496
rect 46716 19456 46722 19468
rect 46753 19465 46765 19468
rect 46799 19465 46811 19499
rect 46753 19459 46811 19465
rect 47026 19456 47032 19508
rect 47084 19456 47090 19508
rect 47302 19456 47308 19508
rect 47360 19496 47366 19508
rect 47360 19468 47624 19496
rect 47360 19456 47366 19468
rect 42705 19431 42763 19437
rect 42705 19428 42717 19431
rect 42168 19400 42717 19428
rect 42061 19391 42119 19397
rect 42705 19397 42717 19400
rect 42751 19397 42763 19431
rect 43438 19428 43444 19440
rect 42705 19391 42763 19397
rect 43272 19400 43444 19428
rect 39669 19363 39727 19369
rect 39669 19329 39681 19363
rect 39715 19360 39727 19363
rect 39850 19360 39856 19372
rect 39715 19332 39856 19360
rect 39715 19329 39727 19332
rect 39669 19323 39727 19329
rect 39850 19320 39856 19332
rect 39908 19320 39914 19372
rect 40402 19320 40408 19372
rect 40460 19360 40466 19372
rect 40862 19360 40868 19372
rect 40460 19332 40868 19360
rect 40460 19320 40466 19332
rect 40862 19320 40868 19332
rect 40920 19320 40926 19372
rect 41322 19320 41328 19372
rect 41380 19320 41386 19372
rect 42429 19363 42487 19369
rect 42429 19329 42441 19363
rect 42475 19360 42487 19363
rect 43272 19360 43300 19400
rect 43438 19388 43444 19400
rect 43496 19388 43502 19440
rect 43622 19388 43628 19440
rect 43680 19428 43686 19440
rect 43901 19431 43959 19437
rect 43901 19428 43913 19431
rect 43680 19400 43913 19428
rect 43680 19388 43686 19400
rect 43901 19397 43913 19400
rect 43947 19397 43959 19431
rect 43901 19391 43959 19397
rect 42475 19332 43300 19360
rect 43349 19363 43407 19369
rect 42475 19329 42487 19332
rect 42429 19323 42487 19329
rect 43349 19329 43361 19363
rect 43395 19360 43407 19363
rect 43714 19360 43720 19372
rect 43395 19332 43720 19360
rect 43395 19329 43407 19332
rect 43349 19323 43407 19329
rect 43714 19320 43720 19332
rect 43772 19320 43778 19372
rect 43809 19363 43867 19369
rect 43809 19329 43821 19363
rect 43855 19334 43867 19363
rect 43993 19363 44051 19369
rect 43855 19329 43944 19334
rect 43809 19323 43944 19329
rect 43993 19329 44005 19363
rect 44039 19360 44051 19363
rect 44468 19360 44496 19456
rect 46293 19363 46351 19369
rect 44039 19332 44496 19360
rect 46032 19332 46244 19360
rect 44039 19329 44051 19332
rect 43993 19323 44051 19329
rect 43824 19306 43944 19323
rect 37516 19264 37688 19292
rect 37516 19252 37522 19264
rect 42518 19252 42524 19304
rect 42576 19292 42582 19304
rect 43441 19295 43499 19301
rect 43441 19292 43453 19295
rect 42576 19264 43453 19292
rect 42576 19252 42582 19264
rect 43441 19261 43453 19264
rect 43487 19261 43499 19295
rect 43441 19255 43499 19261
rect 43530 19252 43536 19304
rect 43588 19252 43594 19304
rect 43916 19292 43944 19306
rect 44082 19292 44088 19304
rect 43916 19264 44088 19292
rect 44082 19252 44088 19264
rect 44140 19252 44146 19304
rect 45465 19295 45523 19301
rect 45465 19261 45477 19295
rect 45511 19292 45523 19295
rect 46032 19292 46060 19332
rect 45511 19264 46060 19292
rect 46109 19295 46167 19301
rect 45511 19261 45523 19264
rect 45465 19255 45523 19261
rect 46109 19261 46121 19295
rect 46155 19261 46167 19295
rect 46216 19292 46244 19332
rect 46293 19329 46305 19363
rect 46339 19360 46351 19363
rect 46842 19360 46848 19372
rect 46339 19332 46848 19360
rect 46339 19329 46351 19332
rect 46293 19323 46351 19329
rect 46584 19304 46612 19332
rect 46842 19320 46848 19332
rect 46900 19320 46906 19372
rect 46934 19320 46940 19372
rect 46992 19320 46998 19372
rect 47044 19369 47072 19456
rect 47596 19437 47624 19468
rect 50154 19456 50160 19508
rect 50212 19456 50218 19508
rect 47581 19431 47639 19437
rect 47581 19397 47593 19431
rect 47627 19397 47639 19431
rect 48774 19428 48780 19440
rect 47581 19391 47639 19397
rect 47780 19400 48780 19428
rect 47780 19372 47808 19400
rect 48774 19388 48780 19400
rect 48832 19428 48838 19440
rect 50525 19431 50583 19437
rect 50525 19428 50537 19431
rect 48832 19400 50537 19428
rect 48832 19388 48838 19400
rect 50525 19397 50537 19400
rect 50571 19397 50583 19431
rect 50525 19391 50583 19397
rect 47029 19363 47087 19369
rect 47029 19329 47041 19363
rect 47075 19329 47087 19363
rect 47029 19323 47087 19329
rect 47302 19320 47308 19372
rect 47360 19320 47366 19372
rect 47762 19320 47768 19372
rect 47820 19320 47826 19372
rect 49786 19320 49792 19372
rect 49844 19320 49850 19372
rect 49970 19320 49976 19372
rect 50028 19360 50034 19372
rect 50341 19363 50399 19369
rect 50341 19360 50353 19363
rect 50028 19332 50353 19360
rect 50028 19320 50034 19332
rect 50341 19329 50353 19332
rect 50387 19329 50399 19363
rect 50341 19323 50399 19329
rect 50617 19363 50675 19369
rect 50617 19329 50629 19363
rect 50663 19360 50675 19363
rect 50663 19332 50844 19360
rect 50663 19329 50675 19332
rect 50617 19323 50675 19329
rect 46382 19292 46388 19304
rect 46216 19264 46388 19292
rect 46109 19255 46167 19261
rect 36354 19184 36360 19236
rect 36412 19224 36418 19236
rect 36412 19196 38332 19224
rect 36412 19184 36418 19196
rect 38304 19168 38332 19196
rect 44266 19184 44272 19236
rect 44324 19224 44330 19236
rect 46124 19224 46152 19255
rect 46382 19252 46388 19264
rect 46440 19252 46446 19304
rect 46566 19252 46572 19304
rect 46624 19252 46630 19304
rect 44324 19196 46152 19224
rect 44324 19184 44330 19196
rect 46198 19184 46204 19236
rect 46256 19224 46262 19236
rect 46477 19227 46535 19233
rect 46477 19224 46489 19227
rect 46256 19196 46489 19224
rect 46256 19184 46262 19196
rect 46477 19193 46489 19196
rect 46523 19224 46535 19227
rect 49804 19224 49832 19320
rect 50816 19304 50844 19332
rect 50798 19252 50804 19304
rect 50856 19252 50862 19304
rect 46523 19196 49832 19224
rect 46523 19193 46535 19196
rect 46477 19187 46535 19193
rect 35342 19156 35348 19168
rect 34256 19128 35348 19156
rect 35342 19116 35348 19128
rect 35400 19116 35406 19168
rect 36170 19116 36176 19168
rect 36228 19156 36234 19168
rect 37921 19159 37979 19165
rect 37921 19156 37933 19159
rect 36228 19128 37933 19156
rect 36228 19116 36234 19128
rect 37921 19125 37933 19128
rect 37967 19125 37979 19159
rect 37921 19119 37979 19125
rect 38286 19116 38292 19168
rect 38344 19116 38350 19168
rect 39758 19116 39764 19168
rect 39816 19116 39822 19168
rect 42610 19116 42616 19168
rect 42668 19116 42674 19168
rect 43530 19116 43536 19168
rect 43588 19156 43594 19168
rect 44284 19156 44312 19184
rect 47412 19168 47440 19196
rect 43588 19128 44312 19156
rect 43588 19116 43594 19128
rect 47210 19116 47216 19168
rect 47268 19116 47274 19168
rect 47394 19116 47400 19168
rect 47452 19116 47458 19168
rect 47946 19116 47952 19168
rect 48004 19116 48010 19168
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 27246 18912 27252 18964
rect 27304 18952 27310 18964
rect 27433 18955 27491 18961
rect 27433 18952 27445 18955
rect 27304 18924 27445 18952
rect 27304 18912 27310 18924
rect 27433 18921 27445 18924
rect 27479 18921 27491 18955
rect 27433 18915 27491 18921
rect 27617 18955 27675 18961
rect 27617 18921 27629 18955
rect 27663 18952 27675 18955
rect 28074 18952 28080 18964
rect 27663 18924 28080 18952
rect 27663 18921 27675 18924
rect 27617 18915 27675 18921
rect 28074 18912 28080 18924
rect 28132 18912 28138 18964
rect 31665 18955 31723 18961
rect 31665 18921 31677 18955
rect 31711 18952 31723 18955
rect 31846 18952 31852 18964
rect 31711 18924 31852 18952
rect 31711 18921 31723 18924
rect 31665 18915 31723 18921
rect 31846 18912 31852 18924
rect 31904 18912 31910 18964
rect 32858 18912 32864 18964
rect 32916 18912 32922 18964
rect 34054 18912 34060 18964
rect 34112 18952 34118 18964
rect 34149 18955 34207 18961
rect 34149 18952 34161 18955
rect 34112 18924 34161 18952
rect 34112 18912 34118 18924
rect 34149 18921 34161 18924
rect 34195 18921 34207 18955
rect 34149 18915 34207 18921
rect 34333 18955 34391 18961
rect 34333 18921 34345 18955
rect 34379 18952 34391 18955
rect 34606 18952 34612 18964
rect 34379 18924 34612 18952
rect 34379 18921 34391 18924
rect 34333 18915 34391 18921
rect 34606 18912 34612 18924
rect 34664 18912 34670 18964
rect 36078 18912 36084 18964
rect 36136 18952 36142 18964
rect 36633 18955 36691 18961
rect 36633 18952 36645 18955
rect 36136 18924 36645 18952
rect 36136 18912 36142 18924
rect 36633 18921 36645 18924
rect 36679 18921 36691 18955
rect 36633 18915 36691 18921
rect 36814 18912 36820 18964
rect 36872 18912 36878 18964
rect 41138 18912 41144 18964
rect 41196 18952 41202 18964
rect 43257 18955 43315 18961
rect 43257 18952 43269 18955
rect 41196 18924 43269 18952
rect 41196 18912 41202 18924
rect 43257 18921 43269 18924
rect 43303 18921 43315 18955
rect 43257 18915 43315 18921
rect 45002 18912 45008 18964
rect 45060 18952 45066 18964
rect 45925 18955 45983 18961
rect 45925 18952 45937 18955
rect 45060 18924 45937 18952
rect 45060 18912 45066 18924
rect 45925 18921 45937 18924
rect 45971 18921 45983 18955
rect 45925 18915 45983 18921
rect 46106 18912 46112 18964
rect 46164 18912 46170 18964
rect 46382 18912 46388 18964
rect 46440 18952 46446 18964
rect 46440 18924 47164 18952
rect 46440 18912 46446 18924
rect 33318 18776 33324 18828
rect 33376 18776 33382 18828
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1581 18751 1639 18757
rect 1581 18748 1593 18751
rect 992 18720 1593 18748
rect 992 18708 998 18720
rect 1581 18717 1593 18720
rect 1627 18717 1639 18751
rect 1581 18711 1639 18717
rect 25222 18708 25228 18760
rect 25280 18748 25286 18760
rect 25593 18751 25651 18757
rect 25593 18748 25605 18751
rect 25280 18720 25605 18748
rect 25280 18708 25286 18720
rect 25593 18717 25605 18720
rect 25639 18717 25651 18751
rect 25593 18711 25651 18717
rect 25860 18751 25918 18757
rect 25860 18717 25872 18751
rect 25906 18748 25918 18751
rect 26234 18748 26240 18760
rect 25906 18720 26240 18748
rect 25906 18717 25918 18720
rect 25860 18711 25918 18717
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 27065 18751 27123 18757
rect 27065 18717 27077 18751
rect 27111 18748 27123 18751
rect 27154 18748 27160 18760
rect 27111 18720 27160 18748
rect 27111 18717 27123 18720
rect 27065 18711 27123 18717
rect 27154 18708 27160 18720
rect 27212 18748 27218 18760
rect 29549 18751 29607 18757
rect 27212 18720 28948 18748
rect 27212 18708 27218 18720
rect 28442 18640 28448 18692
rect 28500 18640 28506 18692
rect 28920 18624 28948 18720
rect 29549 18717 29561 18751
rect 29595 18717 29607 18751
rect 29549 18711 29607 18717
rect 29178 18640 29184 18692
rect 29236 18680 29242 18692
rect 29564 18680 29592 18711
rect 33134 18708 33140 18760
rect 33192 18748 33198 18760
rect 34072 18748 34100 18912
rect 36998 18844 37004 18896
rect 37056 18884 37062 18896
rect 39390 18884 39396 18896
rect 37056 18856 39396 18884
rect 37056 18844 37062 18856
rect 39390 18844 39396 18856
rect 39448 18884 39454 18896
rect 39758 18884 39764 18896
rect 39448 18856 39764 18884
rect 39448 18844 39454 18856
rect 39758 18844 39764 18856
rect 39816 18844 39822 18896
rect 42153 18887 42211 18893
rect 42153 18853 42165 18887
rect 42199 18884 42211 18887
rect 42199 18856 42656 18884
rect 42199 18853 42211 18856
rect 42153 18847 42211 18853
rect 36722 18816 36728 18828
rect 35268 18788 36728 18816
rect 33192 18720 34100 18748
rect 33192 18708 33198 18720
rect 34514 18708 34520 18760
rect 34572 18748 34578 18760
rect 34701 18751 34759 18757
rect 34701 18748 34713 18751
rect 34572 18720 34713 18748
rect 34572 18708 34578 18720
rect 34701 18717 34713 18720
rect 34747 18717 34759 18751
rect 34701 18711 34759 18717
rect 29236 18652 29592 18680
rect 29816 18683 29874 18689
rect 29236 18640 29242 18652
rect 29816 18649 29828 18683
rect 29862 18680 29874 18683
rect 30190 18680 30196 18692
rect 29862 18652 30196 18680
rect 29862 18649 29874 18652
rect 29816 18643 29874 18649
rect 30190 18640 30196 18652
rect 30248 18640 30254 18692
rect 31386 18640 31392 18692
rect 31444 18640 31450 18692
rect 32861 18683 32919 18689
rect 32861 18649 32873 18683
rect 32907 18680 32919 18683
rect 33873 18683 33931 18689
rect 33873 18680 33885 18683
rect 32907 18652 33885 18680
rect 32907 18649 32919 18652
rect 32861 18643 32919 18649
rect 33873 18649 33885 18652
rect 33919 18649 33931 18683
rect 33873 18643 33931 18649
rect 33962 18640 33968 18692
rect 34020 18680 34026 18692
rect 35268 18680 35296 18788
rect 36722 18776 36728 18788
rect 36780 18776 36786 18828
rect 38304 18788 38976 18816
rect 37077 18761 37135 18767
rect 36170 18757 36176 18760
rect 35989 18751 36047 18757
rect 35989 18717 36001 18751
rect 36035 18717 36047 18751
rect 35989 18711 36047 18717
rect 36137 18751 36176 18757
rect 36137 18717 36149 18751
rect 36137 18711 36176 18717
rect 34020 18652 35296 18680
rect 34020 18640 34026 18652
rect 35342 18640 35348 18692
rect 35400 18680 35406 18692
rect 35437 18683 35495 18689
rect 35437 18680 35449 18683
rect 35400 18652 35449 18680
rect 35400 18640 35406 18652
rect 35437 18649 35449 18652
rect 35483 18649 35495 18683
rect 36004 18680 36032 18711
rect 36170 18708 36176 18711
rect 36228 18708 36234 18760
rect 36262 18708 36268 18760
rect 36320 18708 36326 18760
rect 36354 18708 36360 18760
rect 36412 18708 36418 18760
rect 36446 18708 36452 18760
rect 36504 18757 36510 18760
rect 37077 18758 37089 18761
rect 37123 18760 37135 18761
rect 36504 18751 36553 18757
rect 36504 18717 36507 18751
rect 36541 18748 36553 18751
rect 36930 18748 37089 18758
rect 36541 18730 37089 18748
rect 36541 18720 36958 18730
rect 37077 18727 37089 18730
rect 37077 18721 37096 18727
rect 36541 18717 36553 18720
rect 36504 18711 36553 18717
rect 36504 18708 36510 18711
rect 37090 18708 37096 18721
rect 37148 18708 37154 18760
rect 37182 18708 37188 18760
rect 37240 18708 37246 18760
rect 37918 18708 37924 18760
rect 37976 18708 37982 18760
rect 38069 18751 38127 18757
rect 38069 18717 38081 18751
rect 38115 18748 38127 18751
rect 38304 18748 38332 18788
rect 38115 18720 38332 18748
rect 38115 18717 38127 18720
rect 38069 18711 38127 18717
rect 38378 18708 38384 18760
rect 38436 18757 38442 18760
rect 38948 18757 38976 18788
rect 42518 18776 42524 18828
rect 42576 18776 42582 18828
rect 42628 18825 42656 18856
rect 44192 18856 45984 18884
rect 42613 18819 42671 18825
rect 42613 18785 42625 18819
rect 42659 18816 42671 18819
rect 42659 18788 43760 18816
rect 42659 18785 42671 18788
rect 42613 18779 42671 18785
rect 38436 18748 38444 18757
rect 38933 18751 38991 18757
rect 38436 18720 38481 18748
rect 38436 18711 38444 18720
rect 38933 18717 38945 18751
rect 38979 18717 38991 18751
rect 38933 18711 38991 18717
rect 38436 18708 38442 18711
rect 36004 18652 36768 18680
rect 35437 18643 35495 18649
rect 36740 18624 36768 18652
rect 36814 18640 36820 18692
rect 36872 18640 36878 18692
rect 37200 18680 37228 18708
rect 37016 18652 37228 18680
rect 26973 18615 27031 18621
rect 26973 18581 26985 18615
rect 27019 18612 27031 18615
rect 27433 18615 27491 18621
rect 27433 18612 27445 18615
rect 27019 18584 27445 18612
rect 27019 18581 27031 18584
rect 26973 18575 27031 18581
rect 27433 18581 27445 18584
rect 27479 18612 27491 18615
rect 27522 18612 27528 18624
rect 27479 18584 27528 18612
rect 27479 18581 27491 18584
rect 27433 18575 27491 18581
rect 27522 18572 27528 18584
rect 27580 18572 27586 18624
rect 28902 18572 28908 18624
rect 28960 18612 28966 18624
rect 29546 18612 29552 18624
rect 28960 18584 29552 18612
rect 28960 18572 28966 18584
rect 29546 18572 29552 18584
rect 29604 18612 29610 18624
rect 30929 18615 30987 18621
rect 30929 18612 30941 18615
rect 29604 18584 30941 18612
rect 29604 18572 29610 18584
rect 30929 18581 30941 18584
rect 30975 18581 30987 18615
rect 30929 18575 30987 18581
rect 33045 18615 33103 18621
rect 33045 18581 33057 18615
rect 33091 18612 33103 18615
rect 33502 18612 33508 18624
rect 33091 18584 33508 18612
rect 33091 18581 33103 18584
rect 33045 18575 33103 18581
rect 33502 18572 33508 18584
rect 33560 18572 33566 18624
rect 33686 18572 33692 18624
rect 33744 18612 33750 18624
rect 34165 18615 34223 18621
rect 34165 18612 34177 18615
rect 33744 18584 34177 18612
rect 33744 18572 33750 18584
rect 34165 18581 34177 18584
rect 34211 18581 34223 18615
rect 34165 18575 34223 18581
rect 36722 18572 36728 18624
rect 36780 18572 36786 18624
rect 37016 18621 37044 18652
rect 38194 18640 38200 18692
rect 38252 18640 38258 18692
rect 38286 18640 38292 18692
rect 38344 18640 38350 18692
rect 38470 18640 38476 18692
rect 38528 18680 38534 18692
rect 38654 18680 38660 18692
rect 38528 18652 38660 18680
rect 38528 18640 38534 18652
rect 38654 18640 38660 18652
rect 38712 18640 38718 18692
rect 38948 18624 38976 18711
rect 40126 18708 40132 18760
rect 40184 18708 40190 18760
rect 40773 18751 40831 18757
rect 40773 18717 40785 18751
rect 40819 18748 40831 18751
rect 40819 18720 41276 18748
rect 40819 18717 40831 18720
rect 40773 18711 40831 18717
rect 41248 18692 41276 18720
rect 41046 18689 41052 18692
rect 41040 18643 41052 18689
rect 41046 18640 41052 18643
rect 41104 18640 41110 18692
rect 41230 18640 41236 18692
rect 41288 18640 41294 18692
rect 42536 18680 42564 18776
rect 43732 18760 43760 18788
rect 43806 18776 43812 18828
rect 43864 18816 43870 18828
rect 44192 18816 44220 18856
rect 43864 18788 44220 18816
rect 43864 18776 43870 18788
rect 43257 18751 43315 18757
rect 43257 18717 43269 18751
rect 43303 18748 43315 18751
rect 43438 18748 43444 18760
rect 43303 18720 43444 18748
rect 43303 18717 43315 18720
rect 43257 18711 43315 18717
rect 43438 18708 43444 18720
rect 43496 18708 43502 18760
rect 43533 18751 43591 18757
rect 43533 18717 43545 18751
rect 43579 18717 43591 18751
rect 43533 18711 43591 18717
rect 43548 18680 43576 18711
rect 43714 18708 43720 18760
rect 43772 18708 43778 18760
rect 43898 18708 43904 18760
rect 43956 18708 43962 18760
rect 44192 18757 44220 18788
rect 44269 18819 44327 18825
rect 44269 18785 44281 18819
rect 44315 18816 44327 18819
rect 45005 18819 45063 18825
rect 45005 18816 45017 18819
rect 44315 18788 45017 18816
rect 44315 18785 44327 18788
rect 44269 18779 44327 18785
rect 45005 18785 45017 18788
rect 45051 18785 45063 18819
rect 45005 18779 45063 18785
rect 44177 18751 44235 18757
rect 44177 18717 44189 18751
rect 44223 18717 44235 18751
rect 44177 18711 44235 18717
rect 44358 18708 44364 18760
rect 44416 18708 44422 18760
rect 44637 18751 44695 18757
rect 44637 18717 44649 18751
rect 44683 18717 44695 18751
rect 44637 18711 44695 18717
rect 44082 18680 44088 18692
rect 42536 18652 44088 18680
rect 44082 18640 44088 18652
rect 44140 18680 44146 18692
rect 44652 18680 44680 18711
rect 44140 18652 44680 18680
rect 44140 18640 44146 18652
rect 44818 18640 44824 18692
rect 44876 18680 44882 18692
rect 45956 18689 45984 18856
rect 46658 18844 46664 18896
rect 46716 18884 46722 18896
rect 47136 18884 47164 18924
rect 47210 18912 47216 18964
rect 47268 18952 47274 18964
rect 47397 18955 47455 18961
rect 47397 18952 47409 18955
rect 47268 18924 47409 18952
rect 47268 18912 47274 18924
rect 47397 18921 47409 18924
rect 47443 18921 47455 18955
rect 50798 18952 50804 18964
rect 47397 18915 47455 18921
rect 48700 18924 50804 18952
rect 46716 18856 46888 18884
rect 47136 18856 47256 18884
rect 46716 18844 46722 18856
rect 46860 18825 46888 18856
rect 46845 18819 46903 18825
rect 46845 18785 46857 18819
rect 46891 18785 46903 18819
rect 47228 18816 47256 18856
rect 47228 18788 47348 18816
rect 46845 18779 46903 18785
rect 46293 18751 46351 18757
rect 46293 18717 46305 18751
rect 46339 18748 46351 18751
rect 46750 18748 46756 18760
rect 46339 18720 46756 18748
rect 46339 18717 46351 18720
rect 46293 18711 46351 18717
rect 46750 18708 46756 18720
rect 46808 18708 46814 18760
rect 47320 18757 47348 18788
rect 48700 18757 48728 18924
rect 50798 18912 50804 18924
rect 50856 18912 50862 18964
rect 51074 18912 51080 18964
rect 51132 18912 51138 18964
rect 48792 18788 49740 18816
rect 47029 18751 47087 18757
rect 47029 18748 47041 18751
rect 46860 18720 47041 18748
rect 45741 18683 45799 18689
rect 45741 18680 45753 18683
rect 44876 18652 45753 18680
rect 44876 18640 44882 18652
rect 45741 18649 45753 18652
rect 45787 18649 45799 18683
rect 45741 18643 45799 18649
rect 45941 18683 45999 18689
rect 45941 18649 45953 18683
rect 45987 18649 45999 18683
rect 45941 18643 45999 18649
rect 37001 18615 37059 18621
rect 37001 18581 37013 18615
rect 37047 18581 37059 18615
rect 37001 18575 37059 18581
rect 37366 18572 37372 18624
rect 37424 18612 37430 18624
rect 37829 18615 37887 18621
rect 37829 18612 37841 18615
rect 37424 18584 37841 18612
rect 37424 18572 37430 18584
rect 37829 18581 37841 18584
rect 37875 18581 37887 18615
rect 37829 18575 37887 18581
rect 38565 18615 38623 18621
rect 38565 18581 38577 18615
rect 38611 18612 38623 18615
rect 38746 18612 38752 18624
rect 38611 18584 38752 18612
rect 38611 18581 38623 18584
rect 38565 18575 38623 18581
rect 38746 18572 38752 18584
rect 38804 18572 38810 18624
rect 38930 18572 38936 18624
rect 38988 18572 38994 18624
rect 39482 18572 39488 18624
rect 39540 18572 39546 18624
rect 40681 18615 40739 18621
rect 40681 18581 40693 18615
rect 40727 18612 40739 18615
rect 41598 18612 41604 18624
rect 40727 18584 41604 18612
rect 40727 18581 40739 18584
rect 40681 18575 40739 18581
rect 41598 18572 41604 18584
rect 41656 18572 41662 18624
rect 43165 18615 43223 18621
rect 43165 18581 43177 18615
rect 43211 18612 43223 18615
rect 43441 18615 43499 18621
rect 43441 18612 43453 18615
rect 43211 18584 43453 18612
rect 43211 18581 43223 18584
rect 43165 18575 43223 18581
rect 43441 18581 43453 18584
rect 43487 18581 43499 18615
rect 43441 18575 43499 18581
rect 44729 18615 44787 18621
rect 44729 18581 44741 18615
rect 44775 18612 44787 18615
rect 45002 18612 45008 18624
rect 44775 18584 45008 18612
rect 44775 18581 44787 18584
rect 44729 18575 44787 18581
rect 45002 18572 45008 18584
rect 45060 18572 45066 18624
rect 45646 18572 45652 18624
rect 45704 18572 45710 18624
rect 46474 18572 46480 18624
rect 46532 18612 46538 18624
rect 46860 18612 46888 18720
rect 47029 18717 47041 18720
rect 47075 18717 47087 18751
rect 47029 18711 47087 18717
rect 47213 18751 47271 18757
rect 47213 18717 47225 18751
rect 47259 18717 47271 18751
rect 47213 18711 47271 18717
rect 47305 18751 47363 18757
rect 47305 18717 47317 18751
rect 47351 18717 47363 18751
rect 47305 18711 47363 18717
rect 48685 18751 48743 18757
rect 48685 18717 48697 18751
rect 48731 18717 48743 18751
rect 48685 18711 48743 18717
rect 47228 18680 47256 18711
rect 47228 18652 47624 18680
rect 46532 18584 46888 18612
rect 47596 18612 47624 18652
rect 47670 18640 47676 18692
rect 47728 18640 47734 18692
rect 48222 18640 48228 18692
rect 48280 18680 48286 18692
rect 48409 18683 48467 18689
rect 48409 18680 48421 18683
rect 48280 18652 48421 18680
rect 48280 18640 48286 18652
rect 48409 18649 48421 18652
rect 48455 18649 48467 18683
rect 48792 18680 48820 18788
rect 49712 18760 49740 18788
rect 50614 18776 50620 18828
rect 50672 18776 50678 18828
rect 50798 18776 50804 18828
rect 50856 18776 50862 18828
rect 48866 18708 48872 18760
rect 48924 18708 48930 18760
rect 48961 18751 49019 18757
rect 48961 18717 48973 18751
rect 49007 18717 49019 18751
rect 48961 18711 49019 18717
rect 48409 18643 48467 18649
rect 48700 18652 48820 18680
rect 48976 18680 49004 18711
rect 49694 18708 49700 18760
rect 49752 18748 49758 18760
rect 50525 18751 50583 18757
rect 50525 18748 50537 18751
rect 49752 18720 50537 18748
rect 49752 18708 49758 18720
rect 50525 18717 50537 18720
rect 50571 18717 50583 18751
rect 50985 18751 51043 18757
rect 50985 18748 50997 18751
rect 50525 18711 50583 18717
rect 50724 18720 50997 18748
rect 50724 18680 50752 18720
rect 50985 18717 50997 18720
rect 51031 18717 51043 18751
rect 50985 18711 51043 18717
rect 48976 18652 50752 18680
rect 48700 18612 48728 18652
rect 50724 18624 50752 18652
rect 47596 18584 48728 18612
rect 46532 18572 46538 18584
rect 48774 18572 48780 18624
rect 48832 18572 48838 18624
rect 48958 18572 48964 18624
rect 49016 18612 49022 18624
rect 49053 18615 49111 18621
rect 49053 18612 49065 18615
rect 49016 18584 49065 18612
rect 49016 18572 49022 18584
rect 49053 18581 49065 18584
rect 49099 18581 49111 18615
rect 49053 18575 49111 18581
rect 50154 18572 50160 18624
rect 50212 18572 50218 18624
rect 50706 18572 50712 18624
rect 50764 18572 50770 18624
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 26694 18368 26700 18420
rect 26752 18408 26758 18420
rect 30101 18411 30159 18417
rect 30101 18408 30113 18411
rect 26752 18380 30113 18408
rect 26752 18368 26758 18380
rect 30101 18377 30113 18380
rect 30147 18408 30159 18411
rect 31846 18408 31852 18420
rect 30147 18380 31852 18408
rect 30147 18377 30159 18380
rect 30101 18371 30159 18377
rect 31846 18368 31852 18380
rect 31904 18368 31910 18420
rect 33413 18411 33471 18417
rect 33413 18408 33425 18411
rect 32140 18380 33425 18408
rect 29181 18343 29239 18349
rect 29181 18309 29193 18343
rect 29227 18309 29239 18343
rect 29181 18303 29239 18309
rect 27246 18232 27252 18284
rect 27304 18272 27310 18284
rect 27617 18275 27675 18281
rect 27617 18272 27629 18275
rect 27304 18244 27629 18272
rect 27304 18232 27310 18244
rect 27617 18241 27629 18244
rect 27663 18241 27675 18275
rect 27617 18235 27675 18241
rect 29196 18204 29224 18303
rect 29638 18300 29644 18352
rect 29696 18300 29702 18352
rect 30006 18300 30012 18352
rect 30064 18300 30070 18352
rect 30190 18300 30196 18352
rect 30248 18300 30254 18352
rect 31297 18343 31355 18349
rect 31297 18309 31309 18343
rect 31343 18340 31355 18343
rect 31754 18340 31760 18352
rect 31343 18312 31760 18340
rect 31343 18309 31355 18312
rect 31297 18303 31355 18309
rect 31754 18300 31760 18312
rect 31812 18300 31818 18352
rect 29457 18275 29515 18281
rect 29457 18241 29469 18275
rect 29503 18272 29515 18275
rect 29546 18272 29552 18284
rect 29503 18244 29552 18272
rect 29503 18241 29515 18244
rect 29457 18235 29515 18241
rect 29546 18232 29552 18244
rect 29604 18232 29610 18284
rect 30024 18204 30052 18300
rect 29196 18176 30052 18204
rect 27798 18096 27804 18148
rect 27856 18136 27862 18148
rect 28350 18136 28356 18148
rect 27856 18108 28356 18136
rect 27856 18096 27862 18108
rect 28350 18096 28356 18108
rect 28408 18136 28414 18148
rect 28813 18139 28871 18145
rect 28813 18136 28825 18139
rect 28408 18108 28825 18136
rect 28408 18096 28414 18108
rect 28813 18105 28825 18108
rect 28859 18105 28871 18139
rect 29825 18139 29883 18145
rect 29825 18136 29837 18139
rect 28813 18099 28871 18105
rect 29196 18108 29837 18136
rect 27982 18028 27988 18080
rect 28040 18068 28046 18080
rect 29196 18077 29224 18108
rect 29825 18105 29837 18108
rect 29871 18105 29883 18139
rect 30208 18136 30236 18300
rect 30653 18275 30711 18281
rect 30653 18241 30665 18275
rect 30699 18241 30711 18275
rect 30653 18235 30711 18241
rect 31481 18275 31539 18281
rect 31481 18241 31493 18275
rect 31527 18241 31539 18275
rect 31481 18235 31539 18241
rect 30469 18139 30527 18145
rect 30469 18136 30481 18139
rect 30208 18108 30481 18136
rect 29825 18099 29883 18105
rect 30469 18105 30481 18108
rect 30515 18105 30527 18139
rect 30469 18099 30527 18105
rect 28261 18071 28319 18077
rect 28261 18068 28273 18071
rect 28040 18040 28273 18068
rect 28040 18028 28046 18040
rect 28261 18037 28273 18040
rect 28307 18037 28319 18071
rect 28261 18031 28319 18037
rect 29181 18071 29239 18077
rect 29181 18037 29193 18071
rect 29227 18037 29239 18071
rect 29181 18031 29239 18037
rect 29365 18071 29423 18077
rect 29365 18037 29377 18071
rect 29411 18068 29423 18071
rect 30668 18068 30696 18235
rect 31496 18204 31524 18235
rect 31570 18232 31576 18284
rect 31628 18272 31634 18284
rect 31628 18244 32076 18272
rect 31628 18232 31634 18244
rect 32048 18216 32076 18244
rect 32140 18216 32168 18380
rect 31496 18176 31616 18204
rect 31588 18080 31616 18176
rect 32030 18164 32036 18216
rect 32088 18164 32094 18216
rect 32122 18164 32128 18216
rect 32180 18164 32186 18216
rect 32784 18204 32812 18380
rect 33413 18377 33425 18380
rect 33459 18377 33471 18411
rect 33413 18371 33471 18377
rect 33505 18411 33563 18417
rect 33505 18377 33517 18411
rect 33551 18408 33563 18411
rect 33551 18380 33640 18408
rect 33551 18377 33563 18380
rect 33505 18371 33563 18377
rect 33612 18352 33640 18380
rect 33686 18368 33692 18420
rect 33744 18368 33750 18420
rect 33991 18411 34049 18417
rect 33991 18377 34003 18411
rect 34037 18408 34049 18411
rect 34146 18408 34152 18420
rect 34037 18380 34152 18408
rect 34037 18377 34049 18380
rect 33991 18371 34049 18377
rect 34146 18368 34152 18380
rect 34204 18368 34210 18420
rect 38194 18408 38200 18420
rect 36740 18380 38200 18408
rect 32950 18300 32956 18352
rect 33008 18340 33014 18352
rect 33137 18343 33195 18349
rect 33137 18340 33149 18343
rect 33008 18312 33149 18340
rect 33008 18300 33014 18312
rect 33137 18309 33149 18312
rect 33183 18309 33195 18343
rect 33137 18303 33195 18309
rect 33594 18300 33600 18352
rect 33652 18340 33658 18352
rect 33781 18343 33839 18349
rect 33781 18340 33793 18343
rect 33652 18312 33793 18340
rect 33652 18300 33658 18312
rect 33781 18309 33793 18312
rect 33827 18309 33839 18343
rect 33781 18303 33839 18309
rect 32861 18275 32919 18281
rect 32861 18241 32873 18275
rect 32907 18272 32919 18275
rect 32907 18244 33180 18272
rect 32907 18241 32919 18244
rect 32861 18235 32919 18241
rect 32784 18176 33088 18204
rect 32214 18096 32220 18148
rect 32272 18136 32278 18148
rect 32953 18139 33011 18145
rect 32953 18136 32965 18139
rect 32272 18108 32965 18136
rect 32272 18096 32278 18108
rect 32953 18105 32965 18108
rect 32999 18105 33011 18139
rect 32953 18099 33011 18105
rect 29411 18040 30696 18068
rect 29411 18037 29423 18040
rect 29365 18031 29423 18037
rect 31294 18028 31300 18080
rect 31352 18028 31358 18080
rect 31570 18028 31576 18080
rect 31628 18068 31634 18080
rect 32398 18068 32404 18080
rect 31628 18040 32404 18068
rect 31628 18028 31634 18040
rect 32398 18028 32404 18040
rect 32456 18068 32462 18080
rect 32769 18071 32827 18077
rect 32769 18068 32781 18071
rect 32456 18040 32781 18068
rect 32456 18028 32462 18040
rect 32769 18037 32781 18040
rect 32815 18037 32827 18071
rect 32769 18031 32827 18037
rect 32858 18028 32864 18080
rect 32916 18028 32922 18080
rect 33060 18068 33088 18176
rect 33152 18136 33180 18244
rect 33318 18232 33324 18284
rect 33376 18232 33382 18284
rect 35253 18275 35311 18281
rect 35253 18241 35265 18275
rect 35299 18272 35311 18275
rect 35342 18272 35348 18284
rect 35299 18244 35348 18272
rect 35299 18241 35311 18244
rect 35253 18235 35311 18241
rect 35342 18232 35348 18244
rect 35400 18232 35406 18284
rect 35520 18275 35578 18281
rect 35520 18241 35532 18275
rect 35566 18272 35578 18275
rect 35802 18272 35808 18284
rect 35566 18244 35808 18272
rect 35566 18241 35578 18244
rect 35520 18235 35578 18241
rect 35802 18232 35808 18244
rect 35860 18232 35866 18284
rect 36740 18276 36768 18380
rect 38194 18368 38200 18380
rect 38252 18368 38258 18420
rect 38286 18368 38292 18420
rect 38344 18408 38350 18420
rect 38381 18411 38439 18417
rect 38381 18408 38393 18411
rect 38344 18380 38393 18408
rect 38344 18368 38350 18380
rect 38381 18377 38393 18380
rect 38427 18377 38439 18411
rect 38930 18408 38936 18420
rect 38381 18371 38439 18377
rect 38672 18380 38936 18408
rect 36998 18300 37004 18352
rect 37056 18300 37062 18352
rect 37369 18343 37427 18349
rect 37369 18309 37381 18343
rect 37415 18309 37427 18343
rect 37369 18303 37427 18309
rect 37585 18343 37643 18349
rect 37585 18309 37597 18343
rect 37631 18340 37643 18343
rect 37631 18312 38424 18340
rect 37631 18309 37643 18312
rect 37585 18303 37643 18309
rect 36817 18276 36875 18281
rect 36740 18275 36875 18276
rect 36740 18248 36829 18275
rect 36817 18241 36829 18248
rect 36863 18241 36875 18275
rect 37016 18272 37044 18300
rect 36817 18235 36875 18241
rect 36930 18244 37044 18272
rect 37384 18272 37412 18303
rect 38396 18284 38424 18312
rect 37826 18272 37832 18284
rect 37384 18244 37832 18272
rect 33689 18207 33747 18213
rect 33689 18173 33701 18207
rect 33735 18204 33747 18207
rect 34698 18204 34704 18216
rect 33735 18176 34704 18204
rect 33735 18173 33747 18176
rect 33689 18167 33747 18173
rect 34698 18164 34704 18176
rect 34756 18164 34762 18216
rect 36930 18213 36958 18244
rect 37826 18232 37832 18244
rect 37884 18232 37890 18284
rect 38105 18275 38163 18281
rect 38105 18241 38117 18275
rect 38151 18241 38163 18275
rect 38105 18235 38163 18241
rect 36909 18207 36967 18213
rect 36909 18173 36921 18207
rect 36955 18173 36967 18207
rect 36909 18167 36967 18173
rect 37090 18164 37096 18216
rect 37148 18204 37154 18216
rect 37274 18204 37280 18216
rect 37148 18176 37280 18204
rect 37148 18164 37154 18176
rect 37274 18164 37280 18176
rect 37332 18164 37338 18216
rect 34146 18136 34152 18148
rect 33152 18108 34152 18136
rect 34146 18096 34152 18108
rect 34204 18096 34210 18148
rect 36633 18139 36691 18145
rect 36633 18105 36645 18139
rect 36679 18136 36691 18139
rect 37182 18136 37188 18148
rect 36679 18108 37188 18136
rect 36679 18105 36691 18108
rect 36633 18099 36691 18105
rect 37182 18096 37188 18108
rect 37240 18136 37246 18148
rect 38120 18136 38148 18235
rect 38378 18232 38384 18284
rect 38436 18232 38442 18284
rect 38672 18281 38700 18380
rect 38930 18368 38936 18380
rect 38988 18408 38994 18420
rect 40221 18411 40279 18417
rect 40221 18408 40233 18411
rect 38988 18380 40233 18408
rect 38988 18368 38994 18380
rect 40221 18377 40233 18380
rect 40267 18377 40279 18411
rect 40221 18371 40279 18377
rect 41046 18368 41052 18420
rect 41104 18408 41110 18420
rect 41141 18411 41199 18417
rect 41141 18408 41153 18411
rect 41104 18380 41153 18408
rect 41104 18368 41110 18380
rect 41141 18377 41153 18380
rect 41187 18377 41199 18411
rect 41141 18371 41199 18377
rect 42610 18368 42616 18420
rect 42668 18368 42674 18420
rect 44358 18368 44364 18420
rect 44416 18408 44422 18420
rect 44913 18411 44971 18417
rect 44913 18408 44925 18411
rect 44416 18380 44925 18408
rect 44416 18368 44422 18380
rect 44913 18377 44925 18380
rect 44959 18377 44971 18411
rect 44913 18371 44971 18377
rect 45005 18411 45063 18417
rect 45005 18377 45017 18411
rect 45051 18408 45063 18411
rect 45051 18380 45600 18408
rect 45051 18377 45063 18380
rect 45005 18371 45063 18377
rect 39942 18340 39948 18352
rect 38856 18312 39948 18340
rect 38856 18281 38884 18312
rect 39942 18300 39948 18312
rect 40000 18340 40006 18352
rect 42061 18343 42119 18349
rect 42061 18340 42073 18343
rect 40000 18312 42073 18340
rect 40000 18300 40006 18312
rect 42061 18309 42073 18312
rect 42107 18340 42119 18343
rect 42107 18312 42472 18340
rect 42107 18309 42119 18312
rect 42061 18303 42119 18309
rect 38657 18275 38715 18281
rect 38657 18241 38669 18275
rect 38703 18241 38715 18275
rect 38657 18235 38715 18241
rect 38841 18275 38899 18281
rect 38841 18241 38853 18275
rect 38887 18241 38899 18275
rect 38841 18235 38899 18241
rect 38930 18232 38936 18284
rect 38988 18272 38994 18284
rect 39097 18275 39155 18281
rect 39097 18272 39109 18275
rect 38988 18244 39109 18272
rect 38988 18232 38994 18244
rect 39097 18241 39109 18244
rect 39143 18241 39155 18275
rect 39097 18235 39155 18241
rect 41049 18275 41107 18281
rect 41049 18241 41061 18275
rect 41095 18272 41107 18275
rect 41138 18272 41144 18284
rect 41095 18244 41144 18272
rect 41095 18241 41107 18244
rect 41049 18235 41107 18241
rect 41138 18232 41144 18244
rect 41196 18232 41202 18284
rect 41230 18232 41236 18284
rect 41288 18232 41294 18284
rect 41322 18232 41328 18284
rect 41380 18232 41386 18284
rect 42444 18281 42472 18312
rect 42429 18275 42487 18281
rect 42429 18241 42441 18275
rect 42475 18241 42487 18275
rect 42628 18272 42656 18368
rect 42685 18275 42743 18281
rect 42685 18272 42697 18275
rect 42628 18244 42697 18272
rect 42429 18235 42487 18241
rect 42685 18241 42697 18244
rect 42731 18241 42743 18275
rect 42685 18235 42743 18241
rect 44358 18232 44364 18284
rect 44416 18272 44422 18284
rect 44818 18272 44824 18284
rect 44416 18244 44824 18272
rect 44416 18232 44422 18244
rect 44818 18232 44824 18244
rect 44876 18232 44882 18284
rect 45278 18232 45284 18284
rect 45336 18232 45342 18284
rect 45373 18275 45431 18281
rect 45373 18241 45385 18275
rect 45419 18241 45431 18275
rect 45373 18235 45431 18241
rect 41340 18204 41368 18232
rect 40144 18176 41368 18204
rect 37240 18108 38148 18136
rect 37240 18096 37246 18108
rect 33965 18071 34023 18077
rect 33965 18068 33977 18071
rect 33060 18040 33977 18068
rect 33965 18037 33977 18040
rect 34011 18037 34023 18071
rect 33965 18031 34023 18037
rect 36354 18028 36360 18080
rect 36412 18068 36418 18080
rect 36906 18068 36912 18080
rect 36412 18040 36912 18068
rect 36412 18028 36418 18040
rect 36906 18028 36912 18040
rect 36964 18028 36970 18080
rect 37001 18071 37059 18077
rect 37001 18037 37013 18071
rect 37047 18068 37059 18071
rect 37274 18068 37280 18080
rect 37047 18040 37280 18068
rect 37047 18037 37059 18040
rect 37001 18031 37059 18037
rect 37274 18028 37280 18040
rect 37332 18028 37338 18080
rect 37568 18077 37596 18108
rect 38194 18096 38200 18148
rect 38252 18136 38258 18148
rect 38838 18136 38844 18148
rect 38252 18108 38844 18136
rect 38252 18096 38258 18108
rect 38838 18096 38844 18108
rect 38896 18096 38902 18148
rect 37553 18071 37611 18077
rect 37553 18037 37565 18071
rect 37599 18037 37611 18071
rect 37553 18031 37611 18037
rect 37737 18071 37795 18077
rect 37737 18037 37749 18071
rect 37783 18068 37795 18071
rect 38212 18068 38240 18096
rect 37783 18040 38240 18068
rect 37783 18037 37795 18040
rect 37737 18031 37795 18037
rect 38562 18028 38568 18080
rect 38620 18068 38626 18080
rect 40144 18068 40172 18176
rect 43809 18139 43867 18145
rect 43809 18105 43821 18139
rect 43855 18136 43867 18139
rect 43898 18136 43904 18148
rect 43855 18108 43904 18136
rect 43855 18105 43867 18108
rect 43809 18099 43867 18105
rect 43898 18096 43904 18108
rect 43956 18136 43962 18148
rect 45388 18136 45416 18235
rect 45462 18232 45468 18284
rect 45520 18232 45526 18284
rect 43956 18108 45416 18136
rect 45480 18136 45508 18232
rect 45572 18204 45600 18380
rect 45646 18368 45652 18420
rect 45704 18368 45710 18420
rect 46566 18368 46572 18420
rect 46624 18368 46630 18420
rect 47394 18408 47400 18420
rect 47228 18380 47400 18408
rect 45664 18281 45692 18368
rect 46842 18300 46848 18352
rect 46900 18340 46906 18352
rect 47228 18349 47256 18380
rect 47394 18368 47400 18380
rect 47452 18368 47458 18420
rect 47578 18368 47584 18420
rect 47636 18408 47642 18420
rect 50062 18408 50068 18420
rect 47636 18380 50068 18408
rect 47636 18368 47642 18380
rect 47122 18343 47180 18349
rect 47122 18340 47134 18343
rect 46900 18312 47134 18340
rect 46900 18300 46906 18312
rect 47122 18309 47134 18312
rect 47168 18309 47180 18343
rect 47228 18343 47297 18349
rect 47228 18312 47251 18343
rect 47122 18303 47180 18309
rect 47239 18309 47251 18312
rect 47285 18309 47297 18343
rect 47762 18340 47768 18352
rect 47239 18303 47297 18309
rect 47412 18312 47768 18340
rect 45649 18275 45707 18281
rect 45649 18241 45661 18275
rect 45695 18241 45707 18275
rect 46474 18272 46480 18284
rect 45649 18235 45707 18241
rect 45848 18244 46480 18272
rect 45741 18207 45799 18213
rect 45741 18204 45753 18207
rect 45572 18176 45753 18204
rect 45741 18173 45753 18176
rect 45787 18173 45799 18207
rect 45741 18167 45799 18173
rect 45646 18136 45652 18148
rect 45480 18108 45652 18136
rect 43956 18096 43962 18108
rect 45646 18096 45652 18108
rect 45704 18096 45710 18148
rect 38620 18040 40172 18068
rect 38620 18028 38626 18040
rect 44082 18028 44088 18080
rect 44140 18068 44146 18080
rect 45848 18068 45876 18244
rect 46474 18232 46480 18244
rect 46532 18232 46538 18284
rect 46658 18232 46664 18284
rect 46716 18232 46722 18284
rect 46750 18232 46756 18284
rect 46808 18272 46814 18284
rect 46937 18275 46995 18281
rect 46937 18272 46949 18275
rect 46808 18244 46949 18272
rect 46808 18232 46814 18244
rect 46937 18241 46949 18244
rect 46983 18241 46995 18275
rect 46937 18235 46995 18241
rect 47029 18275 47087 18281
rect 47029 18241 47041 18275
rect 47075 18272 47087 18275
rect 47075 18244 47164 18272
rect 47075 18241 47087 18244
rect 47029 18235 47087 18241
rect 47136 18216 47164 18244
rect 47118 18164 47124 18216
rect 47176 18164 47182 18216
rect 47412 18213 47440 18312
rect 47762 18300 47768 18312
rect 47820 18300 47826 18352
rect 47578 18232 47584 18284
rect 47636 18232 47642 18284
rect 48958 18232 48964 18284
rect 49016 18232 49022 18284
rect 49712 18281 49740 18380
rect 50062 18368 50068 18380
rect 50120 18368 50126 18420
rect 50798 18368 50804 18420
rect 50856 18408 50862 18420
rect 50856 18380 51764 18408
rect 50856 18368 50862 18380
rect 51736 18349 51764 18380
rect 51721 18343 51779 18349
rect 51721 18309 51733 18343
rect 51767 18309 51779 18343
rect 51721 18303 51779 18309
rect 49697 18275 49755 18281
rect 49697 18241 49709 18275
rect 49743 18241 49755 18275
rect 49697 18235 49755 18241
rect 51074 18232 51080 18284
rect 51132 18232 51138 18284
rect 47397 18207 47455 18213
rect 47397 18173 47409 18207
rect 47443 18173 47455 18207
rect 47857 18207 47915 18213
rect 47857 18204 47869 18207
rect 47397 18167 47455 18173
rect 47504 18176 47869 18204
rect 47504 18136 47532 18176
rect 47857 18173 47869 18176
rect 47903 18173 47915 18207
rect 47857 18167 47915 18173
rect 47946 18164 47952 18216
rect 48004 18204 48010 18216
rect 48866 18204 48872 18216
rect 48004 18176 48872 18204
rect 48004 18164 48010 18176
rect 48866 18164 48872 18176
rect 48924 18204 48930 18216
rect 49605 18207 49663 18213
rect 49605 18204 49617 18207
rect 48924 18176 49617 18204
rect 48924 18164 48930 18176
rect 49605 18173 49617 18176
rect 49651 18173 49663 18207
rect 49605 18167 49663 18173
rect 49970 18164 49976 18216
rect 50028 18164 50034 18216
rect 46768 18108 47532 18136
rect 44140 18040 45876 18068
rect 44140 18028 44146 18040
rect 46382 18028 46388 18080
rect 46440 18028 46446 18080
rect 46768 18077 46796 18108
rect 46753 18071 46811 18077
rect 46753 18037 46765 18071
rect 46799 18037 46811 18071
rect 46753 18031 46811 18037
rect 46934 18028 46940 18080
rect 46992 18068 46998 18080
rect 47670 18068 47676 18080
rect 46992 18040 47676 18068
rect 46992 18028 46998 18040
rect 47670 18028 47676 18040
rect 47728 18028 47734 18080
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 1820 17836 27200 17864
rect 1820 17824 1826 17836
rect 27172 17796 27200 17836
rect 27246 17824 27252 17876
rect 27304 17864 27310 17876
rect 27433 17867 27491 17873
rect 27433 17864 27445 17867
rect 27304 17836 27445 17864
rect 27304 17824 27310 17836
rect 27433 17833 27445 17836
rect 27479 17833 27491 17867
rect 27433 17827 27491 17833
rect 28000 17836 29684 17864
rect 28000 17796 28028 17836
rect 27172 17768 28028 17796
rect 28077 17799 28135 17805
rect 28077 17765 28089 17799
rect 28123 17765 28135 17799
rect 28077 17759 28135 17765
rect 27798 17688 27804 17740
rect 27856 17688 27862 17740
rect 25222 17620 25228 17672
rect 25280 17660 25286 17672
rect 26053 17663 26111 17669
rect 26053 17660 26065 17663
rect 25280 17632 26065 17660
rect 25280 17620 25286 17632
rect 26053 17629 26065 17632
rect 26099 17629 26111 17663
rect 26053 17623 26111 17629
rect 27709 17663 27767 17669
rect 27709 17629 27721 17663
rect 27755 17660 27767 17663
rect 27982 17660 27988 17672
rect 27755 17632 27988 17660
rect 27755 17629 27767 17632
rect 27709 17623 27767 17629
rect 27982 17620 27988 17632
rect 28040 17620 28046 17672
rect 28092 17660 28120 17759
rect 28169 17663 28227 17669
rect 28169 17660 28181 17663
rect 28092 17632 28181 17660
rect 28169 17629 28181 17632
rect 28215 17629 28227 17663
rect 28169 17623 28227 17629
rect 28350 17620 28356 17672
rect 28408 17620 28414 17672
rect 29656 17660 29684 17836
rect 29730 17824 29736 17876
rect 29788 17864 29794 17876
rect 30561 17867 30619 17873
rect 30561 17864 30573 17867
rect 29788 17836 30573 17864
rect 29788 17824 29794 17836
rect 30561 17833 30573 17836
rect 30607 17864 30619 17867
rect 31386 17864 31392 17876
rect 30607 17836 31392 17864
rect 30607 17833 30619 17836
rect 30561 17827 30619 17833
rect 31386 17824 31392 17836
rect 31444 17824 31450 17876
rect 32122 17824 32128 17876
rect 32180 17824 32186 17876
rect 32214 17824 32220 17876
rect 32272 17824 32278 17876
rect 34054 17824 34060 17876
rect 34112 17824 34118 17876
rect 34146 17824 34152 17876
rect 34204 17864 34210 17876
rect 34425 17867 34483 17873
rect 34425 17864 34437 17867
rect 34204 17836 34437 17864
rect 34204 17824 34210 17836
rect 34425 17833 34437 17836
rect 34471 17833 34483 17867
rect 34425 17827 34483 17833
rect 35802 17824 35808 17876
rect 35860 17824 35866 17876
rect 36446 17824 36452 17876
rect 36504 17824 36510 17876
rect 37366 17864 37372 17876
rect 36648 17836 37372 17864
rect 32030 17756 32036 17808
rect 32088 17796 32094 17808
rect 34072 17796 34100 17824
rect 32088 17768 34100 17796
rect 32088 17756 32094 17768
rect 30285 17663 30343 17669
rect 30285 17660 30297 17663
rect 29656 17632 30297 17660
rect 30285 17629 30297 17632
rect 30331 17629 30343 17663
rect 30285 17623 30343 17629
rect 26320 17595 26378 17601
rect 26320 17561 26332 17595
rect 26366 17592 26378 17595
rect 28261 17595 28319 17601
rect 28261 17592 28273 17595
rect 26366 17564 28273 17592
rect 26366 17561 26378 17564
rect 26320 17555 26378 17561
rect 28261 17561 28273 17564
rect 28307 17561 28319 17595
rect 28261 17555 28319 17561
rect 28997 17595 29055 17601
rect 28997 17561 29009 17595
rect 29043 17592 29055 17595
rect 29270 17592 29276 17604
rect 29043 17564 29276 17592
rect 29043 17561 29055 17564
rect 28997 17555 29055 17561
rect 29270 17552 29276 17564
rect 29328 17592 29334 17604
rect 29730 17592 29736 17604
rect 29328 17564 29736 17592
rect 29328 17552 29334 17564
rect 29730 17552 29736 17564
rect 29788 17552 29794 17604
rect 30101 17595 30159 17601
rect 30101 17561 30113 17595
rect 30147 17592 30159 17595
rect 30190 17592 30196 17604
rect 30147 17564 30196 17592
rect 30147 17561 30159 17564
rect 30101 17555 30159 17561
rect 30190 17552 30196 17564
rect 30248 17552 30254 17604
rect 29089 17527 29147 17533
rect 29089 17493 29101 17527
rect 29135 17524 29147 17527
rect 29362 17524 29368 17536
rect 29135 17496 29368 17524
rect 29135 17493 29147 17496
rect 29089 17487 29147 17493
rect 29362 17484 29368 17496
rect 29420 17524 29426 17536
rect 30006 17524 30012 17536
rect 29420 17496 30012 17524
rect 29420 17484 29426 17496
rect 30006 17484 30012 17496
rect 30064 17484 30070 17536
rect 30300 17524 30328 17623
rect 30742 17620 30748 17672
rect 30800 17620 30806 17672
rect 31012 17663 31070 17669
rect 31012 17629 31024 17663
rect 31058 17660 31070 17663
rect 31294 17660 31300 17672
rect 31058 17632 31300 17660
rect 31058 17629 31070 17632
rect 31012 17623 31070 17629
rect 31294 17620 31300 17632
rect 31352 17620 31358 17672
rect 32398 17620 32404 17672
rect 32456 17620 32462 17672
rect 32493 17663 32551 17669
rect 32493 17629 32505 17663
rect 32539 17660 32551 17663
rect 32591 17660 32619 17768
rect 32677 17731 32735 17737
rect 32677 17697 32689 17731
rect 32723 17728 32735 17731
rect 32858 17728 32864 17740
rect 32723 17700 32864 17728
rect 32723 17697 32735 17700
rect 32677 17691 32735 17697
rect 32858 17688 32864 17700
rect 32916 17688 32922 17740
rect 34517 17731 34575 17737
rect 34517 17697 34529 17731
rect 34563 17728 34575 17731
rect 35345 17731 35403 17737
rect 35345 17728 35357 17731
rect 34563 17700 35357 17728
rect 34563 17697 34575 17700
rect 34517 17691 34575 17697
rect 35345 17697 35357 17700
rect 35391 17697 35403 17731
rect 36464 17728 36492 17824
rect 35345 17691 35403 17697
rect 36280 17700 36492 17728
rect 32539 17632 32619 17660
rect 33413 17663 33471 17669
rect 32539 17629 32551 17632
rect 32493 17623 32551 17629
rect 33413 17629 33425 17663
rect 33459 17660 33471 17663
rect 33594 17660 33600 17672
rect 33459 17632 33600 17660
rect 33459 17629 33471 17632
rect 33413 17623 33471 17629
rect 33594 17620 33600 17632
rect 33652 17620 33658 17672
rect 33962 17620 33968 17672
rect 34020 17660 34026 17672
rect 34057 17663 34115 17669
rect 34057 17660 34069 17663
rect 34020 17632 34069 17660
rect 34020 17620 34026 17632
rect 34057 17629 34069 17632
rect 34103 17629 34115 17663
rect 34057 17623 34115 17629
rect 34241 17663 34299 17669
rect 34241 17629 34253 17663
rect 34287 17660 34299 17663
rect 34422 17660 34428 17672
rect 34287 17632 34428 17660
rect 34287 17629 34299 17632
rect 34241 17623 34299 17629
rect 34422 17620 34428 17632
rect 34480 17620 34486 17672
rect 34698 17620 34704 17672
rect 34756 17620 34762 17672
rect 36280 17669 36308 17700
rect 35989 17663 36047 17669
rect 35989 17629 36001 17663
rect 36035 17629 36047 17663
rect 35989 17623 36047 17629
rect 36265 17663 36323 17669
rect 36265 17629 36277 17663
rect 36311 17629 36323 17663
rect 36265 17623 36323 17629
rect 36449 17663 36507 17669
rect 36449 17629 36461 17663
rect 36495 17660 36507 17663
rect 36648 17660 36676 17836
rect 37366 17824 37372 17836
rect 37424 17824 37430 17876
rect 37826 17824 37832 17876
rect 37884 17864 37890 17876
rect 38565 17867 38623 17873
rect 38565 17864 38577 17867
rect 37884 17836 38577 17864
rect 37884 17824 37890 17836
rect 38565 17833 38577 17836
rect 38611 17833 38623 17867
rect 38565 17827 38623 17833
rect 37182 17756 37188 17808
rect 37240 17756 37246 17808
rect 37200 17728 37228 17756
rect 36832 17700 37228 17728
rect 38580 17728 38608 17827
rect 38654 17824 38660 17876
rect 38712 17864 38718 17876
rect 39301 17867 39359 17873
rect 39301 17864 39313 17867
rect 38712 17836 39313 17864
rect 38712 17824 38718 17836
rect 39301 17833 39313 17836
rect 39347 17833 39359 17867
rect 39301 17827 39359 17833
rect 43349 17867 43407 17873
rect 43349 17833 43361 17867
rect 43395 17864 43407 17867
rect 43438 17864 43444 17876
rect 43395 17836 43444 17864
rect 43395 17833 43407 17836
rect 43349 17827 43407 17833
rect 43438 17824 43444 17836
rect 43496 17824 43502 17876
rect 44082 17824 44088 17876
rect 44140 17864 44146 17876
rect 44140 17836 44312 17864
rect 44140 17824 44146 17836
rect 43714 17756 43720 17808
rect 43772 17796 43778 17808
rect 44284 17805 44312 17836
rect 45278 17824 45284 17876
rect 45336 17864 45342 17876
rect 46474 17864 46480 17876
rect 45336 17836 46480 17864
rect 45336 17824 45342 17836
rect 46474 17824 46480 17836
rect 46532 17824 46538 17876
rect 46842 17824 46848 17876
rect 46900 17864 46906 17876
rect 47305 17867 47363 17873
rect 47305 17864 47317 17867
rect 46900 17836 47317 17864
rect 46900 17824 46906 17836
rect 47305 17833 47317 17836
rect 47351 17833 47363 17867
rect 47305 17827 47363 17833
rect 49237 17867 49295 17873
rect 49237 17833 49249 17867
rect 49283 17864 49295 17867
rect 49970 17864 49976 17876
rect 49283 17836 49976 17864
rect 49283 17833 49295 17836
rect 49237 17827 49295 17833
rect 49970 17824 49976 17836
rect 50028 17824 50034 17876
rect 50617 17867 50675 17873
rect 50617 17833 50629 17867
rect 50663 17864 50675 17867
rect 51074 17864 51080 17876
rect 50663 17836 51080 17864
rect 50663 17833 50675 17836
rect 50617 17827 50675 17833
rect 51074 17824 51080 17836
rect 51132 17824 51138 17876
rect 44177 17799 44235 17805
rect 44177 17796 44189 17799
rect 43772 17768 44189 17796
rect 43772 17756 43778 17768
rect 44177 17765 44189 17768
rect 44223 17765 44235 17799
rect 44177 17759 44235 17765
rect 44269 17799 44327 17805
rect 44269 17765 44281 17799
rect 44315 17765 44327 17799
rect 44269 17759 44327 17765
rect 38657 17731 38715 17737
rect 38657 17728 38669 17731
rect 38580 17700 38669 17728
rect 36832 17669 36860 17700
rect 38657 17697 38669 17700
rect 38703 17697 38715 17731
rect 38657 17691 38715 17697
rect 39112 17700 39620 17728
rect 36495 17632 36676 17660
rect 36725 17663 36783 17669
rect 36495 17629 36507 17632
rect 36449 17623 36507 17629
rect 36725 17629 36737 17663
rect 36771 17629 36783 17663
rect 36725 17623 36783 17629
rect 36817 17663 36875 17669
rect 36817 17629 36829 17663
rect 36863 17629 36875 17663
rect 36817 17623 36875 17629
rect 32217 17595 32275 17601
rect 32217 17561 32229 17595
rect 32263 17592 32275 17595
rect 36004 17592 36032 17623
rect 36541 17595 36599 17601
rect 36541 17592 36553 17595
rect 32263 17564 34008 17592
rect 36004 17564 36553 17592
rect 32263 17561 32275 17564
rect 32217 17555 32275 17561
rect 33134 17524 33140 17536
rect 30300 17496 33140 17524
rect 33134 17484 33140 17496
rect 33192 17484 33198 17536
rect 33226 17484 33232 17536
rect 33284 17484 33290 17536
rect 33980 17533 34008 17564
rect 36541 17561 36553 17564
rect 36587 17561 36599 17595
rect 36541 17555 36599 17561
rect 36630 17552 36636 17604
rect 36688 17592 36694 17604
rect 36740 17592 36768 17623
rect 36906 17620 36912 17672
rect 36964 17660 36970 17672
rect 37001 17663 37059 17669
rect 37001 17660 37013 17663
rect 36964 17632 37013 17660
rect 36964 17620 36970 17632
rect 37001 17629 37013 17632
rect 37047 17629 37059 17663
rect 37001 17623 37059 17629
rect 37093 17663 37151 17669
rect 37093 17629 37105 17663
rect 37139 17629 37151 17663
rect 37093 17623 37151 17629
rect 36688 17564 36768 17592
rect 37108 17592 37136 17623
rect 37182 17620 37188 17672
rect 37240 17620 37246 17672
rect 37274 17620 37280 17672
rect 37332 17660 37338 17672
rect 37441 17663 37499 17669
rect 37441 17660 37453 17663
rect 37332 17632 37453 17660
rect 37332 17620 37338 17632
rect 37441 17629 37453 17632
rect 37487 17629 37499 17663
rect 37441 17623 37499 17629
rect 37918 17620 37924 17672
rect 37976 17620 37982 17672
rect 37936 17592 37964 17620
rect 37108 17564 37964 17592
rect 36688 17552 36694 17564
rect 33965 17527 34023 17533
rect 33965 17493 33977 17527
rect 34011 17493 34023 17527
rect 33965 17487 34023 17493
rect 36170 17484 36176 17536
rect 36228 17524 36234 17536
rect 39112 17524 39140 17700
rect 39592 17669 39620 17700
rect 43548 17700 43944 17728
rect 43548 17669 43576 17700
rect 43916 17672 43944 17700
rect 46584 17700 46796 17728
rect 39393 17663 39451 17669
rect 39393 17629 39405 17663
rect 39439 17629 39451 17663
rect 39393 17623 39451 17629
rect 39577 17663 39635 17669
rect 39577 17629 39589 17663
rect 39623 17629 39635 17663
rect 39577 17623 39635 17629
rect 43533 17663 43591 17669
rect 43533 17629 43545 17663
rect 43579 17629 43591 17663
rect 43533 17623 43591 17629
rect 39408 17592 39436 17623
rect 43806 17620 43812 17672
rect 43864 17620 43870 17672
rect 43898 17620 43904 17672
rect 43956 17660 43962 17672
rect 44085 17663 44143 17669
rect 44085 17660 44097 17663
rect 43956 17632 44097 17660
rect 43956 17620 43962 17632
rect 44085 17629 44097 17632
rect 44131 17629 44143 17663
rect 44085 17623 44143 17629
rect 44358 17620 44364 17672
rect 44416 17620 44422 17672
rect 44450 17620 44456 17672
rect 44508 17660 44514 17672
rect 45097 17663 45155 17669
rect 45097 17660 45109 17663
rect 44508 17632 45109 17660
rect 44508 17620 44514 17632
rect 45097 17629 45109 17632
rect 45143 17660 45155 17663
rect 46584 17660 46612 17700
rect 46768 17672 46796 17700
rect 47578 17688 47584 17740
rect 47636 17728 47642 17740
rect 48133 17731 48191 17737
rect 48133 17728 48145 17731
rect 47636 17700 48145 17728
rect 47636 17688 47642 17700
rect 48133 17697 48145 17700
rect 48179 17697 48191 17731
rect 48133 17691 48191 17697
rect 49053 17731 49111 17737
rect 49053 17697 49065 17731
rect 49099 17728 49111 17731
rect 49234 17728 49240 17740
rect 49099 17700 49240 17728
rect 49099 17697 49111 17700
rect 49053 17691 49111 17697
rect 49234 17688 49240 17700
rect 49292 17688 49298 17740
rect 45143 17632 46612 17660
rect 45143 17629 45155 17632
rect 45097 17623 45155 17629
rect 46658 17620 46664 17672
rect 46716 17620 46722 17672
rect 46750 17620 46756 17672
rect 46808 17620 46814 17672
rect 46934 17620 46940 17672
rect 46992 17660 46998 17672
rect 47397 17663 47455 17669
rect 47397 17660 47409 17663
rect 46992 17632 47409 17660
rect 46992 17620 46998 17632
rect 47397 17629 47409 17632
rect 47443 17629 47455 17663
rect 47397 17623 47455 17629
rect 49421 17663 49479 17669
rect 49421 17629 49433 17663
rect 49467 17660 49479 17663
rect 50154 17660 50160 17672
rect 49467 17632 50160 17660
rect 49467 17629 49479 17632
rect 49421 17623 49479 17629
rect 50154 17620 50160 17632
rect 50212 17620 50218 17672
rect 50525 17663 50583 17669
rect 50525 17629 50537 17663
rect 50571 17660 50583 17663
rect 50706 17660 50712 17672
rect 50571 17632 50712 17660
rect 50571 17629 50583 17632
rect 50525 17623 50583 17629
rect 41598 17592 41604 17604
rect 39408 17564 41604 17592
rect 41598 17552 41604 17564
rect 41656 17552 41662 17604
rect 43717 17595 43775 17601
rect 43717 17561 43729 17595
rect 43763 17592 43775 17595
rect 44376 17592 44404 17620
rect 43763 17564 44404 17592
rect 45364 17595 45422 17601
rect 43763 17561 43775 17564
rect 43717 17555 43775 17561
rect 45364 17561 45376 17595
rect 45410 17592 45422 17595
rect 46382 17592 46388 17604
rect 45410 17564 46388 17592
rect 45410 17561 45422 17564
rect 45364 17555 45422 17561
rect 46382 17552 46388 17564
rect 46440 17552 46446 17604
rect 50540 17592 50568 17623
rect 50706 17620 50712 17632
rect 50764 17620 50770 17672
rect 50080 17564 50568 17592
rect 50080 17536 50108 17564
rect 36228 17496 39140 17524
rect 39485 17527 39543 17533
rect 36228 17484 36234 17496
rect 39485 17493 39497 17527
rect 39531 17524 39543 17527
rect 39574 17524 39580 17536
rect 39531 17496 39580 17524
rect 39531 17493 39543 17496
rect 39485 17487 39543 17493
rect 39574 17484 39580 17496
rect 39632 17484 39638 17536
rect 43162 17484 43168 17536
rect 43220 17524 43226 17536
rect 43901 17527 43959 17533
rect 43901 17524 43913 17527
rect 43220 17496 43913 17524
rect 43220 17484 43226 17496
rect 43901 17493 43913 17496
rect 43947 17493 43959 17527
rect 43901 17487 43959 17493
rect 48406 17484 48412 17536
rect 48464 17484 48470 17536
rect 48774 17484 48780 17536
rect 48832 17484 48838 17536
rect 48866 17484 48872 17536
rect 48924 17484 48930 17536
rect 50062 17484 50068 17536
rect 50120 17484 50126 17536
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 29365 17323 29423 17329
rect 29365 17289 29377 17323
rect 29411 17289 29423 17323
rect 29365 17283 29423 17289
rect 29178 17252 29184 17264
rect 27908 17224 29184 17252
rect 26145 17187 26203 17193
rect 26145 17153 26157 17187
rect 26191 17184 26203 17187
rect 26602 17184 26608 17196
rect 26191 17156 26608 17184
rect 26191 17153 26203 17156
rect 26145 17147 26203 17153
rect 26602 17144 26608 17156
rect 26660 17144 26666 17196
rect 27522 17076 27528 17128
rect 27580 17116 27586 17128
rect 27908 17125 27936 17224
rect 29178 17212 29184 17224
rect 29236 17212 29242 17264
rect 28160 17187 28218 17193
rect 28160 17153 28172 17187
rect 28206 17184 28218 17187
rect 29380 17184 29408 17283
rect 31754 17280 31760 17332
rect 31812 17320 31818 17332
rect 31849 17323 31907 17329
rect 31849 17320 31861 17323
rect 31812 17292 31861 17320
rect 31812 17280 31818 17292
rect 31849 17289 31861 17292
rect 31895 17289 31907 17323
rect 31849 17283 31907 17289
rect 33594 17280 33600 17332
rect 33652 17280 33658 17332
rect 34698 17280 34704 17332
rect 34756 17320 34762 17332
rect 35069 17323 35127 17329
rect 35069 17320 35081 17323
rect 34756 17292 35081 17320
rect 34756 17280 34762 17292
rect 35069 17289 35081 17292
rect 35115 17289 35127 17323
rect 35069 17283 35127 17289
rect 36265 17323 36323 17329
rect 36265 17289 36277 17323
rect 36311 17320 36323 17323
rect 36354 17320 36360 17332
rect 36311 17292 36360 17320
rect 36311 17289 36323 17292
rect 36265 17283 36323 17289
rect 36354 17280 36360 17292
rect 36412 17280 36418 17332
rect 38746 17280 38752 17332
rect 38804 17280 38810 17332
rect 38838 17280 38844 17332
rect 38896 17320 38902 17332
rect 39482 17320 39488 17332
rect 38896 17292 39160 17320
rect 38896 17280 38902 17292
rect 35342 17252 35348 17264
rect 32232 17224 35348 17252
rect 28206 17156 29408 17184
rect 29549 17187 29607 17193
rect 28206 17153 28218 17156
rect 28160 17147 28218 17153
rect 29549 17153 29561 17187
rect 29595 17153 29607 17187
rect 29549 17147 29607 17153
rect 30469 17187 30527 17193
rect 30469 17153 30481 17187
rect 30515 17153 30527 17187
rect 30469 17147 30527 17153
rect 27893 17119 27951 17125
rect 27893 17116 27905 17119
rect 27580 17088 27905 17116
rect 27580 17076 27586 17088
rect 27893 17085 27905 17088
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 28902 17076 28908 17128
rect 28960 17116 28966 17128
rect 29564 17116 29592 17147
rect 28960 17088 29592 17116
rect 30484 17116 30512 17147
rect 31570 17144 31576 17196
rect 31628 17144 31634 17196
rect 31665 17187 31723 17193
rect 31665 17153 31677 17187
rect 31711 17184 31723 17187
rect 32030 17184 32036 17196
rect 31711 17156 32036 17184
rect 31711 17153 31723 17156
rect 31665 17147 31723 17153
rect 32030 17144 32036 17156
rect 32088 17144 32094 17196
rect 32232 17193 32260 17224
rect 32217 17187 32275 17193
rect 32217 17153 32229 17187
rect 32263 17153 32275 17187
rect 32217 17147 32275 17153
rect 32484 17187 32542 17193
rect 32484 17153 32496 17187
rect 32530 17184 32542 17187
rect 33226 17184 33232 17196
rect 32530 17156 33232 17184
rect 32530 17153 32542 17156
rect 32484 17147 32542 17153
rect 33226 17144 33232 17156
rect 33284 17144 33290 17196
rect 33704 17193 33732 17224
rect 35342 17212 35348 17224
rect 35400 17212 35406 17264
rect 36081 17255 36139 17261
rect 36081 17221 36093 17255
rect 36127 17252 36139 17255
rect 37826 17252 37832 17264
rect 36127 17224 37832 17252
rect 36127 17221 36139 17224
rect 36081 17215 36139 17221
rect 37826 17212 37832 17224
rect 37884 17212 37890 17264
rect 33962 17193 33968 17196
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17153 33747 17187
rect 33956 17184 33968 17193
rect 33923 17156 33968 17184
rect 33689 17147 33747 17153
rect 33956 17147 33968 17156
rect 33962 17144 33968 17147
rect 34020 17144 34026 17196
rect 35713 17187 35771 17193
rect 35713 17153 35725 17187
rect 35759 17153 35771 17187
rect 35713 17147 35771 17153
rect 31754 17116 31760 17128
rect 30484 17088 31760 17116
rect 28960 17076 28966 17088
rect 31754 17076 31760 17088
rect 31812 17076 31818 17128
rect 31846 17076 31852 17128
rect 31904 17116 31910 17128
rect 35728 17116 35756 17147
rect 35894 17144 35900 17196
rect 35952 17184 35958 17196
rect 36170 17184 36176 17196
rect 35952 17156 36176 17184
rect 35952 17144 35958 17156
rect 36170 17144 36176 17156
rect 36228 17144 36234 17196
rect 36357 17187 36415 17193
rect 36357 17153 36369 17187
rect 36403 17184 36415 17187
rect 36446 17184 36452 17196
rect 36403 17156 36452 17184
rect 36403 17153 36415 17156
rect 36357 17147 36415 17153
rect 36446 17144 36452 17156
rect 36504 17144 36510 17196
rect 38764 17184 38792 17280
rect 39132 17193 39160 17292
rect 39316 17292 39488 17320
rect 39316 17193 39344 17292
rect 39482 17280 39488 17292
rect 39540 17280 39546 17332
rect 41598 17280 41604 17332
rect 41656 17280 41662 17332
rect 44177 17323 44235 17329
rect 44177 17289 44189 17323
rect 44223 17320 44235 17323
rect 44358 17320 44364 17332
rect 44223 17292 44364 17320
rect 44223 17289 44235 17292
rect 44177 17283 44235 17289
rect 44358 17280 44364 17292
rect 44416 17280 44422 17332
rect 46474 17280 46480 17332
rect 46532 17280 46538 17332
rect 46845 17323 46903 17329
rect 46845 17289 46857 17323
rect 46891 17320 46903 17323
rect 47026 17320 47032 17332
rect 46891 17292 47032 17320
rect 46891 17289 46903 17292
rect 46845 17283 46903 17289
rect 47026 17280 47032 17292
rect 47084 17280 47090 17332
rect 39942 17252 39948 17264
rect 39500 17224 39948 17252
rect 39500 17193 39528 17224
rect 39942 17212 39948 17224
rect 40000 17212 40006 17264
rect 38841 17187 38899 17193
rect 38841 17184 38853 17187
rect 38764 17156 38853 17184
rect 38841 17153 38853 17156
rect 38887 17153 38899 17187
rect 38841 17147 38899 17153
rect 39117 17187 39175 17193
rect 39117 17153 39129 17187
rect 39163 17153 39175 17187
rect 39117 17147 39175 17153
rect 39301 17187 39359 17193
rect 39301 17153 39313 17187
rect 39347 17153 39359 17187
rect 39301 17147 39359 17153
rect 39485 17187 39543 17193
rect 39485 17153 39497 17187
rect 39531 17153 39543 17187
rect 39485 17147 39543 17153
rect 39574 17144 39580 17196
rect 39632 17184 39638 17196
rect 39741 17187 39799 17193
rect 39741 17184 39753 17187
rect 39632 17156 39753 17184
rect 39632 17144 39638 17156
rect 39741 17153 39753 17156
rect 39787 17153 39799 17187
rect 39741 17147 39799 17153
rect 43064 17187 43122 17193
rect 43064 17153 43076 17187
rect 43110 17184 43122 17187
rect 43898 17184 43904 17196
rect 43110 17156 43904 17184
rect 43110 17153 43122 17156
rect 43064 17147 43122 17153
rect 43898 17144 43904 17156
rect 43956 17144 43962 17196
rect 45646 17144 45652 17196
rect 45704 17184 45710 17196
rect 46382 17184 46388 17196
rect 45704 17156 46388 17184
rect 45704 17144 45710 17156
rect 46382 17144 46388 17156
rect 46440 17144 46446 17196
rect 46492 17184 46520 17280
rect 50157 17255 50215 17261
rect 50157 17252 50169 17255
rect 49726 17224 50169 17252
rect 50157 17221 50169 17224
rect 50203 17221 50215 17255
rect 50157 17215 50215 17221
rect 46753 17187 46811 17193
rect 46753 17184 46765 17187
rect 46492 17156 46765 17184
rect 46753 17153 46765 17156
rect 46799 17153 46811 17187
rect 50062 17184 50068 17196
rect 46753 17147 46811 17153
rect 49804 17156 50068 17184
rect 38657 17119 38715 17125
rect 31904 17088 32168 17116
rect 35728 17088 36124 17116
rect 31904 17076 31910 17088
rect 32140 17060 32168 17088
rect 32122 17008 32128 17060
rect 32180 17008 32186 17060
rect 36096 17057 36124 17088
rect 38657 17085 38669 17119
rect 38703 17116 38715 17119
rect 38930 17116 38936 17128
rect 38703 17088 38936 17116
rect 38703 17085 38715 17088
rect 38657 17079 38715 17085
rect 38930 17076 38936 17088
rect 38988 17076 38994 17128
rect 40954 17076 40960 17128
rect 41012 17076 41018 17128
rect 42794 17076 42800 17128
rect 42852 17076 42858 17128
rect 44361 17119 44419 17125
rect 44361 17085 44373 17119
rect 44407 17116 44419 17119
rect 46661 17119 46719 17125
rect 46661 17116 46673 17119
rect 44407 17088 46673 17116
rect 44407 17085 44419 17088
rect 44361 17079 44419 17085
rect 46661 17085 46673 17088
rect 46707 17116 46719 17119
rect 47302 17116 47308 17128
rect 46707 17088 47308 17116
rect 46707 17085 46719 17088
rect 46661 17079 46719 17085
rect 36081 17051 36139 17057
rect 34624 17020 36032 17048
rect 25774 16940 25780 16992
rect 25832 16980 25838 16992
rect 25961 16983 26019 16989
rect 25961 16980 25973 16983
rect 25832 16952 25973 16980
rect 25832 16940 25838 16952
rect 25961 16949 25973 16952
rect 26007 16949 26019 16983
rect 25961 16943 26019 16949
rect 28810 16940 28816 16992
rect 28868 16980 28874 16992
rect 29273 16983 29331 16989
rect 29273 16980 29285 16983
rect 28868 16952 29285 16980
rect 28868 16940 28874 16952
rect 29273 16949 29285 16952
rect 29319 16949 29331 16983
rect 29273 16943 29331 16949
rect 30282 16940 30288 16992
rect 30340 16940 30346 16992
rect 30374 16940 30380 16992
rect 30432 16980 30438 16992
rect 34624 16980 34652 17020
rect 30432 16952 34652 16980
rect 30432 16940 30438 16952
rect 35618 16940 35624 16992
rect 35676 16980 35682 16992
rect 35713 16983 35771 16989
rect 35713 16980 35725 16983
rect 35676 16952 35725 16980
rect 35676 16940 35682 16952
rect 35713 16949 35725 16952
rect 35759 16949 35771 16983
rect 36004 16980 36032 17020
rect 36081 17017 36093 17051
rect 36127 17017 36139 17051
rect 41230 17048 41236 17060
rect 36081 17011 36139 17017
rect 40420 17020 41236 17048
rect 40420 16980 40448 17020
rect 41230 17008 41236 17020
rect 41288 17008 41294 17060
rect 36004 16952 40448 16980
rect 35713 16943 35771 16949
rect 40862 16940 40868 16992
rect 40920 16980 40926 16992
rect 44376 16980 44404 17079
rect 47302 17076 47308 17088
rect 47360 17076 47366 17128
rect 48222 17076 48228 17128
rect 48280 17076 48286 17128
rect 48498 17076 48504 17128
rect 48556 17076 48562 17128
rect 49804 17060 49832 17156
rect 50062 17144 50068 17156
rect 50120 17144 50126 17196
rect 46566 17048 46572 17060
rect 45940 17020 46572 17048
rect 45940 16992 45968 17020
rect 46566 17008 46572 17020
rect 46624 17008 46630 17060
rect 49786 17008 49792 17060
rect 49844 17008 49850 17060
rect 68462 17008 68468 17060
rect 68520 17008 68526 17060
rect 40920 16952 44404 16980
rect 40920 16940 40926 16952
rect 44910 16940 44916 16992
rect 44968 16940 44974 16992
rect 45922 16940 45928 16992
rect 45980 16940 45986 16992
rect 46198 16940 46204 16992
rect 46256 16940 46262 16992
rect 49234 16940 49240 16992
rect 49292 16980 49298 16992
rect 49973 16983 50031 16989
rect 49973 16980 49985 16983
rect 49292 16952 49985 16980
rect 49292 16940 49298 16952
rect 49973 16949 49985 16952
rect 50019 16949 50031 16983
rect 49973 16943 50031 16949
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 28169 16779 28227 16785
rect 28169 16745 28181 16779
rect 28215 16776 28227 16779
rect 28718 16776 28724 16788
rect 28215 16748 28724 16776
rect 28215 16745 28227 16748
rect 28169 16739 28227 16745
rect 28718 16736 28724 16748
rect 28776 16736 28782 16788
rect 28810 16736 28816 16788
rect 28868 16736 28874 16788
rect 33042 16736 33048 16788
rect 33100 16776 33106 16788
rect 33100 16748 37320 16776
rect 33100 16736 33106 16748
rect 27525 16643 27583 16649
rect 27525 16609 27537 16643
rect 27571 16640 27583 16643
rect 28445 16643 28503 16649
rect 27571 16612 28396 16640
rect 27571 16609 27583 16612
rect 27525 16603 27583 16609
rect 25222 16532 25228 16584
rect 25280 16572 25286 16584
rect 25774 16581 25780 16584
rect 25501 16575 25559 16581
rect 25501 16572 25513 16575
rect 25280 16544 25513 16572
rect 25280 16532 25286 16544
rect 25501 16541 25513 16544
rect 25547 16541 25559 16575
rect 25768 16572 25780 16581
rect 25735 16544 25780 16572
rect 25501 16535 25559 16541
rect 25768 16535 25780 16544
rect 25774 16532 25780 16535
rect 25832 16532 25838 16584
rect 27801 16575 27859 16581
rect 27801 16572 27813 16575
rect 27448 16544 27813 16572
rect 27448 16513 27476 16544
rect 27801 16541 27813 16544
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 27982 16532 27988 16584
rect 28040 16532 28046 16584
rect 27433 16507 27491 16513
rect 27433 16504 27445 16507
rect 26896 16476 27445 16504
rect 26896 16448 26924 16476
rect 27433 16473 27445 16476
rect 27479 16473 27491 16507
rect 28368 16504 28396 16612
rect 28445 16609 28457 16643
rect 28491 16640 28503 16643
rect 28828 16640 28856 16736
rect 36725 16711 36783 16717
rect 36725 16677 36737 16711
rect 36771 16708 36783 16711
rect 37292 16708 37320 16748
rect 37826 16736 37832 16788
rect 37884 16736 37890 16788
rect 39390 16736 39396 16788
rect 39448 16776 39454 16788
rect 39485 16779 39543 16785
rect 39485 16776 39497 16779
rect 39448 16748 39497 16776
rect 39448 16736 39454 16748
rect 39485 16745 39497 16748
rect 39531 16745 39543 16779
rect 44821 16779 44879 16785
rect 44821 16776 44833 16779
rect 39485 16739 39543 16745
rect 39592 16748 44833 16776
rect 39592 16708 39620 16748
rect 44821 16745 44833 16748
rect 44867 16745 44879 16779
rect 45922 16776 45928 16788
rect 44821 16739 44879 16745
rect 44928 16748 45928 16776
rect 36771 16680 37228 16708
rect 37292 16680 38700 16708
rect 36771 16677 36783 16680
rect 36725 16671 36783 16677
rect 28491 16612 28856 16640
rect 28491 16609 28503 16612
rect 28445 16603 28503 16609
rect 29178 16600 29184 16652
rect 29236 16640 29242 16652
rect 37200 16649 37228 16680
rect 38672 16649 38700 16680
rect 38856 16680 39620 16708
rect 39669 16711 39727 16717
rect 29733 16643 29791 16649
rect 29733 16640 29745 16643
rect 29236 16612 29745 16640
rect 29236 16600 29242 16612
rect 29472 16584 29500 16612
rect 29733 16609 29745 16612
rect 29779 16609 29791 16643
rect 29733 16603 29791 16609
rect 37185 16643 37243 16649
rect 37185 16609 37197 16643
rect 37231 16609 37243 16643
rect 37185 16603 37243 16609
rect 38657 16643 38715 16649
rect 38657 16609 38669 16643
rect 38703 16609 38715 16643
rect 38657 16603 38715 16609
rect 28718 16532 28724 16584
rect 28776 16572 28782 16584
rect 29273 16575 29331 16581
rect 29273 16572 29285 16575
rect 28776 16544 29285 16572
rect 28776 16532 28782 16544
rect 29273 16541 29285 16544
rect 29319 16541 29331 16575
rect 29273 16535 29331 16541
rect 29365 16575 29423 16581
rect 29365 16541 29377 16575
rect 29411 16541 29423 16575
rect 29365 16535 29423 16541
rect 28902 16504 28908 16516
rect 28368 16476 28908 16504
rect 27433 16467 27491 16473
rect 28902 16464 28908 16476
rect 28960 16464 28966 16516
rect 28997 16507 29055 16513
rect 28997 16473 29009 16507
rect 29043 16504 29055 16507
rect 29089 16507 29147 16513
rect 29089 16504 29101 16507
rect 29043 16476 29101 16504
rect 29043 16473 29055 16476
rect 28997 16467 29055 16473
rect 29089 16473 29101 16476
rect 29135 16473 29147 16507
rect 29089 16467 29147 16473
rect 29380 16448 29408 16535
rect 29454 16532 29460 16584
rect 29512 16532 29518 16584
rect 30000 16575 30058 16581
rect 30000 16541 30012 16575
rect 30046 16572 30058 16575
rect 30282 16572 30288 16584
rect 30046 16544 30288 16572
rect 30046 16541 30058 16544
rect 30000 16535 30058 16541
rect 30282 16532 30288 16544
rect 30340 16532 30346 16584
rect 35618 16581 35624 16584
rect 35345 16575 35403 16581
rect 35345 16541 35357 16575
rect 35391 16541 35403 16575
rect 35612 16572 35624 16581
rect 35579 16544 35624 16572
rect 35345 16535 35403 16541
rect 35612 16535 35624 16544
rect 35360 16448 35388 16535
rect 35618 16532 35624 16535
rect 35676 16532 35682 16584
rect 38856 16581 38884 16680
rect 39669 16677 39681 16711
rect 39715 16677 39727 16711
rect 39669 16671 39727 16677
rect 39853 16711 39911 16717
rect 39853 16677 39865 16711
rect 39899 16708 39911 16711
rect 41509 16711 41567 16717
rect 39899 16680 40172 16708
rect 39899 16677 39911 16680
rect 39853 16671 39911 16677
rect 39117 16643 39175 16649
rect 39117 16609 39129 16643
rect 39163 16640 39175 16643
rect 39684 16640 39712 16671
rect 40144 16640 40172 16680
rect 41509 16677 41521 16711
rect 41555 16677 41567 16711
rect 43162 16708 43168 16720
rect 41509 16671 41567 16677
rect 42536 16680 43168 16708
rect 41524 16640 41552 16671
rect 41601 16643 41659 16649
rect 41601 16640 41613 16643
rect 39163 16612 39620 16640
rect 39684 16612 39896 16640
rect 40144 16612 40264 16640
rect 41524 16612 41613 16640
rect 39163 16609 39175 16612
rect 39117 16603 39175 16609
rect 38105 16575 38163 16581
rect 38105 16572 38117 16575
rect 38028 16544 38117 16572
rect 38028 16448 38056 16544
rect 38105 16541 38117 16544
rect 38151 16541 38163 16575
rect 38105 16535 38163 16541
rect 38841 16575 38899 16581
rect 38841 16541 38853 16575
rect 38887 16541 38899 16575
rect 38841 16535 38899 16541
rect 38194 16464 38200 16516
rect 38252 16464 38258 16516
rect 26878 16396 26884 16448
rect 26936 16396 26942 16448
rect 26970 16396 26976 16448
rect 27028 16396 27034 16448
rect 27338 16396 27344 16448
rect 27396 16396 27402 16448
rect 28626 16396 28632 16448
rect 28684 16436 28690 16448
rect 29187 16439 29245 16445
rect 29187 16436 29199 16439
rect 28684 16408 29199 16436
rect 28684 16396 28690 16408
rect 29187 16405 29199 16408
rect 29233 16405 29245 16439
rect 29187 16399 29245 16405
rect 29362 16396 29368 16448
rect 29420 16396 29426 16448
rect 30282 16396 30288 16448
rect 30340 16436 30346 16448
rect 31113 16439 31171 16445
rect 31113 16436 31125 16439
rect 30340 16408 31125 16436
rect 30340 16396 30346 16408
rect 31113 16405 31125 16408
rect 31159 16405 31171 16439
rect 31113 16399 31171 16405
rect 35342 16396 35348 16448
rect 35400 16396 35406 16448
rect 38010 16396 38016 16448
rect 38068 16396 38074 16448
rect 39022 16396 39028 16448
rect 39080 16396 39086 16448
rect 39482 16396 39488 16448
rect 39540 16396 39546 16448
rect 39592 16436 39620 16612
rect 39868 16572 39896 16612
rect 40037 16575 40095 16581
rect 40037 16572 40049 16575
rect 39868 16544 40049 16572
rect 40037 16541 40049 16544
rect 40083 16541 40095 16575
rect 40037 16535 40095 16541
rect 40129 16575 40187 16581
rect 40129 16541 40141 16575
rect 40175 16541 40187 16575
rect 40129 16535 40187 16541
rect 39942 16464 39948 16516
rect 40000 16504 40006 16516
rect 40144 16504 40172 16535
rect 40000 16476 40172 16504
rect 40236 16504 40264 16612
rect 41601 16609 41613 16612
rect 41647 16609 41659 16643
rect 41601 16603 41659 16609
rect 42429 16575 42487 16581
rect 42429 16541 42441 16575
rect 42475 16572 42487 16575
rect 42536 16572 42564 16680
rect 43162 16668 43168 16680
rect 43220 16668 43226 16720
rect 44177 16711 44235 16717
rect 44177 16677 44189 16711
rect 44223 16708 44235 16711
rect 44928 16708 44956 16748
rect 45922 16736 45928 16748
rect 45980 16736 45986 16788
rect 46198 16736 46204 16788
rect 46256 16736 46262 16788
rect 48225 16779 48283 16785
rect 48225 16745 48237 16779
rect 48271 16776 48283 16779
rect 48498 16776 48504 16788
rect 48271 16748 48504 16776
rect 48271 16745 48283 16748
rect 48225 16739 48283 16745
rect 48498 16736 48504 16748
rect 48556 16736 48562 16788
rect 48774 16736 48780 16788
rect 48832 16776 48838 16788
rect 49145 16779 49203 16785
rect 49145 16776 49157 16779
rect 48832 16748 49157 16776
rect 48832 16736 48838 16748
rect 49145 16745 49157 16748
rect 49191 16745 49203 16779
rect 49145 16739 49203 16745
rect 44223 16680 44956 16708
rect 45005 16711 45063 16717
rect 44223 16677 44235 16680
rect 44177 16671 44235 16677
rect 45005 16677 45017 16711
rect 45051 16677 45063 16711
rect 45005 16671 45063 16677
rect 42610 16600 42616 16652
rect 42668 16640 42674 16652
rect 42797 16643 42855 16649
rect 42797 16640 42809 16643
rect 42668 16612 42809 16640
rect 42668 16600 42674 16612
rect 42797 16609 42809 16612
rect 42843 16609 42855 16643
rect 42797 16603 42855 16609
rect 43625 16643 43683 16649
rect 43625 16609 43637 16643
rect 43671 16640 43683 16643
rect 44082 16640 44088 16652
rect 43671 16612 44088 16640
rect 43671 16609 43683 16612
rect 43625 16603 43683 16609
rect 44082 16600 44088 16612
rect 44140 16600 44146 16652
rect 44192 16612 44404 16640
rect 42475 16544 42564 16572
rect 42705 16575 42763 16581
rect 42475 16541 42487 16544
rect 42429 16535 42487 16541
rect 42705 16541 42717 16575
rect 42751 16541 42763 16575
rect 42705 16535 42763 16541
rect 40374 16507 40432 16513
rect 40374 16504 40386 16507
rect 40236 16476 40386 16504
rect 40000 16464 40006 16476
rect 40374 16473 40386 16476
rect 40420 16473 40432 16507
rect 42720 16504 42748 16535
rect 43806 16532 43812 16584
rect 43864 16572 43870 16584
rect 44192 16572 44220 16612
rect 43864 16544 44220 16572
rect 43864 16532 43870 16544
rect 44266 16532 44272 16584
rect 44324 16532 44330 16584
rect 44376 16572 44404 16612
rect 44637 16575 44695 16581
rect 44637 16572 44649 16575
rect 44376 16544 44649 16572
rect 44637 16541 44649 16544
rect 44683 16541 44695 16575
rect 45020 16572 45048 16671
rect 46109 16643 46167 16649
rect 46109 16609 46121 16643
rect 46155 16640 46167 16643
rect 46216 16640 46244 16736
rect 48133 16711 48191 16717
rect 48133 16677 48145 16711
rect 48179 16708 48191 16711
rect 48179 16680 48544 16708
rect 48179 16677 48191 16680
rect 48133 16671 48191 16677
rect 46658 16640 46664 16652
rect 46155 16612 46244 16640
rect 46584 16612 46664 16640
rect 46155 16609 46167 16612
rect 46109 16603 46167 16609
rect 44637 16535 44695 16541
rect 44744 16544 45048 16572
rect 45281 16575 45339 16581
rect 42886 16504 42892 16516
rect 42720 16476 42892 16504
rect 40374 16467 40432 16473
rect 42886 16464 42892 16476
rect 42944 16464 42950 16516
rect 44453 16507 44511 16513
rect 43364 16476 44312 16504
rect 40218 16436 40224 16448
rect 39592 16408 40224 16436
rect 40218 16396 40224 16408
rect 40276 16396 40282 16448
rect 42242 16396 42248 16448
rect 42300 16396 42306 16448
rect 42518 16396 42524 16448
rect 42576 16445 42582 16448
rect 42576 16399 42585 16445
rect 42613 16439 42671 16445
rect 42613 16405 42625 16439
rect 42659 16436 42671 16439
rect 43364 16436 43392 16476
rect 44284 16448 44312 16476
rect 44453 16473 44465 16507
rect 44499 16473 44511 16507
rect 44453 16467 44511 16473
rect 42659 16408 43392 16436
rect 42659 16405 42671 16408
rect 42613 16399 42671 16405
rect 42576 16396 42582 16399
rect 43438 16396 43444 16448
rect 43496 16396 43502 16448
rect 44266 16396 44272 16448
rect 44324 16396 44330 16448
rect 44468 16436 44496 16467
rect 44542 16464 44548 16516
rect 44600 16464 44606 16516
rect 44744 16448 44772 16544
rect 45281 16541 45293 16575
rect 45327 16541 45339 16575
rect 45281 16535 45339 16541
rect 45002 16464 45008 16516
rect 45060 16464 45066 16516
rect 45296 16504 45324 16535
rect 45370 16532 45376 16584
rect 45428 16532 45434 16584
rect 45557 16575 45615 16581
rect 45557 16541 45569 16575
rect 45603 16572 45615 16575
rect 46584 16572 46612 16612
rect 46658 16600 46664 16612
rect 46716 16600 46722 16652
rect 48516 16649 48544 16680
rect 48501 16643 48559 16649
rect 48501 16609 48513 16643
rect 48547 16609 48559 16643
rect 48501 16603 48559 16609
rect 48774 16600 48780 16652
rect 48832 16640 48838 16652
rect 49234 16640 49240 16652
rect 48832 16612 49240 16640
rect 48832 16600 48838 16612
rect 49234 16600 49240 16612
rect 49292 16600 49298 16652
rect 45603 16544 46612 16572
rect 45603 16541 45615 16544
rect 45557 16535 45615 16541
rect 45664 16516 45692 16544
rect 46750 16532 46756 16584
rect 46808 16532 46814 16584
rect 48406 16532 48412 16584
rect 48464 16532 48470 16584
rect 51261 16575 51319 16581
rect 51261 16541 51273 16575
rect 51307 16541 51319 16575
rect 51261 16535 51319 16541
rect 45465 16507 45523 16513
rect 45465 16504 45477 16507
rect 45296 16476 45477 16504
rect 45465 16473 45477 16476
rect 45511 16473 45523 16507
rect 45465 16467 45523 16473
rect 45646 16464 45652 16516
rect 45704 16464 45710 16516
rect 46661 16507 46719 16513
rect 46661 16473 46673 16507
rect 46707 16504 46719 16507
rect 46998 16507 47056 16513
rect 46998 16504 47010 16507
rect 46707 16476 47010 16504
rect 46707 16473 46719 16476
rect 46661 16467 46719 16473
rect 46998 16473 47010 16476
rect 47044 16473 47056 16507
rect 46998 16467 47056 16473
rect 49786 16464 49792 16516
rect 49844 16504 49850 16516
rect 51276 16504 51304 16535
rect 51810 16532 51816 16584
rect 51868 16532 51874 16584
rect 49844 16476 52776 16504
rect 49844 16464 49850 16476
rect 52748 16448 52776 16476
rect 44634 16436 44640 16448
rect 44468 16408 44640 16436
rect 44634 16396 44640 16408
rect 44692 16396 44698 16448
rect 44726 16396 44732 16448
rect 44784 16396 44790 16448
rect 45186 16396 45192 16448
rect 45244 16396 45250 16448
rect 49694 16396 49700 16448
rect 49752 16436 49758 16448
rect 49881 16439 49939 16445
rect 49881 16436 49893 16439
rect 49752 16408 49893 16436
rect 49752 16396 49758 16408
rect 49881 16405 49893 16408
rect 49927 16405 49939 16439
rect 49881 16399 49939 16405
rect 51353 16439 51411 16445
rect 51353 16405 51365 16439
rect 51399 16436 51411 16439
rect 51442 16436 51448 16448
rect 51399 16408 51448 16436
rect 51399 16405 51411 16408
rect 51353 16399 51411 16405
rect 51442 16396 51448 16408
rect 51500 16396 51506 16448
rect 52362 16396 52368 16448
rect 52420 16396 52426 16448
rect 52730 16396 52736 16448
rect 52788 16396 52794 16448
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 26252 16204 26464 16232
rect 25961 16167 26019 16173
rect 25961 16133 25973 16167
rect 26007 16164 26019 16167
rect 26142 16164 26148 16176
rect 26007 16136 26148 16164
rect 26007 16133 26019 16136
rect 25961 16127 26019 16133
rect 26142 16124 26148 16136
rect 26200 16124 26206 16176
rect 25777 16099 25835 16105
rect 25777 16065 25789 16099
rect 25823 16065 25835 16099
rect 25777 16059 25835 16065
rect 25792 16028 25820 16059
rect 26050 16056 26056 16108
rect 26108 16056 26114 16108
rect 26142 16028 26148 16040
rect 25792 16000 26148 16028
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 26252 16037 26280 16204
rect 26436 16164 26464 16204
rect 26602 16192 26608 16244
rect 26660 16192 26666 16244
rect 26694 16192 26700 16244
rect 26752 16192 26758 16244
rect 26970 16192 26976 16244
rect 27028 16192 27034 16244
rect 27338 16192 27344 16244
rect 27396 16192 27402 16244
rect 27982 16192 27988 16244
rect 28040 16232 28046 16244
rect 28902 16232 28908 16244
rect 28040 16204 28908 16232
rect 28040 16192 28046 16204
rect 28902 16192 28908 16204
rect 28960 16232 28966 16244
rect 29181 16235 29239 16241
rect 29181 16232 29193 16235
rect 28960 16204 29193 16232
rect 28960 16192 28966 16204
rect 29181 16201 29193 16204
rect 29227 16201 29239 16235
rect 29181 16195 29239 16201
rect 29362 16192 29368 16244
rect 29420 16232 29426 16244
rect 29420 16204 29592 16232
rect 29420 16192 29426 16204
rect 26712 16164 26740 16192
rect 26436 16136 26740 16164
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16096 26479 16099
rect 26988 16096 27016 16192
rect 27356 16164 27384 16192
rect 27356 16136 29500 16164
rect 26467 16068 27016 16096
rect 27792 16099 27850 16105
rect 26467 16065 26479 16068
rect 26421 16059 26479 16065
rect 27792 16065 27804 16099
rect 27838 16096 27850 16099
rect 28810 16096 28816 16108
rect 27838 16068 28816 16096
rect 27838 16065 27850 16068
rect 27792 16059 27850 16065
rect 28810 16056 28816 16068
rect 28868 16056 28874 16108
rect 29089 16099 29147 16105
rect 29089 16096 29101 16099
rect 29012 16068 29101 16096
rect 29012 16040 29040 16068
rect 29089 16065 29101 16068
rect 29135 16065 29147 16099
rect 29089 16059 29147 16065
rect 29270 16056 29276 16108
rect 29328 16056 29334 16108
rect 29472 16105 29500 16136
rect 29457 16099 29515 16105
rect 29457 16065 29469 16099
rect 29503 16065 29515 16099
rect 29564 16096 29592 16204
rect 30006 16192 30012 16244
rect 30064 16232 30070 16244
rect 30064 16204 31524 16232
rect 30064 16192 30070 16204
rect 31496 16176 31524 16204
rect 31754 16192 31760 16244
rect 31812 16232 31818 16244
rect 32493 16235 32551 16241
rect 32493 16232 32505 16235
rect 31812 16204 32505 16232
rect 31812 16192 31818 16204
rect 32493 16201 32505 16204
rect 32539 16201 32551 16235
rect 32493 16195 32551 16201
rect 39942 16192 39948 16244
rect 40000 16192 40006 16244
rect 40862 16192 40868 16244
rect 40920 16192 40926 16244
rect 42242 16232 42248 16244
rect 41386 16204 42248 16232
rect 30837 16167 30895 16173
rect 30837 16164 30849 16167
rect 30668 16136 30849 16164
rect 30668 16108 30696 16136
rect 30837 16133 30849 16136
rect 30883 16133 30895 16167
rect 30837 16127 30895 16133
rect 31478 16124 31484 16176
rect 31536 16164 31542 16176
rect 37553 16167 37611 16173
rect 31536 16136 37136 16164
rect 31536 16124 31542 16136
rect 30561 16099 30619 16105
rect 30561 16096 30573 16099
rect 29564 16068 30573 16096
rect 29457 16059 29515 16065
rect 30561 16065 30573 16068
rect 30607 16065 30619 16099
rect 30561 16059 30619 16065
rect 26237 16031 26295 16037
rect 26237 15997 26249 16031
rect 26283 15997 26295 16031
rect 26237 15991 26295 15997
rect 27522 15988 27528 16040
rect 27580 15988 27586 16040
rect 28994 15988 29000 16040
rect 29052 16028 29058 16040
rect 29362 16028 29368 16040
rect 29052 16000 29368 16028
rect 29052 15988 29058 16000
rect 29362 15988 29368 16000
rect 29420 15988 29426 16040
rect 29472 16028 29500 16059
rect 30650 16056 30656 16108
rect 30708 16056 30714 16108
rect 30745 16099 30803 16105
rect 30745 16065 30757 16099
rect 30791 16065 30803 16099
rect 30745 16059 30803 16065
rect 30929 16099 30987 16105
rect 30929 16065 30941 16099
rect 30975 16096 30987 16099
rect 31110 16096 31116 16108
rect 30975 16068 31116 16096
rect 30975 16065 30987 16068
rect 30929 16059 30987 16065
rect 29914 16028 29920 16040
rect 29472 16000 29920 16028
rect 29914 15988 29920 16000
rect 29972 16028 29978 16040
rect 30282 16028 30288 16040
rect 29972 16000 30288 16028
rect 29972 15988 29978 16000
rect 30282 15988 30288 16000
rect 30340 16028 30346 16040
rect 30760 16028 30788 16059
rect 31110 16056 31116 16068
rect 31168 16056 31174 16108
rect 32309 16099 32367 16105
rect 32309 16096 32321 16099
rect 31726 16068 32321 16096
rect 30340 16000 30788 16028
rect 30340 15988 30346 16000
rect 31202 15988 31208 16040
rect 31260 15988 31266 16040
rect 25222 15920 25228 15972
rect 25280 15960 25286 15972
rect 27540 15960 27568 15988
rect 25280 15932 27568 15960
rect 25280 15920 25286 15932
rect 28534 15920 28540 15972
rect 28592 15960 28598 15972
rect 30101 15963 30159 15969
rect 30101 15960 30113 15963
rect 28592 15932 30113 15960
rect 28592 15920 28598 15932
rect 30101 15929 30113 15932
rect 30147 15929 30159 15963
rect 30101 15923 30159 15929
rect 31113 15963 31171 15969
rect 31113 15929 31125 15963
rect 31159 15960 31171 15963
rect 31726 15960 31754 16068
rect 32309 16065 32321 16068
rect 32355 16065 32367 16099
rect 32309 16059 32367 16065
rect 33042 16056 33048 16108
rect 33100 16056 33106 16108
rect 33321 16099 33379 16105
rect 33321 16065 33333 16099
rect 33367 16065 33379 16099
rect 33321 16059 33379 16065
rect 32122 15988 32128 16040
rect 32180 16028 32186 16040
rect 33060 16028 33088 16056
rect 32180 16000 33088 16028
rect 32180 15988 32186 16000
rect 31159 15932 31754 15960
rect 33336 15960 33364 16059
rect 33410 16056 33416 16108
rect 33468 16056 33474 16108
rect 33612 16105 33640 16136
rect 37108 16108 37136 16136
rect 37553 16133 37565 16167
rect 37599 16164 37611 16167
rect 37826 16164 37832 16176
rect 37599 16136 37832 16164
rect 37599 16133 37611 16136
rect 37553 16127 37611 16133
rect 37826 16124 37832 16136
rect 37884 16124 37890 16176
rect 38102 16124 38108 16176
rect 38160 16124 38166 16176
rect 39960 16164 39988 16192
rect 39132 16136 39988 16164
rect 33597 16099 33655 16105
rect 33597 16065 33609 16099
rect 33643 16065 33655 16099
rect 33597 16059 33655 16065
rect 33689 16099 33747 16105
rect 33689 16065 33701 16099
rect 33735 16096 33747 16099
rect 34425 16099 34483 16105
rect 34425 16096 34437 16099
rect 33735 16068 34437 16096
rect 33735 16065 33747 16068
rect 33689 16059 33747 16065
rect 34425 16065 34437 16068
rect 34471 16096 34483 16099
rect 34514 16096 34520 16108
rect 34471 16068 34520 16096
rect 34471 16065 34483 16068
rect 34425 16059 34483 16065
rect 34514 16056 34520 16068
rect 34572 16056 34578 16108
rect 37090 16056 37096 16108
rect 37148 16056 37154 16108
rect 39132 16105 39160 16136
rect 39390 16105 39396 16108
rect 39117 16099 39175 16105
rect 39117 16065 39129 16099
rect 39163 16065 39175 16099
rect 39117 16059 39175 16065
rect 39384 16059 39396 16105
rect 39390 16056 39396 16059
rect 39448 16056 39454 16108
rect 39960 16096 39988 16136
rect 40681 16167 40739 16173
rect 40681 16133 40693 16167
rect 40727 16164 40739 16167
rect 41386 16164 41414 16204
rect 42242 16192 42248 16204
rect 42300 16192 42306 16244
rect 42518 16192 42524 16244
rect 42576 16232 42582 16244
rect 42576 16204 43576 16232
rect 42576 16192 42582 16204
rect 42794 16164 42800 16176
rect 40727 16136 41414 16164
rect 42444 16136 42800 16164
rect 40727 16133 40739 16136
rect 40681 16127 40739 16133
rect 39960 16068 40172 16096
rect 33778 15988 33784 16040
rect 33836 15988 33842 16040
rect 37274 15988 37280 16040
rect 37332 15988 37338 16040
rect 40144 16028 40172 16068
rect 40218 16056 40224 16108
rect 40276 16096 40282 16108
rect 40957 16099 41015 16105
rect 40957 16096 40969 16099
rect 40276 16068 40969 16096
rect 40276 16056 40282 16068
rect 40957 16065 40969 16068
rect 41003 16096 41015 16099
rect 41046 16096 41052 16108
rect 41003 16068 41052 16096
rect 41003 16065 41015 16068
rect 40957 16059 41015 16065
rect 41046 16056 41052 16068
rect 41104 16056 41110 16108
rect 42444 16105 42472 16136
rect 42794 16124 42800 16136
rect 42852 16124 42858 16176
rect 43438 16124 43444 16176
rect 43496 16124 43502 16176
rect 42429 16099 42487 16105
rect 42429 16096 42441 16099
rect 41386 16068 42441 16096
rect 41386 16028 41414 16068
rect 42429 16065 42441 16068
rect 42475 16065 42487 16099
rect 42429 16059 42487 16065
rect 42696 16099 42754 16105
rect 42696 16065 42708 16099
rect 42742 16096 42754 16099
rect 43456 16096 43484 16124
rect 42742 16068 43484 16096
rect 43548 16096 43576 16204
rect 43898 16192 43904 16244
rect 43956 16232 43962 16244
rect 43993 16235 44051 16241
rect 43993 16232 44005 16235
rect 43956 16204 44005 16232
rect 43956 16192 43962 16204
rect 43993 16201 44005 16204
rect 44039 16201 44051 16235
rect 43993 16195 44051 16201
rect 44082 16192 44088 16244
rect 44140 16232 44146 16244
rect 44634 16232 44640 16244
rect 44140 16204 44640 16232
rect 44140 16192 44146 16204
rect 44634 16192 44640 16204
rect 44692 16192 44698 16244
rect 44910 16192 44916 16244
rect 44968 16232 44974 16244
rect 44968 16204 46060 16232
rect 44968 16192 44974 16204
rect 44100 16164 44128 16192
rect 44008 16136 44128 16164
rect 43901 16099 43959 16105
rect 43901 16096 43913 16099
rect 43548 16068 43913 16096
rect 42742 16065 42754 16068
rect 42696 16059 42754 16065
rect 43901 16065 43913 16068
rect 43947 16065 43959 16099
rect 43901 16059 43959 16065
rect 40144 16000 41414 16028
rect 34606 15960 34612 15972
rect 33336 15932 34612 15960
rect 31159 15929 31171 15932
rect 31113 15923 31171 15929
rect 34606 15920 34612 15932
rect 34664 15920 34670 15972
rect 40681 15963 40739 15969
rect 40681 15929 40693 15963
rect 40727 15960 40739 15963
rect 40954 15960 40960 15972
rect 40727 15932 40960 15960
rect 40727 15929 40739 15932
rect 40681 15923 40739 15929
rect 40954 15920 40960 15932
rect 41012 15920 41018 15972
rect 44008 15960 44036 16136
rect 44726 16124 44732 16176
rect 44784 16124 44790 16176
rect 45738 16124 45744 16176
rect 45796 16124 45802 16176
rect 44082 16056 44088 16108
rect 44140 16056 44146 16108
rect 44450 15988 44456 16040
rect 44508 15988 44514 16040
rect 46032 16028 46060 16204
rect 51810 16192 51816 16244
rect 51868 16232 51874 16244
rect 51905 16235 51963 16241
rect 51905 16232 51917 16235
rect 51868 16204 51917 16232
rect 51868 16192 51874 16204
rect 51905 16201 51917 16204
rect 51951 16201 51963 16235
rect 51905 16195 51963 16201
rect 51442 16124 51448 16176
rect 51500 16124 51506 16176
rect 46474 16056 46480 16108
rect 46532 16056 46538 16108
rect 46566 16056 46572 16108
rect 46624 16096 46630 16108
rect 47029 16099 47087 16105
rect 47029 16096 47041 16099
rect 46624 16068 47041 16096
rect 46624 16056 46630 16068
rect 47029 16065 47041 16068
rect 47075 16065 47087 16099
rect 47029 16059 47087 16065
rect 47213 16099 47271 16105
rect 47213 16065 47225 16099
rect 47259 16096 47271 16099
rect 48498 16096 48504 16108
rect 47259 16068 48504 16096
rect 47259 16065 47271 16068
rect 47213 16059 47271 16065
rect 48498 16056 48504 16068
rect 48556 16056 48562 16108
rect 46753 16031 46811 16037
rect 46753 16028 46765 16031
rect 46032 16000 46765 16028
rect 46753 15997 46765 16000
rect 46799 15997 46811 16031
rect 46753 15991 46811 15997
rect 50157 16031 50215 16037
rect 50157 15997 50169 16031
rect 50203 15997 50215 16031
rect 50157 15991 50215 15997
rect 43732 15932 44036 15960
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 992 15864 1593 15892
rect 992 15852 998 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 24854 15852 24860 15904
rect 24912 15892 24918 15904
rect 25777 15895 25835 15901
rect 25777 15892 25789 15895
rect 24912 15864 25789 15892
rect 24912 15852 24918 15864
rect 25777 15861 25789 15864
rect 25823 15861 25835 15895
rect 25777 15855 25835 15861
rect 28718 15852 28724 15904
rect 28776 15892 28782 15904
rect 28905 15895 28963 15901
rect 28905 15892 28917 15895
rect 28776 15864 28917 15892
rect 28776 15852 28782 15864
rect 28905 15861 28917 15864
rect 28951 15861 28963 15895
rect 28905 15855 28963 15861
rect 31846 15852 31852 15904
rect 31904 15852 31910 15904
rect 33134 15852 33140 15904
rect 33192 15852 33198 15904
rect 38654 15852 38660 15904
rect 38712 15892 38718 15904
rect 39025 15895 39083 15901
rect 39025 15892 39037 15895
rect 38712 15864 39037 15892
rect 38712 15852 38718 15864
rect 39025 15861 39037 15864
rect 39071 15861 39083 15895
rect 39025 15855 39083 15861
rect 39482 15852 39488 15904
rect 39540 15892 39546 15904
rect 40497 15895 40555 15901
rect 40497 15892 40509 15895
rect 39540 15864 40509 15892
rect 39540 15852 39546 15864
rect 40497 15861 40509 15864
rect 40543 15892 40555 15895
rect 43732 15892 43760 15932
rect 40543 15864 43760 15892
rect 40543 15861 40555 15864
rect 40497 15855 40555 15861
rect 43806 15852 43812 15904
rect 43864 15852 43870 15904
rect 45738 15852 45744 15904
rect 45796 15892 45802 15904
rect 46201 15895 46259 15901
rect 46201 15892 46213 15895
rect 45796 15864 46213 15892
rect 45796 15852 45802 15864
rect 46201 15861 46213 15864
rect 46247 15861 46259 15895
rect 46201 15855 46259 15861
rect 46290 15852 46296 15904
rect 46348 15852 46354 15904
rect 46661 15895 46719 15901
rect 46661 15861 46673 15895
rect 46707 15892 46719 15895
rect 47029 15895 47087 15901
rect 47029 15892 47041 15895
rect 46707 15864 47041 15892
rect 46707 15861 46719 15864
rect 46661 15855 46719 15861
rect 47029 15861 47041 15864
rect 47075 15861 47087 15895
rect 47029 15855 47087 15861
rect 48222 15852 48228 15904
rect 48280 15892 48286 15904
rect 48958 15892 48964 15904
rect 48280 15864 48964 15892
rect 48280 15852 48286 15864
rect 48958 15852 48964 15864
rect 49016 15892 49022 15904
rect 50172 15892 50200 15991
rect 50430 15988 50436 16040
rect 50488 15988 50494 16040
rect 52270 15892 52276 15904
rect 49016 15864 52276 15892
rect 49016 15852 49022 15864
rect 52270 15852 52276 15864
rect 52328 15852 52334 15904
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 26050 15648 26056 15700
rect 26108 15688 26114 15700
rect 27338 15688 27344 15700
rect 26108 15660 27344 15688
rect 26108 15648 26114 15660
rect 27338 15648 27344 15660
rect 27396 15688 27402 15700
rect 27433 15691 27491 15697
rect 27433 15688 27445 15691
rect 27396 15660 27445 15688
rect 27396 15648 27402 15660
rect 27433 15657 27445 15660
rect 27479 15657 27491 15691
rect 28534 15688 28540 15700
rect 27433 15651 27491 15657
rect 27540 15660 28540 15688
rect 27540 15629 27568 15660
rect 28534 15648 28540 15660
rect 28592 15648 28598 15700
rect 28810 15648 28816 15700
rect 28868 15688 28874 15700
rect 29825 15691 29883 15697
rect 29825 15688 29837 15691
rect 28868 15660 29837 15688
rect 28868 15648 28874 15660
rect 29825 15657 29837 15660
rect 29871 15657 29883 15691
rect 29825 15651 29883 15657
rect 31110 15648 31116 15700
rect 31168 15688 31174 15700
rect 32125 15691 32183 15697
rect 32125 15688 32137 15691
rect 31168 15660 32137 15688
rect 31168 15648 31174 15660
rect 32125 15657 32137 15660
rect 32171 15657 32183 15691
rect 32125 15651 32183 15657
rect 32950 15648 32956 15700
rect 33008 15688 33014 15700
rect 37458 15688 37464 15700
rect 33008 15660 37464 15688
rect 33008 15648 33014 15660
rect 37458 15648 37464 15660
rect 37516 15648 37522 15700
rect 38102 15648 38108 15700
rect 38160 15648 38166 15700
rect 38654 15648 38660 15700
rect 38712 15648 38718 15700
rect 39301 15691 39359 15697
rect 39301 15657 39313 15691
rect 39347 15688 39359 15691
rect 39390 15688 39396 15700
rect 39347 15660 39396 15688
rect 39347 15657 39359 15660
rect 39301 15651 39359 15657
rect 39390 15648 39396 15660
rect 39448 15648 39454 15700
rect 42886 15648 42892 15700
rect 42944 15648 42950 15700
rect 44910 15688 44916 15700
rect 42996 15660 44916 15688
rect 27525 15623 27583 15629
rect 27525 15589 27537 15623
rect 27571 15589 27583 15623
rect 29362 15620 29368 15632
rect 27525 15583 27583 15589
rect 28552 15592 29368 15620
rect 26234 15512 26240 15564
rect 26292 15552 26298 15564
rect 27246 15552 27252 15564
rect 26292 15524 27252 15552
rect 26292 15512 26298 15524
rect 27246 15512 27252 15524
rect 27304 15552 27310 15564
rect 28552 15552 28580 15592
rect 29362 15580 29368 15592
rect 29420 15620 29426 15632
rect 30190 15620 30196 15632
rect 29420 15592 30196 15620
rect 29420 15580 29426 15592
rect 30190 15580 30196 15592
rect 30248 15580 30254 15632
rect 27304 15524 28580 15552
rect 27304 15512 27310 15524
rect 28626 15512 28632 15564
rect 28684 15512 28690 15564
rect 28718 15512 28724 15564
rect 28776 15512 28782 15564
rect 29638 15552 29644 15564
rect 28828 15524 29644 15552
rect 25130 15444 25136 15496
rect 25188 15444 25194 15496
rect 26050 15444 26056 15496
rect 26108 15444 26114 15496
rect 26789 15487 26847 15493
rect 26789 15453 26801 15487
rect 26835 15484 26847 15487
rect 26878 15484 26884 15496
rect 26835 15456 26884 15484
rect 26835 15453 26847 15456
rect 26789 15447 26847 15453
rect 26878 15444 26884 15456
rect 26936 15444 26942 15496
rect 27433 15487 27491 15493
rect 27433 15453 27445 15487
rect 27479 15484 27491 15487
rect 27614 15484 27620 15496
rect 27479 15456 27620 15484
rect 27479 15453 27491 15456
rect 27433 15447 27491 15453
rect 27614 15444 27620 15456
rect 27672 15444 27678 15496
rect 27893 15487 27951 15493
rect 27893 15453 27905 15487
rect 27939 15484 27951 15487
rect 28074 15484 28080 15496
rect 27939 15456 28080 15484
rect 27939 15453 27951 15456
rect 27893 15447 27951 15453
rect 28074 15444 28080 15456
rect 28132 15484 28138 15496
rect 28736 15484 28764 15512
rect 28132 15456 28764 15484
rect 28132 15444 28138 15456
rect 26970 15376 26976 15428
rect 27028 15416 27034 15428
rect 27709 15419 27767 15425
rect 27709 15416 27721 15419
rect 27028 15388 27721 15416
rect 27028 15376 27034 15388
rect 27709 15385 27721 15388
rect 27755 15416 27767 15419
rect 28828 15416 28856 15524
rect 29638 15512 29644 15524
rect 29696 15512 29702 15564
rect 29086 15444 29092 15496
rect 29144 15484 29150 15496
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29144 15456 29745 15484
rect 29144 15444 29150 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 29825 15487 29883 15493
rect 29825 15453 29837 15487
rect 29871 15453 29883 15487
rect 29825 15447 29883 15453
rect 30009 15487 30067 15493
rect 30009 15453 30021 15487
rect 30055 15484 30067 15487
rect 30098 15484 30104 15496
rect 30055 15456 30104 15484
rect 30055 15453 30067 15456
rect 30009 15447 30067 15453
rect 27755 15388 28856 15416
rect 29181 15419 29239 15425
rect 27755 15385 27767 15388
rect 27709 15379 27767 15385
rect 29181 15385 29193 15419
rect 29227 15416 29239 15419
rect 29840 15416 29868 15447
rect 30098 15444 30104 15456
rect 30156 15444 30162 15496
rect 30742 15444 30748 15496
rect 30800 15444 30806 15496
rect 32306 15444 32312 15496
rect 32364 15484 32370 15496
rect 32585 15487 32643 15493
rect 32585 15484 32597 15487
rect 32364 15456 32597 15484
rect 32364 15444 32370 15456
rect 32585 15453 32597 15456
rect 32631 15484 32643 15487
rect 34701 15487 34759 15493
rect 34701 15484 34713 15487
rect 32631 15456 34713 15484
rect 32631 15453 32643 15456
rect 32585 15447 32643 15453
rect 34701 15453 34713 15456
rect 34747 15484 34759 15487
rect 35342 15484 35348 15496
rect 34747 15456 35348 15484
rect 34747 15453 34759 15456
rect 34701 15447 34759 15453
rect 35342 15444 35348 15456
rect 35400 15484 35406 15496
rect 37274 15484 37280 15496
rect 35400 15456 37280 15484
rect 35400 15444 35406 15456
rect 37274 15444 37280 15456
rect 37332 15444 37338 15496
rect 37476 15493 37504 15648
rect 38672 15620 38700 15648
rect 40126 15620 40132 15632
rect 38672 15592 40132 15620
rect 40126 15580 40132 15592
rect 40184 15580 40190 15632
rect 42061 15623 42119 15629
rect 42061 15589 42073 15623
rect 42107 15620 42119 15623
rect 42996 15620 43024 15660
rect 44910 15648 44916 15660
rect 44968 15648 44974 15700
rect 45370 15648 45376 15700
rect 45428 15688 45434 15700
rect 45741 15691 45799 15697
rect 45741 15688 45753 15691
rect 45428 15660 45753 15688
rect 45428 15648 45434 15660
rect 45741 15657 45753 15660
rect 45787 15657 45799 15691
rect 45741 15651 45799 15657
rect 46290 15648 46296 15700
rect 46348 15648 46354 15700
rect 46750 15648 46756 15700
rect 46808 15688 46814 15700
rect 48222 15688 48228 15700
rect 46808 15660 48228 15688
rect 46808 15648 46814 15660
rect 48222 15648 48228 15660
rect 48280 15648 48286 15700
rect 50430 15648 50436 15700
rect 50488 15688 50494 15700
rect 51353 15691 51411 15697
rect 51353 15688 51365 15691
rect 50488 15660 51365 15688
rect 50488 15648 50494 15660
rect 51353 15657 51365 15660
rect 51399 15657 51411 15691
rect 51994 15688 52000 15700
rect 51353 15651 51411 15657
rect 51644 15660 52000 15688
rect 42107 15592 42288 15620
rect 42107 15589 42119 15592
rect 42061 15583 42119 15589
rect 39298 15552 39304 15564
rect 38856 15524 39304 15552
rect 38856 15496 38884 15524
rect 39298 15512 39304 15524
rect 39356 15512 39362 15564
rect 39942 15512 39948 15564
rect 40000 15552 40006 15564
rect 42260 15561 42288 15592
rect 42720 15592 43024 15620
rect 40681 15555 40739 15561
rect 40681 15552 40693 15555
rect 40000 15524 40693 15552
rect 40000 15512 40006 15524
rect 40681 15521 40693 15524
rect 40727 15521 40739 15555
rect 40681 15515 40739 15521
rect 42245 15555 42303 15561
rect 42245 15521 42257 15555
rect 42291 15521 42303 15555
rect 42245 15515 42303 15521
rect 37461 15487 37519 15493
rect 37461 15453 37473 15487
rect 37507 15453 37519 15487
rect 38010 15484 38016 15496
rect 37461 15447 37519 15453
rect 37752 15456 38016 15484
rect 29227 15388 29868 15416
rect 31012 15419 31070 15425
rect 29227 15385 29239 15388
rect 29181 15379 29239 15385
rect 31012 15385 31024 15419
rect 31058 15416 31070 15419
rect 31662 15416 31668 15428
rect 31058 15388 31668 15416
rect 31058 15385 31070 15388
rect 31012 15379 31070 15385
rect 31662 15376 31668 15388
rect 31720 15376 31726 15428
rect 32852 15419 32910 15425
rect 32852 15385 32864 15419
rect 32898 15416 32910 15419
rect 33134 15416 33140 15428
rect 32898 15388 33140 15416
rect 32898 15385 32910 15388
rect 32852 15379 32910 15385
rect 33134 15376 33140 15388
rect 33192 15376 33198 15428
rect 33888 15388 34744 15416
rect 25685 15351 25743 15357
rect 25685 15317 25697 15351
rect 25731 15348 25743 15351
rect 26234 15348 26240 15360
rect 25731 15320 26240 15348
rect 25731 15317 25743 15320
rect 25685 15311 25743 15317
rect 26234 15308 26240 15320
rect 26292 15308 26298 15360
rect 26602 15308 26608 15360
rect 26660 15308 26666 15360
rect 27062 15308 27068 15360
rect 27120 15348 27126 15360
rect 27341 15351 27399 15357
rect 27341 15348 27353 15351
rect 27120 15320 27353 15348
rect 27120 15308 27126 15320
rect 27341 15317 27353 15320
rect 27387 15317 27399 15351
rect 27341 15311 27399 15317
rect 28445 15351 28503 15357
rect 28445 15317 28457 15351
rect 28491 15348 28503 15351
rect 28718 15348 28724 15360
rect 28491 15320 28724 15348
rect 28491 15317 28503 15320
rect 28445 15311 28503 15317
rect 28718 15308 28724 15320
rect 28776 15308 28782 15360
rect 29546 15308 29552 15360
rect 29604 15308 29610 15360
rect 30650 15308 30656 15360
rect 30708 15348 30714 15360
rect 33888 15348 33916 15388
rect 34716 15360 34744 15388
rect 34790 15376 34796 15428
rect 34848 15416 34854 15428
rect 34946 15419 35004 15425
rect 34946 15416 34958 15419
rect 34848 15388 34958 15416
rect 34848 15376 34854 15388
rect 34946 15385 34958 15388
rect 34992 15385 35004 15419
rect 34946 15379 35004 15385
rect 37550 15376 37556 15428
rect 37608 15416 37614 15428
rect 37752 15425 37780 15456
rect 38010 15444 38016 15456
rect 38068 15444 38074 15496
rect 38838 15444 38844 15496
rect 38896 15444 38902 15496
rect 39022 15444 39028 15496
rect 39080 15484 39086 15496
rect 39485 15487 39543 15493
rect 39485 15484 39497 15487
rect 39080 15456 39497 15484
rect 39080 15444 39086 15456
rect 39485 15453 39497 15456
rect 39531 15453 39543 15487
rect 39485 15447 39543 15453
rect 40218 15444 40224 15496
rect 40276 15484 40282 15496
rect 40313 15487 40371 15493
rect 40313 15484 40325 15487
rect 40276 15456 40325 15484
rect 40276 15444 40282 15456
rect 40313 15453 40325 15456
rect 40359 15453 40371 15487
rect 40313 15447 40371 15453
rect 40402 15444 40408 15496
rect 40460 15444 40466 15496
rect 40497 15487 40555 15493
rect 40497 15453 40509 15487
rect 40543 15484 40555 15487
rect 42720 15484 42748 15592
rect 42794 15512 42800 15564
rect 42852 15552 42858 15564
rect 42981 15555 43039 15561
rect 42981 15552 42993 15555
rect 42852 15524 42993 15552
rect 42852 15512 42858 15524
rect 42981 15521 42993 15524
rect 43027 15521 43039 15555
rect 42981 15515 43039 15521
rect 43349 15555 43407 15561
rect 43349 15521 43361 15555
rect 43395 15552 43407 15555
rect 43622 15552 43628 15564
rect 43395 15524 43628 15552
rect 43395 15521 43407 15524
rect 43349 15515 43407 15521
rect 43622 15512 43628 15524
rect 43680 15512 43686 15564
rect 44726 15512 44732 15564
rect 44784 15561 44790 15564
rect 44784 15555 44833 15561
rect 44784 15521 44787 15555
rect 44821 15552 44833 15555
rect 45097 15555 45155 15561
rect 45097 15552 45109 15555
rect 44821 15524 45109 15552
rect 44821 15521 44833 15524
rect 44784 15515 44833 15521
rect 45097 15521 45109 15524
rect 45143 15521 45155 15555
rect 45097 15515 45155 15521
rect 46109 15555 46167 15561
rect 46109 15521 46121 15555
rect 46155 15552 46167 15555
rect 46308 15552 46336 15648
rect 46768 15561 46796 15648
rect 46155 15524 46336 15552
rect 46753 15555 46811 15561
rect 46155 15521 46167 15524
rect 46109 15515 46167 15521
rect 46753 15521 46765 15555
rect 46799 15521 46811 15555
rect 46753 15515 46811 15521
rect 44784 15512 44790 15515
rect 51644 15503 51672 15660
rect 51994 15648 52000 15660
rect 52052 15648 52058 15700
rect 52362 15648 52368 15700
rect 52420 15648 52426 15700
rect 52089 15555 52147 15561
rect 52089 15521 52101 15555
rect 52135 15552 52147 15555
rect 52380 15552 52408 15648
rect 52546 15580 52552 15632
rect 52604 15620 52610 15632
rect 52604 15592 53420 15620
rect 52604 15580 52610 15592
rect 52135 15524 52408 15552
rect 52135 15521 52147 15524
rect 52089 15515 52147 15521
rect 51638 15497 51696 15503
rect 40543 15456 42748 15484
rect 40543 15453 40555 15456
rect 40497 15447 40555 15453
rect 44634 15444 44640 15496
rect 44692 15484 44698 15496
rect 47394 15484 47400 15496
rect 44692 15456 47400 15484
rect 44692 15444 44698 15456
rect 47394 15444 47400 15456
rect 47452 15444 47458 15496
rect 48225 15487 48283 15493
rect 48225 15484 48237 15487
rect 48148 15456 48237 15484
rect 37737 15419 37795 15425
rect 37737 15416 37749 15419
rect 37608 15388 37749 15416
rect 37608 15376 37614 15388
rect 37737 15385 37749 15388
rect 37783 15385 37795 15419
rect 37737 15379 37795 15385
rect 39206 15376 39212 15428
rect 39264 15376 39270 15428
rect 40129 15419 40187 15425
rect 40129 15385 40141 15419
rect 40175 15416 40187 15419
rect 40926 15419 40984 15425
rect 40926 15416 40938 15419
rect 40175 15388 40938 15416
rect 40175 15385 40187 15388
rect 40129 15379 40187 15385
rect 40926 15385 40938 15388
rect 40972 15385 40984 15419
rect 40926 15379 40984 15385
rect 44358 15376 44364 15428
rect 44416 15376 44422 15428
rect 46661 15419 46719 15425
rect 46661 15385 46673 15419
rect 46707 15416 46719 15419
rect 46998 15419 47056 15425
rect 46998 15416 47010 15419
rect 46707 15388 47010 15416
rect 46707 15385 46719 15388
rect 46661 15379 46719 15385
rect 46998 15385 47010 15388
rect 47044 15385 47056 15419
rect 46998 15379 47056 15385
rect 30708 15320 33916 15348
rect 30708 15308 30714 15320
rect 33962 15308 33968 15360
rect 34020 15308 34026 15360
rect 34698 15308 34704 15360
rect 34756 15348 34762 15360
rect 36078 15348 36084 15360
rect 34756 15320 36084 15348
rect 34756 15308 34762 15320
rect 36078 15308 36084 15320
rect 36136 15308 36142 15360
rect 44174 15308 44180 15360
rect 44232 15348 44238 15360
rect 45830 15348 45836 15360
rect 44232 15320 45836 15348
rect 44232 15308 44238 15320
rect 45830 15308 45836 15320
rect 45888 15308 45894 15360
rect 48148 15357 48176 15456
rect 48225 15453 48237 15456
rect 48271 15453 48283 15487
rect 48225 15447 48283 15453
rect 49786 15444 49792 15496
rect 49844 15444 49850 15496
rect 50801 15487 50859 15493
rect 50801 15453 50813 15487
rect 50847 15484 50859 15487
rect 51445 15487 51503 15493
rect 51445 15484 51457 15487
rect 50847 15456 51457 15484
rect 50847 15453 50859 15456
rect 50801 15447 50859 15453
rect 51445 15453 51457 15456
rect 51491 15453 51503 15487
rect 51638 15463 51650 15497
rect 51684 15463 51696 15497
rect 51638 15457 51696 15463
rect 51445 15447 51503 15453
rect 51810 15444 51816 15496
rect 51868 15444 51874 15496
rect 51951 15487 52009 15493
rect 51951 15453 51963 15487
rect 51997 15484 52009 15487
rect 52549 15487 52607 15493
rect 52549 15484 52561 15487
rect 51997 15456 52561 15484
rect 51997 15453 52009 15456
rect 51951 15447 52009 15453
rect 52104 15428 52132 15456
rect 52549 15453 52561 15456
rect 52595 15453 52607 15487
rect 52549 15447 52607 15453
rect 52638 15444 52644 15496
rect 52696 15444 52702 15496
rect 53392 15493 53420 15592
rect 52825 15487 52883 15493
rect 52825 15453 52837 15487
rect 52871 15453 52883 15487
rect 52825 15447 52883 15453
rect 53377 15487 53435 15493
rect 53377 15453 53389 15487
rect 53423 15484 53435 15487
rect 54478 15484 54484 15496
rect 53423 15456 54484 15484
rect 53423 15453 53435 15456
rect 53377 15447 53435 15453
rect 51626 15376 51632 15428
rect 51684 15416 51690 15428
rect 51722 15419 51780 15425
rect 51722 15416 51734 15419
rect 51684 15388 51734 15416
rect 51684 15376 51690 15388
rect 51722 15385 51734 15388
rect 51768 15385 51780 15419
rect 51722 15379 51780 15385
rect 52086 15376 52092 15428
rect 52144 15376 52150 15428
rect 52178 15376 52184 15428
rect 52236 15376 52242 15428
rect 52365 15419 52423 15425
rect 52365 15385 52377 15419
rect 52411 15416 52423 15419
rect 52733 15419 52791 15425
rect 52733 15416 52745 15419
rect 52411 15388 52745 15416
rect 52411 15385 52423 15388
rect 52365 15379 52423 15385
rect 52733 15385 52745 15388
rect 52779 15385 52791 15419
rect 52733 15379 52791 15385
rect 48133 15351 48191 15357
rect 48133 15317 48145 15351
rect 48179 15317 48191 15351
rect 48133 15311 48191 15317
rect 48317 15351 48375 15357
rect 48317 15317 48329 15351
rect 48363 15348 48375 15351
rect 48498 15348 48504 15360
rect 48363 15320 48504 15348
rect 48363 15317 48375 15320
rect 48317 15311 48375 15317
rect 48498 15308 48504 15320
rect 48556 15308 48562 15360
rect 49878 15308 49884 15360
rect 49936 15308 49942 15360
rect 51994 15308 52000 15360
rect 52052 15348 52058 15360
rect 52380 15348 52408 15379
rect 52052 15320 52408 15348
rect 52052 15308 52058 15320
rect 52454 15308 52460 15360
rect 52512 15348 52518 15360
rect 52840 15348 52868 15447
rect 54478 15444 54484 15456
rect 54536 15444 54542 15496
rect 52512 15320 52868 15348
rect 52512 15308 52518 15320
rect 53926 15308 53932 15360
rect 53984 15308 53990 15360
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 26050 15104 26056 15156
rect 26108 15144 26114 15156
rect 26605 15147 26663 15153
rect 26605 15144 26617 15147
rect 26108 15116 26617 15144
rect 26108 15104 26114 15116
rect 26605 15113 26617 15116
rect 26651 15113 26663 15147
rect 26605 15107 26663 15113
rect 27065 15147 27123 15153
rect 27065 15113 27077 15147
rect 27111 15113 27123 15147
rect 27065 15107 27123 15113
rect 25492 15079 25550 15085
rect 23768 15048 25176 15076
rect 23768 15017 23796 15048
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 14977 23811 15011
rect 23753 14971 23811 14977
rect 24020 15011 24078 15017
rect 24020 14977 24032 15011
rect 24066 15008 24078 15011
rect 24854 15008 24860 15020
rect 24066 14980 24860 15008
rect 24066 14977 24078 14980
rect 24020 14971 24078 14977
rect 24854 14968 24860 14980
rect 24912 14968 24918 15020
rect 25148 14940 25176 15048
rect 25492 15045 25504 15079
rect 25538 15076 25550 15079
rect 27080 15076 27108 15107
rect 27614 15104 27620 15156
rect 27672 15144 27678 15156
rect 28629 15147 28687 15153
rect 28629 15144 28641 15147
rect 27672 15116 28641 15144
rect 27672 15104 27678 15116
rect 28629 15113 28641 15116
rect 28675 15113 28687 15147
rect 28629 15107 28687 15113
rect 25538 15048 27108 15076
rect 25538 15045 25550 15048
rect 25492 15039 25550 15045
rect 26973 15011 27031 15017
rect 26973 14977 26985 15011
rect 27019 15008 27031 15011
rect 27062 15008 27068 15020
rect 27019 14980 27068 15008
rect 27019 14977 27031 14980
rect 26973 14971 27031 14977
rect 27062 14968 27068 14980
rect 27120 14968 27126 15020
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 15008 27215 15011
rect 27246 15008 27252 15020
rect 27203 14980 27252 15008
rect 27203 14977 27215 14980
rect 27157 14971 27215 14977
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 27338 14968 27344 15020
rect 27396 14968 27402 15020
rect 28074 14968 28080 15020
rect 28132 14968 28138 15020
rect 25222 14940 25228 14952
rect 25148 14912 25228 14940
rect 25222 14900 25228 14912
rect 25280 14900 25286 14952
rect 28644 14940 28672 15107
rect 28902 15104 28908 15156
rect 28960 15104 28966 15156
rect 29086 15104 29092 15156
rect 29144 15104 29150 15156
rect 30837 15147 30895 15153
rect 30837 15113 30849 15147
rect 30883 15144 30895 15147
rect 31202 15144 31208 15156
rect 30883 15116 31208 15144
rect 30883 15113 30895 15116
rect 30837 15107 30895 15113
rect 31202 15104 31208 15116
rect 31260 15104 31266 15156
rect 31662 15104 31668 15156
rect 31720 15104 31726 15156
rect 31846 15104 31852 15156
rect 31904 15104 31910 15156
rect 33689 15147 33747 15153
rect 33689 15113 33701 15147
rect 33735 15144 33747 15147
rect 33778 15144 33784 15156
rect 33735 15116 33784 15144
rect 33735 15113 33747 15116
rect 33689 15107 33747 15113
rect 33778 15104 33784 15116
rect 33836 15104 33842 15156
rect 34422 15104 34428 15156
rect 34480 15104 34486 15156
rect 38654 15144 38660 15156
rect 34532 15116 38660 15144
rect 28718 14968 28724 15020
rect 28776 14968 28782 15020
rect 28920 15017 28948 15104
rect 29546 15036 29552 15088
rect 29604 15076 29610 15088
rect 29702 15079 29760 15085
rect 29702 15076 29714 15079
rect 29604 15048 29714 15076
rect 29604 15036 29610 15048
rect 29702 15045 29714 15048
rect 29748 15045 29760 15079
rect 29702 15039 29760 15045
rect 28905 15011 28963 15017
rect 28905 14977 28917 15011
rect 28951 14977 28963 15011
rect 28905 14971 28963 14977
rect 29181 15011 29239 15017
rect 29181 14977 29193 15011
rect 29227 14977 29239 15011
rect 29181 14971 29239 14977
rect 29196 14940 29224 14971
rect 29454 14968 29460 15020
rect 29512 15008 29518 15020
rect 30742 15008 30748 15020
rect 29512 14980 30748 15008
rect 29512 14968 29518 14980
rect 30742 14968 30748 14980
rect 30800 14968 30806 15020
rect 31757 15011 31815 15017
rect 31757 14977 31769 15011
rect 31803 15008 31815 15011
rect 31864 15008 31892 15104
rect 34532 15076 34560 15116
rect 38654 15104 38660 15116
rect 38712 15104 38718 15156
rect 40402 15104 40408 15156
rect 40460 15144 40466 15156
rect 42429 15147 42487 15153
rect 40460 15116 41276 15144
rect 40460 15104 40466 15116
rect 34440 15048 34560 15076
rect 31803 14980 31892 15008
rect 32576 15011 32634 15017
rect 31803 14977 31815 14980
rect 31757 14971 31815 14977
rect 32576 14977 32588 15011
rect 32622 15008 32634 15011
rect 33134 15008 33140 15020
rect 32622 14980 33140 15008
rect 32622 14977 32634 14980
rect 32576 14971 32634 14977
rect 33134 14968 33140 14980
rect 33192 14968 33198 15020
rect 33410 14968 33416 15020
rect 33468 14968 33474 15020
rect 34440 15017 34468 15048
rect 34698 15036 34704 15088
rect 34756 15076 34762 15088
rect 38473 15079 38531 15085
rect 34756 15048 35020 15076
rect 34756 15036 34762 15048
rect 34422 15011 34480 15017
rect 34422 14977 34434 15011
rect 34468 14977 34480 15011
rect 34422 14971 34480 14977
rect 34514 14968 34520 15020
rect 34572 15008 34578 15020
rect 34992 15017 35020 15048
rect 38473 15045 38485 15079
rect 38519 15076 38531 15079
rect 38838 15076 38844 15088
rect 38519 15048 38844 15076
rect 38519 15045 38531 15048
rect 38473 15039 38531 15045
rect 38838 15036 38844 15048
rect 38896 15036 38902 15088
rect 41248 15085 41276 15116
rect 42429 15113 42441 15147
rect 42475 15144 42487 15147
rect 42610 15144 42616 15156
rect 42475 15116 42616 15144
rect 42475 15113 42487 15116
rect 42429 15107 42487 15113
rect 42610 15104 42616 15116
rect 42668 15104 42674 15156
rect 44358 15104 44364 15156
rect 44416 15144 44422 15156
rect 44545 15147 44603 15153
rect 44545 15144 44557 15147
rect 44416 15116 44557 15144
rect 44416 15104 44422 15116
rect 44545 15113 44557 15116
rect 44591 15113 44603 15147
rect 44545 15107 44603 15113
rect 45186 15104 45192 15156
rect 45244 15144 45250 15156
rect 45373 15147 45431 15153
rect 45373 15144 45385 15147
rect 45244 15116 45385 15144
rect 45244 15104 45250 15116
rect 45373 15113 45385 15116
rect 45419 15113 45431 15147
rect 45373 15107 45431 15113
rect 48958 15104 48964 15156
rect 49016 15104 49022 15156
rect 51718 15144 51724 15156
rect 51276 15116 51724 15144
rect 41233 15079 41291 15085
rect 40144 15048 40632 15076
rect 34885 15011 34943 15017
rect 34885 15008 34897 15011
rect 34572 14980 34897 15008
rect 34572 14968 34578 14980
rect 34885 14977 34897 14980
rect 34931 14977 34943 15011
rect 34885 14971 34943 14977
rect 34977 15011 35035 15017
rect 34977 14977 34989 15011
rect 35023 14977 35035 15011
rect 34977 14971 35035 14977
rect 35342 14968 35348 15020
rect 35400 15017 35406 15020
rect 35400 15008 35410 15017
rect 35612 15011 35670 15017
rect 35400 14980 35445 15008
rect 35400 14971 35410 14980
rect 35612 14977 35624 15011
rect 35658 15008 35670 15011
rect 36446 15008 36452 15020
rect 35658 14980 36452 15008
rect 35658 14977 35670 14980
rect 35612 14971 35670 14977
rect 35400 14968 35406 14971
rect 36446 14968 36452 14980
rect 36504 14968 36510 15020
rect 36817 15011 36875 15017
rect 36817 14977 36829 15011
rect 36863 14977 36875 15011
rect 36817 14971 36875 14977
rect 37001 15011 37059 15017
rect 37001 14977 37013 15011
rect 37047 14977 37059 15011
rect 37001 14971 37059 14977
rect 28644 14912 29224 14940
rect 31018 14900 31024 14952
rect 31076 14900 31082 14952
rect 32306 14900 32312 14952
rect 32364 14900 32370 14952
rect 33428 14940 33456 14968
rect 34238 14940 34244 14952
rect 33428 14912 34244 14940
rect 34238 14900 34244 14912
rect 34296 14940 34302 14952
rect 34793 14943 34851 14949
rect 34793 14940 34805 14943
rect 34296 14912 34805 14940
rect 34296 14900 34302 14912
rect 34793 14909 34805 14912
rect 34839 14909 34851 14943
rect 36832 14940 36860 14971
rect 34793 14903 34851 14909
rect 36372 14912 36860 14940
rect 36372 14816 36400 14912
rect 37016 14872 37044 14971
rect 36556 14844 37044 14872
rect 38856 14872 38884 15036
rect 39482 14968 39488 15020
rect 39540 14968 39546 15020
rect 39945 15011 40003 15017
rect 39945 15008 39957 15011
rect 39592 14980 39957 15008
rect 39206 14900 39212 14952
rect 39264 14940 39270 14952
rect 39592 14940 39620 14980
rect 39945 14977 39957 14980
rect 39991 14977 40003 15011
rect 39945 14971 40003 14977
rect 39264 14912 39620 14940
rect 39761 14943 39819 14949
rect 39264 14900 39270 14912
rect 39761 14909 39773 14943
rect 39807 14909 39819 14943
rect 39761 14903 39819 14909
rect 39776 14872 39804 14903
rect 38856 14844 39804 14872
rect 36556 14816 36584 14844
rect 40144 14816 40172 15048
rect 40221 15011 40279 15017
rect 40221 14977 40233 15011
rect 40267 14977 40279 15011
rect 40221 14971 40279 14977
rect 40236 14940 40264 14971
rect 40402 14968 40408 15020
rect 40460 14968 40466 15020
rect 40494 14968 40500 15020
rect 40552 14968 40558 15020
rect 40604 15017 40632 15048
rect 41233 15045 41245 15079
rect 41279 15076 41291 15079
rect 43806 15076 43812 15088
rect 41279 15048 41414 15076
rect 41279 15045 41291 15048
rect 41233 15039 41291 15045
rect 40589 15011 40647 15017
rect 40589 14977 40601 15011
rect 40635 14977 40647 15011
rect 40589 14971 40647 14977
rect 40770 14968 40776 15020
rect 40828 15008 40834 15020
rect 40957 15011 41015 15017
rect 40957 15008 40969 15011
rect 40828 14980 40969 15008
rect 40828 14968 40834 14980
rect 40957 14977 40969 14980
rect 41003 14977 41015 15011
rect 40957 14971 41015 14977
rect 40236 14912 40724 14940
rect 40696 14816 40724 14912
rect 41386 14872 41414 15048
rect 42628 15048 43812 15076
rect 42628 15017 42656 15048
rect 43806 15036 43812 15048
rect 43864 15036 43870 15088
rect 48774 15076 48780 15088
rect 45940 15048 46796 15076
rect 42613 15011 42671 15017
rect 42613 14977 42625 15011
rect 42659 14977 42671 15011
rect 42613 14971 42671 14977
rect 42705 15011 42763 15017
rect 42705 14977 42717 15011
rect 42751 15008 42763 15011
rect 42794 15008 42800 15020
rect 42751 14980 42800 15008
rect 42751 14977 42763 14980
rect 42705 14971 42763 14977
rect 42794 14968 42800 14980
rect 42852 14968 42858 15020
rect 42886 14968 42892 15020
rect 42944 14968 42950 15020
rect 42981 15011 43039 15017
rect 42981 14977 42993 15011
rect 43027 14977 43039 15011
rect 42981 14971 43039 14977
rect 44453 15011 44511 15017
rect 44453 14977 44465 15011
rect 44499 14977 44511 15011
rect 44453 14971 44511 14977
rect 42242 14900 42248 14952
rect 42300 14940 42306 14952
rect 42996 14940 43024 14971
rect 42300 14912 43024 14940
rect 42300 14900 42306 14912
rect 43806 14900 43812 14952
rect 43864 14900 43870 14952
rect 44082 14900 44088 14952
rect 44140 14900 44146 14952
rect 44266 14900 44272 14952
rect 44324 14940 44330 14952
rect 44361 14943 44419 14949
rect 44361 14940 44373 14943
rect 44324 14912 44373 14940
rect 44324 14900 44330 14912
rect 44361 14909 44373 14912
rect 44407 14909 44419 14943
rect 44361 14903 44419 14909
rect 44100 14872 44128 14900
rect 41386 14844 44128 14872
rect 25130 14764 25136 14816
rect 25188 14764 25194 14816
rect 27890 14764 27896 14816
rect 27948 14764 27954 14816
rect 29270 14764 29276 14816
rect 29328 14764 29334 14816
rect 31849 14807 31907 14813
rect 31849 14773 31861 14807
rect 31895 14804 31907 14807
rect 33594 14804 33600 14816
rect 31895 14776 33600 14804
rect 31895 14773 31907 14776
rect 31849 14767 31907 14773
rect 33594 14764 33600 14776
rect 33652 14764 33658 14816
rect 33686 14764 33692 14816
rect 33744 14804 33750 14816
rect 34241 14807 34299 14813
rect 34241 14804 34253 14807
rect 33744 14776 34253 14804
rect 33744 14764 33750 14776
rect 34241 14773 34253 14776
rect 34287 14773 34299 14807
rect 34241 14767 34299 14773
rect 35069 14807 35127 14813
rect 35069 14773 35081 14807
rect 35115 14804 35127 14807
rect 35250 14804 35256 14816
rect 35115 14776 35256 14804
rect 35115 14773 35127 14776
rect 35069 14767 35127 14773
rect 35250 14764 35256 14776
rect 35308 14764 35314 14816
rect 36354 14764 36360 14816
rect 36412 14764 36418 14816
rect 36538 14764 36544 14816
rect 36596 14764 36602 14816
rect 36722 14764 36728 14816
rect 36780 14764 36786 14816
rect 36814 14764 36820 14816
rect 36872 14764 36878 14816
rect 38749 14807 38807 14813
rect 38749 14773 38761 14807
rect 38795 14804 38807 14807
rect 38930 14804 38936 14816
rect 38795 14776 38936 14804
rect 38795 14773 38807 14776
rect 38749 14767 38807 14773
rect 38930 14764 38936 14776
rect 38988 14764 38994 14816
rect 39574 14764 39580 14816
rect 39632 14764 39638 14816
rect 40126 14764 40132 14816
rect 40184 14764 40190 14816
rect 40678 14764 40684 14816
rect 40736 14764 40742 14816
rect 40773 14807 40831 14813
rect 40773 14773 40785 14807
rect 40819 14804 40831 14807
rect 40954 14804 40960 14816
rect 40819 14776 40960 14804
rect 40819 14773 40831 14776
rect 40773 14767 40831 14773
rect 40954 14764 40960 14776
rect 41012 14764 41018 14816
rect 44174 14764 44180 14816
rect 44232 14804 44238 14816
rect 44476 14804 44504 14971
rect 44726 14968 44732 15020
rect 44784 15008 44790 15020
rect 45005 15011 45063 15017
rect 45005 15008 45017 15011
rect 44784 14980 45017 15008
rect 44784 14968 44790 14980
rect 45005 14977 45017 14980
rect 45051 14977 45063 15011
rect 45005 14971 45063 14977
rect 45189 15011 45247 15017
rect 45189 14977 45201 15011
rect 45235 15008 45247 15011
rect 45646 15008 45652 15020
rect 45235 14980 45652 15008
rect 45235 14977 45247 14980
rect 45189 14971 45247 14977
rect 45646 14968 45652 14980
rect 45704 14968 45710 15020
rect 45940 15017 45968 15048
rect 46768 15020 46796 15048
rect 48424 15048 48780 15076
rect 45925 15011 45983 15017
rect 45925 14977 45937 15011
rect 45971 14977 45983 15011
rect 45925 14971 45983 14977
rect 46192 15011 46250 15017
rect 46192 14977 46204 15011
rect 46238 15008 46250 15011
rect 46566 15008 46572 15020
rect 46238 14980 46572 15008
rect 46238 14977 46250 14980
rect 46192 14971 46250 14977
rect 46566 14968 46572 14980
rect 46624 14968 46630 15020
rect 46750 14968 46756 15020
rect 46808 14968 46814 15020
rect 48424 15017 48452 15048
rect 48774 15036 48780 15048
rect 48832 15036 48838 15088
rect 48976 15076 49004 15104
rect 51276 15088 51304 15116
rect 51718 15104 51724 15116
rect 51776 15104 51782 15156
rect 53926 15144 53932 15156
rect 52012 15116 53932 15144
rect 48884 15048 49004 15076
rect 48884 15017 48912 15048
rect 49878 15036 49884 15088
rect 49936 15036 49942 15088
rect 51258 15036 51264 15088
rect 51316 15036 51322 15088
rect 51626 15076 51632 15088
rect 51476 15048 51632 15076
rect 51476 15045 51549 15048
rect 48409 15011 48467 15017
rect 48409 14977 48421 15011
rect 48455 14977 48467 15011
rect 48409 14971 48467 14977
rect 48501 15011 48559 15017
rect 48501 14977 48513 15011
rect 48547 15008 48559 15011
rect 48869 15011 48927 15017
rect 48547 14980 48636 15008
rect 48547 14977 48559 14980
rect 48501 14971 48559 14977
rect 48608 14952 48636 14980
rect 48869 14977 48881 15011
rect 48915 14977 48927 15011
rect 51476 15011 51503 15045
rect 51537 15011 51549 15045
rect 51626 15036 51632 15048
rect 51684 15036 51690 15088
rect 52012 15017 52040 15116
rect 53926 15104 53932 15116
rect 53984 15104 53990 15156
rect 54478 15104 54484 15156
rect 54536 15104 54542 15156
rect 52270 15036 52276 15088
rect 52328 15076 52334 15088
rect 52328 15048 52776 15076
rect 52328 15036 52334 15048
rect 51476 15008 51549 15011
rect 51721 15011 51779 15017
rect 51721 15008 51733 15011
rect 48869 14971 48927 14977
rect 51460 15005 51549 15008
rect 51460 14980 51504 15005
rect 51644 14980 51733 15008
rect 51460 14952 51488 14980
rect 47578 14940 47584 14952
rect 47320 14912 47584 14940
rect 47320 14881 47348 14912
rect 47578 14900 47584 14912
rect 47636 14900 47642 14952
rect 48590 14900 48596 14952
rect 48648 14900 48654 14952
rect 48682 14900 48688 14952
rect 48740 14900 48746 14952
rect 49142 14900 49148 14952
rect 49200 14900 49206 14952
rect 51442 14900 51448 14952
rect 51500 14900 51506 14952
rect 51644 14881 51672 14980
rect 51721 14977 51733 14980
rect 51767 14977 51779 15011
rect 51721 14971 51779 14977
rect 51905 15011 51963 15017
rect 51905 14977 51917 15011
rect 51951 14977 51963 15011
rect 51905 14971 51963 14977
rect 51997 15011 52055 15017
rect 51997 14977 52009 15011
rect 52043 14977 52055 15011
rect 51997 14971 52055 14977
rect 51920 14940 51948 14971
rect 52086 14968 52092 15020
rect 52144 14968 52150 15020
rect 52365 15011 52423 15017
rect 52365 14977 52377 15011
rect 52411 15008 52423 15011
rect 52454 15008 52460 15020
rect 52411 14980 52460 15008
rect 52411 14977 52423 14980
rect 52365 14971 52423 14977
rect 52454 14968 52460 14980
rect 52512 14968 52518 15020
rect 52546 14968 52552 15020
rect 52604 14968 52610 15020
rect 52748 15017 52776 15048
rect 53466 15036 53472 15088
rect 53524 15036 53530 15088
rect 52733 15011 52791 15017
rect 52733 14977 52745 15011
rect 52779 14977 52791 15011
rect 52733 14971 52791 14977
rect 53009 14943 53067 14949
rect 53009 14940 53021 14943
rect 51920 14912 52224 14940
rect 47305 14875 47363 14881
rect 47305 14841 47317 14875
rect 47351 14841 47363 14875
rect 51629 14875 51687 14881
rect 47305 14835 47363 14841
rect 47412 14844 49004 14872
rect 47412 14804 47440 14844
rect 44232 14776 47440 14804
rect 44232 14764 44238 14776
rect 47486 14764 47492 14816
rect 47544 14804 47550 14816
rect 48225 14807 48283 14813
rect 48225 14804 48237 14807
rect 47544 14776 48237 14804
rect 47544 14764 47550 14776
rect 48225 14773 48237 14776
rect 48271 14773 48283 14807
rect 48225 14767 48283 14773
rect 48314 14764 48320 14816
rect 48372 14804 48378 14816
rect 48682 14804 48688 14816
rect 48372 14776 48688 14804
rect 48372 14764 48378 14776
rect 48682 14764 48688 14776
rect 48740 14764 48746 14816
rect 48976 14804 49004 14844
rect 51629 14841 51641 14875
rect 51675 14841 51687 14875
rect 51629 14835 51687 14841
rect 49786 14804 49792 14816
rect 48976 14776 49792 14804
rect 49786 14764 49792 14776
rect 49844 14764 49850 14816
rect 50617 14807 50675 14813
rect 50617 14773 50629 14807
rect 50663 14804 50675 14807
rect 50706 14804 50712 14816
rect 50663 14776 50712 14804
rect 50663 14773 50675 14776
rect 50617 14767 50675 14773
rect 50706 14764 50712 14776
rect 50764 14804 50770 14816
rect 51445 14807 51503 14813
rect 51445 14804 51457 14807
rect 50764 14776 51457 14804
rect 50764 14764 50770 14776
rect 51445 14773 51457 14776
rect 51491 14804 51503 14807
rect 51534 14804 51540 14816
rect 51491 14776 51540 14804
rect 51491 14773 51503 14776
rect 51445 14767 51503 14773
rect 51534 14764 51540 14776
rect 51592 14764 51598 14816
rect 51644 14804 51672 14835
rect 51994 14804 52000 14816
rect 51644 14776 52000 14804
rect 51994 14764 52000 14776
rect 52052 14764 52058 14816
rect 52196 14804 52224 14912
rect 52748 14912 53021 14940
rect 52273 14875 52331 14881
rect 52273 14841 52285 14875
rect 52319 14872 52331 14875
rect 52748 14872 52776 14912
rect 53009 14909 53021 14912
rect 53055 14909 53067 14943
rect 53009 14903 53067 14909
rect 52319 14844 52776 14872
rect 52319 14841 52331 14844
rect 52273 14835 52331 14841
rect 52365 14807 52423 14813
rect 52365 14804 52377 14807
rect 52196 14776 52377 14804
rect 52365 14773 52377 14776
rect 52411 14773 52423 14807
rect 52365 14767 52423 14773
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 26326 14560 26332 14612
rect 26384 14560 26390 14612
rect 26878 14560 26884 14612
rect 26936 14560 26942 14612
rect 29270 14560 29276 14612
rect 29328 14560 29334 14612
rect 31018 14560 31024 14612
rect 31076 14560 31082 14612
rect 31846 14600 31852 14612
rect 31726 14572 31852 14600
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 25961 14467 26019 14473
rect 25961 14464 25973 14467
rect 24912 14436 25973 14464
rect 24912 14424 24918 14436
rect 25961 14433 25973 14436
rect 26007 14433 26019 14467
rect 25961 14427 26019 14433
rect 26050 14424 26056 14476
rect 26108 14424 26114 14476
rect 27249 14467 27307 14473
rect 27249 14464 27261 14467
rect 27080 14436 27261 14464
rect 25130 14356 25136 14408
rect 25188 14396 25194 14408
rect 25777 14399 25835 14405
rect 25777 14396 25789 14399
rect 25188 14368 25789 14396
rect 25188 14356 25194 14368
rect 25777 14365 25789 14368
rect 25823 14365 25835 14399
rect 25777 14359 25835 14365
rect 25869 14399 25927 14405
rect 25869 14365 25881 14399
rect 25915 14396 25927 14399
rect 26068 14396 26096 14424
rect 27080 14408 27108 14436
rect 27249 14433 27261 14436
rect 27295 14433 27307 14467
rect 29288 14464 29316 14560
rect 29914 14492 29920 14544
rect 29972 14492 29978 14544
rect 29288 14436 30052 14464
rect 27249 14427 27307 14433
rect 25915 14368 26096 14396
rect 25915 14365 25927 14368
rect 25869 14359 25927 14365
rect 26234 14356 26240 14408
rect 26292 14356 26298 14408
rect 26602 14356 26608 14408
rect 26660 14356 26666 14408
rect 26881 14399 26939 14405
rect 26881 14365 26893 14399
rect 26927 14396 26939 14399
rect 26970 14396 26976 14408
rect 26927 14368 26976 14396
rect 26927 14365 26939 14368
rect 26881 14359 26939 14365
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27062 14356 27068 14408
rect 27120 14356 27126 14408
rect 27157 14399 27215 14405
rect 27157 14365 27169 14399
rect 27203 14396 27215 14399
rect 27338 14396 27344 14408
rect 27203 14368 27344 14396
rect 27203 14365 27215 14368
rect 27157 14359 27215 14365
rect 27338 14356 27344 14368
rect 27396 14356 27402 14408
rect 28813 14399 28871 14405
rect 28813 14365 28825 14399
rect 28859 14396 28871 14399
rect 29549 14399 29607 14405
rect 29549 14396 29561 14399
rect 28859 14368 29561 14396
rect 28859 14365 28871 14368
rect 28813 14359 28871 14365
rect 29549 14365 29561 14368
rect 29595 14365 29607 14399
rect 29549 14359 29607 14365
rect 29638 14356 29644 14408
rect 29696 14396 29702 14408
rect 30024 14405 30052 14436
rect 30742 14424 30748 14476
rect 30800 14464 30806 14476
rect 30800 14436 31340 14464
rect 30800 14424 30806 14436
rect 29733 14399 29791 14405
rect 29733 14396 29745 14399
rect 29696 14368 29745 14396
rect 29696 14356 29702 14368
rect 29733 14365 29745 14368
rect 29779 14365 29791 14399
rect 29733 14359 29791 14365
rect 29825 14399 29883 14405
rect 29825 14365 29837 14399
rect 29871 14365 29883 14399
rect 29825 14359 29883 14365
rect 30009 14399 30067 14405
rect 30009 14365 30021 14399
rect 30055 14365 30067 14399
rect 30009 14359 30067 14365
rect 30193 14399 30251 14405
rect 30193 14365 30205 14399
rect 30239 14365 30251 14399
rect 30193 14359 30251 14365
rect 25409 14263 25467 14269
rect 25409 14229 25421 14263
rect 25455 14260 25467 14263
rect 25958 14260 25964 14272
rect 25455 14232 25964 14260
rect 25455 14229 25467 14232
rect 25409 14223 25467 14229
rect 25958 14220 25964 14232
rect 26016 14220 26022 14272
rect 26620 14260 26648 14356
rect 27516 14331 27574 14337
rect 27516 14297 27528 14331
rect 27562 14328 27574 14331
rect 29365 14331 29423 14337
rect 29365 14328 29377 14331
rect 27562 14300 29377 14328
rect 27562 14297 27574 14300
rect 27516 14291 27574 14297
rect 29365 14297 29377 14300
rect 29411 14297 29423 14331
rect 29365 14291 29423 14297
rect 27065 14263 27123 14269
rect 27065 14260 27077 14263
rect 26620 14232 27077 14260
rect 27065 14229 27077 14232
rect 27111 14229 27123 14263
rect 27065 14223 27123 14229
rect 28626 14220 28632 14272
rect 28684 14260 28690 14272
rect 29840 14260 29868 14359
rect 30208 14328 30236 14359
rect 31110 14356 31116 14408
rect 31168 14396 31174 14408
rect 31312 14405 31340 14436
rect 31205 14399 31263 14405
rect 31205 14396 31217 14399
rect 31168 14368 31217 14396
rect 31168 14356 31174 14368
rect 31205 14365 31217 14368
rect 31251 14365 31263 14399
rect 31205 14359 31263 14365
rect 31297 14399 31355 14405
rect 31297 14365 31309 14399
rect 31343 14365 31355 14399
rect 31297 14359 31355 14365
rect 31478 14356 31484 14408
rect 31536 14356 31542 14408
rect 31573 14399 31631 14405
rect 31573 14365 31585 14399
rect 31619 14396 31631 14399
rect 31726 14396 31754 14572
rect 31846 14560 31852 14572
rect 31904 14560 31910 14612
rect 33134 14560 33140 14612
rect 33192 14560 33198 14612
rect 33594 14560 33600 14612
rect 33652 14560 33658 14612
rect 34422 14560 34428 14612
rect 34480 14560 34486 14612
rect 34517 14603 34575 14609
rect 34517 14569 34529 14603
rect 34563 14600 34575 14603
rect 34606 14600 34612 14612
rect 34563 14572 34612 14600
rect 34563 14569 34575 14572
rect 34517 14563 34575 14569
rect 34606 14560 34612 14572
rect 34664 14560 34670 14612
rect 34701 14603 34759 14609
rect 34701 14569 34713 14603
rect 34747 14600 34759 14603
rect 34790 14600 34796 14612
rect 34747 14572 34796 14600
rect 34747 14569 34759 14572
rect 34701 14563 34759 14569
rect 34790 14560 34796 14572
rect 34848 14560 34854 14612
rect 36446 14560 36452 14612
rect 36504 14560 36510 14612
rect 37090 14560 37096 14612
rect 37148 14600 37154 14612
rect 37148 14572 39620 14600
rect 37148 14560 37154 14572
rect 31619 14368 31754 14396
rect 31619 14365 31631 14368
rect 31573 14359 31631 14365
rect 31938 14356 31944 14408
rect 31996 14356 32002 14408
rect 32585 14399 32643 14405
rect 32585 14365 32597 14399
rect 32631 14396 32643 14399
rect 32950 14396 32956 14408
rect 32631 14368 32956 14396
rect 32631 14365 32643 14368
rect 32585 14359 32643 14365
rect 32950 14356 32956 14368
rect 33008 14356 33014 14408
rect 33318 14356 33324 14408
rect 33376 14356 33382 14408
rect 30208 14300 32628 14328
rect 28684 14232 29868 14260
rect 28684 14220 28690 14232
rect 32490 14220 32496 14272
rect 32548 14220 32554 14272
rect 32600 14260 32628 14300
rect 32674 14288 32680 14340
rect 32732 14328 32738 14340
rect 32861 14331 32919 14337
rect 32861 14328 32873 14331
rect 32732 14300 32873 14328
rect 32732 14288 32738 14300
rect 32861 14297 32873 14300
rect 32907 14297 32919 14331
rect 33612 14328 33640 14560
rect 34440 14532 34468 14560
rect 34440 14504 39436 14532
rect 33962 14424 33968 14476
rect 34020 14424 34026 14476
rect 36354 14464 36360 14476
rect 34532 14436 35011 14464
rect 34532 14408 34560 14436
rect 34514 14356 34520 14408
rect 34572 14356 34578 14408
rect 34698 14356 34704 14408
rect 34756 14396 34762 14408
rect 34885 14399 34943 14405
rect 34885 14396 34897 14399
rect 34756 14368 34897 14396
rect 34756 14356 34762 14368
rect 34885 14365 34897 14368
rect 34931 14365 34943 14399
rect 34983 14396 35011 14436
rect 36188 14436 36360 14464
rect 35187 14399 35245 14405
rect 35187 14396 35199 14399
rect 34983 14368 35199 14396
rect 34885 14359 34943 14365
rect 35187 14365 35199 14368
rect 35233 14365 35245 14399
rect 35187 14359 35245 14365
rect 35342 14356 35348 14408
rect 35400 14356 35406 14408
rect 36188 14405 36216 14436
rect 36354 14424 36360 14436
rect 36412 14424 36418 14476
rect 36722 14424 36728 14476
rect 36780 14424 36786 14476
rect 36173 14399 36231 14405
rect 36173 14396 36185 14399
rect 35452 14368 36185 14396
rect 34977 14331 35035 14337
rect 34977 14328 34989 14331
rect 33612 14300 34989 14328
rect 32861 14291 32919 14297
rect 34977 14297 34989 14300
rect 35023 14297 35035 14331
rect 34977 14291 35035 14297
rect 32766 14260 32772 14272
rect 32600 14232 32772 14260
rect 32766 14220 32772 14232
rect 32824 14220 32830 14272
rect 34992 14260 35020 14291
rect 35066 14288 35072 14340
rect 35124 14288 35130 14340
rect 35452 14260 35480 14368
rect 36173 14365 36185 14368
rect 36219 14365 36231 14399
rect 36173 14359 36231 14365
rect 36265 14399 36323 14405
rect 36265 14365 36277 14399
rect 36311 14396 36323 14399
rect 36998 14396 37004 14408
rect 36311 14368 37004 14396
rect 36311 14365 36323 14368
rect 36265 14359 36323 14365
rect 36998 14356 37004 14368
rect 37056 14396 37062 14408
rect 37277 14399 37335 14405
rect 37277 14396 37289 14399
rect 37056 14368 37289 14396
rect 37056 14356 37062 14368
rect 37277 14365 37289 14368
rect 37323 14365 37335 14399
rect 37277 14359 37335 14365
rect 37458 14288 37464 14340
rect 37516 14288 37522 14340
rect 39408 14328 39436 14504
rect 39482 14492 39488 14544
rect 39540 14492 39546 14544
rect 39592 14532 39620 14572
rect 39758 14560 39764 14612
rect 39816 14600 39822 14612
rect 40494 14600 40500 14612
rect 39816 14572 40500 14600
rect 39816 14560 39822 14572
rect 40494 14560 40500 14572
rect 40552 14560 40558 14612
rect 40678 14560 40684 14612
rect 40736 14600 40742 14612
rect 42153 14603 42211 14609
rect 42153 14600 42165 14603
rect 40736 14572 42165 14600
rect 40736 14560 40742 14572
rect 42153 14569 42165 14572
rect 42199 14569 42211 14603
rect 42153 14563 42211 14569
rect 42242 14560 42248 14612
rect 42300 14560 42306 14612
rect 42886 14560 42892 14612
rect 42944 14560 42950 14612
rect 46566 14560 46572 14612
rect 46624 14600 46630 14612
rect 46937 14603 46995 14609
rect 46937 14600 46949 14603
rect 46624 14572 46949 14600
rect 46624 14560 46630 14572
rect 46937 14569 46949 14572
rect 46983 14569 46995 14603
rect 46937 14563 46995 14569
rect 47210 14560 47216 14612
rect 47268 14560 47274 14612
rect 47486 14560 47492 14612
rect 47544 14560 47550 14612
rect 47578 14560 47584 14612
rect 47636 14560 47642 14612
rect 47765 14603 47823 14609
rect 47765 14569 47777 14603
rect 47811 14600 47823 14603
rect 48958 14600 48964 14612
rect 47811 14572 48964 14600
rect 47811 14569 47823 14572
rect 47765 14563 47823 14569
rect 48958 14560 48964 14572
rect 49016 14560 49022 14612
rect 49142 14560 49148 14612
rect 49200 14600 49206 14612
rect 49513 14603 49571 14609
rect 49513 14600 49525 14603
rect 49200 14572 49525 14600
rect 49200 14560 49206 14572
rect 49513 14569 49525 14572
rect 49559 14569 49571 14603
rect 49513 14563 49571 14569
rect 49694 14560 49700 14612
rect 49752 14560 49758 14612
rect 51077 14603 51135 14609
rect 51077 14569 51089 14603
rect 51123 14600 51135 14603
rect 51258 14600 51264 14612
rect 51123 14572 51264 14600
rect 51123 14569 51135 14572
rect 51077 14563 51135 14569
rect 51258 14560 51264 14572
rect 51316 14560 51322 14612
rect 51994 14560 52000 14612
rect 52052 14600 52058 14612
rect 52638 14600 52644 14612
rect 52052 14572 52644 14600
rect 52052 14560 52058 14572
rect 52638 14560 52644 14572
rect 52696 14560 52702 14612
rect 52825 14603 52883 14609
rect 52825 14569 52837 14603
rect 52871 14600 52883 14603
rect 53466 14600 53472 14612
rect 52871 14572 53472 14600
rect 52871 14569 52883 14572
rect 52825 14563 52883 14569
rect 53466 14560 53472 14572
rect 53524 14560 53530 14612
rect 42260 14532 42288 14560
rect 39592 14504 42288 14532
rect 42337 14535 42395 14541
rect 42337 14501 42349 14535
rect 42383 14532 42395 14535
rect 42702 14532 42708 14544
rect 42383 14504 42708 14532
rect 42383 14501 42395 14504
rect 42337 14495 42395 14501
rect 42702 14492 42708 14504
rect 42760 14492 42766 14544
rect 42794 14492 42800 14544
rect 42852 14532 42858 14544
rect 43717 14535 43775 14541
rect 43717 14532 43729 14535
rect 42852 14504 43729 14532
rect 42852 14492 42858 14504
rect 39500 14464 39528 14492
rect 40218 14464 40224 14476
rect 39500 14436 40224 14464
rect 40218 14424 40224 14436
rect 40276 14464 40282 14476
rect 40589 14467 40647 14473
rect 40589 14464 40601 14467
rect 40276 14436 40601 14464
rect 40276 14424 40282 14436
rect 40589 14433 40601 14436
rect 40635 14433 40647 14467
rect 40589 14427 40647 14433
rect 39666 14356 39672 14408
rect 39724 14396 39730 14408
rect 39853 14399 39911 14405
rect 39853 14396 39865 14399
rect 39724 14368 39865 14396
rect 39724 14356 39730 14368
rect 39853 14365 39865 14368
rect 39899 14365 39911 14399
rect 39853 14359 39911 14365
rect 41601 14399 41659 14405
rect 41601 14365 41613 14399
rect 41647 14396 41659 14399
rect 42518 14396 42524 14408
rect 41647 14368 42288 14396
rect 42479 14368 42524 14396
rect 41647 14365 41659 14368
rect 41601 14359 41659 14365
rect 40310 14328 40316 14340
rect 39408 14300 40316 14328
rect 40310 14288 40316 14300
rect 40368 14288 40374 14340
rect 42260 14272 42288 14368
rect 42518 14356 42524 14368
rect 42576 14356 42582 14408
rect 42904 14396 42932 14504
rect 43717 14501 43729 14504
rect 43763 14532 43775 14535
rect 47228 14532 47256 14560
rect 43763 14504 47256 14532
rect 43763 14501 43775 14504
rect 43717 14495 43775 14501
rect 47302 14492 47308 14544
rect 47360 14492 47366 14544
rect 47394 14492 47400 14544
rect 47452 14492 47458 14544
rect 45554 14464 45560 14476
rect 43180 14436 45560 14464
rect 42981 14399 43039 14405
rect 42981 14396 42993 14399
rect 42904 14368 42993 14396
rect 42981 14365 42993 14368
rect 43027 14365 43039 14399
rect 42981 14359 43039 14365
rect 43070 14356 43076 14408
rect 43128 14356 43134 14408
rect 43180 14328 43208 14436
rect 45554 14424 45560 14436
rect 45612 14424 45618 14476
rect 46474 14424 46480 14476
rect 46532 14464 46538 14476
rect 46750 14464 46756 14476
rect 46532 14436 46756 14464
rect 46532 14424 46538 14436
rect 46750 14424 46756 14436
rect 46808 14464 46814 14476
rect 47504 14464 47532 14560
rect 46808 14436 47164 14464
rect 46808 14424 46814 14436
rect 43257 14399 43315 14405
rect 43257 14365 43269 14399
rect 43303 14365 43315 14399
rect 43257 14359 43315 14365
rect 43625 14399 43683 14405
rect 43625 14365 43637 14399
rect 43671 14396 43683 14399
rect 43806 14396 43812 14408
rect 43671 14368 43812 14396
rect 43671 14365 43683 14368
rect 43625 14359 43683 14365
rect 42536 14300 43208 14328
rect 43272 14328 43300 14359
rect 43806 14356 43812 14368
rect 43864 14356 43870 14408
rect 44082 14356 44088 14408
rect 44140 14356 44146 14408
rect 46385 14399 46443 14405
rect 46385 14365 46397 14399
rect 46431 14396 46443 14399
rect 47029 14399 47087 14405
rect 47029 14396 47041 14399
rect 46431 14368 47041 14396
rect 46431 14365 46443 14368
rect 46385 14359 46443 14365
rect 47029 14365 47041 14368
rect 47075 14365 47087 14399
rect 47029 14359 47087 14365
rect 44100 14328 44128 14356
rect 43272 14300 44128 14328
rect 47136 14328 47164 14436
rect 47228 14436 47532 14464
rect 47228 14405 47256 14436
rect 47213 14399 47271 14405
rect 47213 14365 47225 14399
rect 47259 14365 47271 14399
rect 47213 14359 47271 14365
rect 47489 14399 47547 14405
rect 47489 14365 47501 14399
rect 47535 14365 47547 14399
rect 47596 14396 47624 14560
rect 48682 14492 48688 14544
rect 48740 14532 48746 14544
rect 48866 14532 48872 14544
rect 48740 14504 48872 14532
rect 48740 14492 48746 14504
rect 48866 14492 48872 14504
rect 48924 14532 48930 14544
rect 49237 14535 49295 14541
rect 49237 14532 49249 14535
rect 48924 14504 49249 14532
rect 48924 14492 48930 14504
rect 49237 14501 49249 14504
rect 49283 14501 49295 14535
rect 49237 14495 49295 14501
rect 49712 14464 49740 14560
rect 48240 14436 49740 14464
rect 51092 14436 52592 14464
rect 47673 14399 47731 14405
rect 47673 14396 47685 14399
rect 47596 14368 47685 14396
rect 47489 14359 47547 14365
rect 47673 14365 47685 14368
rect 47719 14365 47731 14399
rect 47673 14359 47731 14365
rect 48133 14399 48191 14405
rect 48133 14365 48145 14399
rect 48179 14365 48191 14399
rect 48240 14398 48268 14436
rect 48317 14399 48375 14405
rect 48317 14398 48329 14399
rect 48240 14370 48329 14398
rect 48133 14359 48191 14365
rect 48317 14365 48329 14370
rect 48363 14365 48375 14399
rect 48317 14359 48375 14365
rect 48409 14399 48467 14405
rect 48409 14365 48421 14399
rect 48455 14365 48467 14399
rect 48409 14359 48467 14365
rect 48593 14399 48651 14405
rect 48593 14365 48605 14399
rect 48639 14396 48651 14399
rect 48866 14396 48872 14408
rect 48639 14368 48872 14396
rect 48639 14365 48651 14368
rect 48593 14359 48651 14365
rect 47504 14328 47532 14359
rect 47136 14300 47532 14328
rect 48148 14328 48176 14359
rect 48424 14328 48452 14359
rect 48866 14356 48872 14368
rect 48924 14356 48930 14408
rect 49053 14399 49111 14405
rect 49053 14365 49065 14399
rect 49099 14365 49111 14399
rect 49053 14359 49111 14365
rect 48682 14328 48688 14340
rect 48148 14300 48688 14328
rect 34992 14232 35480 14260
rect 35805 14263 35863 14269
rect 35805 14229 35817 14263
rect 35851 14260 35863 14263
rect 36722 14260 36728 14272
rect 35851 14232 36728 14260
rect 35851 14229 35863 14232
rect 35805 14223 35863 14229
rect 36722 14220 36728 14232
rect 36780 14220 36786 14272
rect 38562 14220 38568 14272
rect 38620 14260 38626 14272
rect 38749 14263 38807 14269
rect 38749 14260 38761 14263
rect 38620 14232 38761 14260
rect 38620 14220 38626 14232
rect 38749 14229 38761 14232
rect 38795 14229 38807 14263
rect 38749 14223 38807 14229
rect 40494 14220 40500 14272
rect 40552 14220 40558 14272
rect 41230 14220 41236 14272
rect 41288 14220 41294 14272
rect 42242 14220 42248 14272
rect 42300 14260 42306 14272
rect 42536 14269 42564 14300
rect 42521 14263 42579 14269
rect 42521 14260 42533 14263
rect 42300 14232 42533 14260
rect 42300 14220 42306 14232
rect 42521 14229 42533 14232
rect 42567 14229 42579 14263
rect 42521 14223 42579 14229
rect 43162 14220 43168 14272
rect 43220 14220 43226 14272
rect 45830 14220 45836 14272
rect 45888 14260 45894 14272
rect 48148 14260 48176 14300
rect 48682 14288 48688 14300
rect 48740 14288 48746 14340
rect 49068 14328 49096 14359
rect 49694 14356 49700 14408
rect 49752 14356 49758 14408
rect 49786 14356 49792 14408
rect 49844 14396 49850 14408
rect 49844 14368 50844 14396
rect 49844 14356 49850 14368
rect 50816 14340 50844 14368
rect 50982 14356 50988 14408
rect 51040 14356 51046 14408
rect 51092 14405 51120 14436
rect 52564 14408 52592 14436
rect 51077 14399 51135 14405
rect 51077 14365 51089 14399
rect 51123 14365 51135 14399
rect 51077 14359 51135 14365
rect 51442 14356 51448 14408
rect 51500 14396 51506 14408
rect 51537 14399 51595 14405
rect 51537 14396 51549 14399
rect 51500 14368 51549 14396
rect 51500 14356 51506 14368
rect 51537 14365 51549 14368
rect 51583 14365 51595 14399
rect 51537 14359 51595 14365
rect 51721 14399 51779 14405
rect 51721 14365 51733 14399
rect 51767 14396 51779 14399
rect 52454 14396 52460 14408
rect 51767 14368 52460 14396
rect 51767 14365 51779 14368
rect 51721 14359 51779 14365
rect 50154 14328 50160 14340
rect 49068 14300 50160 14328
rect 50154 14288 50160 14300
rect 50212 14288 50218 14340
rect 50614 14288 50620 14340
rect 50672 14288 50678 14340
rect 50798 14288 50804 14340
rect 50856 14288 50862 14340
rect 51736 14328 51764 14359
rect 52454 14356 52460 14368
rect 52512 14356 52518 14408
rect 52546 14356 52552 14408
rect 52604 14356 52610 14408
rect 52730 14356 52736 14408
rect 52788 14396 52794 14408
rect 52788 14368 53512 14396
rect 52788 14356 52794 14368
rect 53484 14340 53512 14368
rect 68462 14356 68468 14408
rect 68520 14356 68526 14408
rect 51046 14300 51764 14328
rect 45888 14232 48176 14260
rect 45888 14220 45894 14232
rect 48222 14220 48228 14272
rect 48280 14220 48286 14272
rect 48590 14220 48596 14272
rect 48648 14260 48654 14272
rect 51046 14260 51074 14300
rect 53466 14288 53472 14340
rect 53524 14288 53530 14340
rect 48648 14232 51074 14260
rect 48648 14220 48654 14232
rect 51258 14220 51264 14272
rect 51316 14220 51322 14272
rect 51626 14220 51632 14272
rect 51684 14220 51690 14272
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 27890 14016 27896 14068
rect 27948 14016 27954 14068
rect 28626 14016 28632 14068
rect 28684 14016 28690 14068
rect 31938 14016 31944 14068
rect 31996 14056 32002 14068
rect 33505 14059 33563 14065
rect 33505 14056 33517 14059
rect 31996 14028 33517 14056
rect 31996 14016 32002 14028
rect 33505 14025 33517 14028
rect 33551 14025 33563 14059
rect 33505 14019 33563 14025
rect 33597 14059 33655 14065
rect 33597 14025 33609 14059
rect 33643 14025 33655 14059
rect 33597 14019 33655 14025
rect 34333 14059 34391 14065
rect 34333 14025 34345 14059
rect 34379 14056 34391 14059
rect 34606 14056 34612 14068
rect 34379 14028 34612 14056
rect 34379 14025 34391 14028
rect 34333 14019 34391 14025
rect 23934 13948 23940 14000
rect 23992 13948 23998 14000
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13920 27859 13923
rect 27908 13920 27936 14016
rect 27847 13892 27936 13920
rect 27985 13923 28043 13929
rect 27847 13889 27859 13892
rect 27801 13883 27859 13889
rect 27985 13889 27997 13923
rect 28031 13889 28043 13923
rect 27985 13883 28043 13889
rect 28077 13923 28135 13929
rect 28077 13889 28089 13923
rect 28123 13920 28135 13923
rect 28644 13920 28672 14016
rect 33042 13988 33048 14000
rect 32140 13960 33048 13988
rect 29730 13929 29736 13932
rect 28123 13892 28672 13920
rect 28123 13889 28135 13892
rect 28077 13883 28135 13889
rect 29724 13883 29736 13929
rect 22370 13812 22376 13864
rect 22428 13852 22434 13864
rect 22925 13855 22983 13861
rect 22925 13852 22937 13855
rect 22428 13824 22937 13852
rect 22428 13812 22434 13824
rect 22925 13821 22937 13824
rect 22971 13821 22983 13855
rect 22925 13815 22983 13821
rect 23198 13812 23204 13864
rect 23256 13812 23262 13864
rect 24854 13812 24860 13864
rect 24912 13852 24918 13864
rect 24949 13855 25007 13861
rect 24949 13852 24961 13855
rect 24912 13824 24961 13852
rect 24912 13812 24918 13824
rect 24949 13821 24961 13824
rect 24995 13821 25007 13855
rect 28000 13852 28028 13883
rect 29730 13880 29736 13883
rect 29788 13880 29794 13932
rect 32140 13929 32168 13960
rect 33042 13948 33048 13960
rect 33100 13948 33106 14000
rect 32125 13923 32183 13929
rect 32125 13889 32137 13923
rect 32171 13889 32183 13923
rect 32125 13883 32183 13889
rect 32214 13880 32220 13932
rect 32272 13880 32278 13932
rect 32392 13923 32450 13929
rect 32392 13889 32404 13923
rect 32438 13920 32450 13923
rect 33612 13920 33640 14019
rect 34606 14016 34612 14028
rect 34664 14056 34670 14068
rect 35342 14056 35348 14068
rect 34664 14028 35348 14056
rect 34664 14016 34670 14028
rect 35342 14016 35348 14028
rect 35400 14016 35406 14068
rect 38657 14059 38715 14065
rect 38657 14056 38669 14059
rect 36464 14028 38669 14056
rect 32438 13892 33640 13920
rect 32438 13889 32450 13892
rect 32392 13883 32450 13889
rect 33778 13880 33784 13932
rect 33836 13880 33842 13932
rect 33873 13923 33931 13929
rect 33873 13889 33885 13923
rect 33919 13920 33931 13923
rect 33962 13920 33968 13932
rect 33919 13892 33968 13920
rect 33919 13889 33931 13892
rect 33873 13883 33931 13889
rect 33962 13880 33968 13892
rect 34020 13880 34026 13932
rect 34057 13923 34115 13929
rect 34057 13889 34069 13923
rect 34103 13889 34115 13923
rect 34057 13883 34115 13889
rect 28000 13824 28120 13852
rect 24949 13815 25007 13821
rect 28092 13784 28120 13824
rect 28166 13812 28172 13864
rect 28224 13812 28230 13864
rect 28350 13852 28356 13864
rect 28276 13824 28356 13852
rect 28276 13784 28304 13824
rect 28350 13812 28356 13824
rect 28408 13852 28414 13864
rect 28408 13824 28948 13852
rect 28408 13812 28414 13824
rect 28092 13756 28304 13784
rect 28920 13784 28948 13824
rect 28994 13812 29000 13864
rect 29052 13852 29058 13864
rect 29457 13855 29515 13861
rect 29457 13852 29469 13855
rect 29052 13824 29469 13852
rect 29052 13812 29058 13824
rect 29457 13821 29469 13824
rect 29503 13821 29515 13855
rect 31205 13855 31263 13861
rect 31205 13852 31217 13855
rect 29457 13815 29515 13821
rect 30852 13824 31217 13852
rect 30852 13793 30880 13824
rect 31205 13821 31217 13824
rect 31251 13852 31263 13855
rect 32232 13852 32260 13880
rect 31251 13824 32260 13852
rect 31251 13821 31263 13824
rect 31205 13815 31263 13821
rect 33226 13812 33232 13864
rect 33284 13852 33290 13864
rect 34072 13852 34100 13883
rect 34238 13880 34244 13932
rect 34296 13880 34302 13932
rect 34425 13923 34483 13929
rect 34425 13889 34437 13923
rect 34471 13889 34483 13923
rect 34425 13883 34483 13889
rect 34146 13852 34152 13864
rect 33284 13824 34152 13852
rect 33284 13812 33290 13824
rect 34146 13812 34152 13824
rect 34204 13812 34210 13864
rect 34440 13852 34468 13883
rect 36078 13880 36084 13932
rect 36136 13920 36142 13932
rect 36357 13923 36415 13929
rect 36357 13920 36369 13923
rect 36136 13892 36369 13920
rect 36136 13880 36142 13892
rect 36357 13889 36369 13892
rect 36403 13889 36415 13923
rect 36464 13920 36492 14028
rect 38657 14025 38669 14028
rect 38703 14056 38715 14059
rect 39022 14056 39028 14068
rect 38703 14028 39028 14056
rect 38703 14025 38715 14028
rect 38657 14019 38715 14025
rect 39022 14016 39028 14028
rect 39080 14056 39086 14068
rect 39758 14056 39764 14068
rect 39080 14028 39764 14056
rect 39080 14016 39086 14028
rect 39758 14016 39764 14028
rect 39816 14016 39822 14068
rect 40218 14016 40224 14068
rect 40276 14016 40282 14068
rect 40494 14016 40500 14068
rect 40552 14016 40558 14068
rect 42242 14016 42248 14068
rect 42300 14016 42306 14068
rect 43162 14016 43168 14068
rect 43220 14016 43226 14068
rect 44726 14016 44732 14068
rect 44784 14016 44790 14068
rect 45557 14059 45615 14065
rect 45557 14025 45569 14059
rect 45603 14056 45615 14059
rect 45646 14056 45652 14068
rect 45603 14028 45652 14056
rect 45603 14025 45615 14028
rect 45557 14019 45615 14025
rect 45646 14016 45652 14028
rect 45704 14016 45710 14068
rect 49602 14056 49608 14068
rect 48056 14028 49608 14056
rect 36541 13991 36599 13997
rect 36541 13957 36553 13991
rect 36587 13988 36599 13991
rect 36814 13988 36820 14000
rect 36587 13960 36820 13988
rect 36587 13957 36599 13960
rect 36541 13951 36599 13957
rect 36814 13948 36820 13960
rect 36872 13948 36878 14000
rect 36906 13948 36912 14000
rect 36964 13988 36970 14000
rect 37522 13991 37580 13997
rect 37522 13988 37534 13991
rect 36964 13960 37534 13988
rect 36964 13948 36970 13960
rect 37522 13957 37534 13960
rect 37568 13957 37580 13991
rect 37522 13951 37580 13957
rect 39108 13991 39166 13997
rect 39108 13957 39120 13991
rect 39154 13988 39166 13991
rect 40512 13988 40540 14016
rect 42696 13991 42754 13997
rect 39154 13960 40540 13988
rect 40880 13960 42472 13988
rect 39154 13957 39166 13960
rect 39108 13951 39166 13957
rect 36633 13923 36691 13929
rect 36633 13920 36645 13923
rect 36464 13892 36645 13920
rect 36357 13883 36415 13889
rect 36633 13889 36645 13892
rect 36679 13889 36691 13923
rect 36633 13883 36691 13889
rect 36722 13880 36728 13932
rect 36780 13920 36786 13932
rect 36780 13892 36958 13920
rect 36780 13880 36786 13892
rect 36538 13852 36544 13864
rect 34440 13824 36544 13852
rect 36538 13812 36544 13824
rect 36596 13852 36602 13864
rect 36930 13852 36958 13892
rect 37274 13880 37280 13932
rect 37332 13880 37338 13932
rect 38654 13920 38660 13932
rect 37375 13892 38660 13920
rect 37375 13852 37403 13892
rect 38654 13880 38660 13892
rect 38712 13880 38718 13932
rect 36596 13824 36860 13852
rect 36930 13824 37403 13852
rect 36596 13812 36602 13824
rect 30837 13787 30895 13793
rect 28920 13756 29040 13784
rect 27798 13676 27804 13728
rect 27856 13676 27862 13728
rect 29012 13716 29040 13756
rect 30837 13753 30849 13787
rect 30883 13753 30895 13787
rect 34330 13784 34336 13796
rect 30837 13747 30895 13753
rect 31128 13756 32168 13784
rect 31128 13728 31156 13756
rect 30098 13716 30104 13728
rect 29012 13688 30104 13716
rect 30098 13676 30104 13688
rect 30156 13676 30162 13728
rect 31110 13676 31116 13728
rect 31168 13676 31174 13728
rect 31662 13676 31668 13728
rect 31720 13716 31726 13728
rect 31757 13719 31815 13725
rect 31757 13716 31769 13719
rect 31720 13688 31769 13716
rect 31720 13676 31726 13688
rect 31757 13685 31769 13688
rect 31803 13685 31815 13719
rect 32140 13716 32168 13756
rect 33060 13756 34336 13784
rect 33060 13716 33088 13756
rect 34330 13744 34336 13756
rect 34388 13744 34394 13796
rect 32140 13688 33088 13716
rect 31757 13679 31815 13685
rect 33870 13676 33876 13728
rect 33928 13676 33934 13728
rect 36832 13716 36860 13824
rect 38838 13812 38844 13864
rect 38896 13812 38902 13864
rect 39850 13812 39856 13864
rect 39908 13852 39914 13864
rect 40880 13861 40908 13960
rect 40954 13880 40960 13932
rect 41012 13920 41018 13932
rect 41121 13923 41179 13929
rect 41121 13920 41133 13923
rect 41012 13892 41133 13920
rect 41012 13880 41018 13892
rect 41121 13889 41133 13892
rect 41167 13889 41179 13923
rect 41121 13883 41179 13889
rect 42444 13861 42472 13960
rect 42696 13957 42708 13991
rect 42742 13988 42754 13991
rect 43180 13988 43208 14016
rect 42742 13960 43208 13988
rect 44836 13960 46244 13988
rect 42742 13957 42754 13960
rect 42696 13951 42754 13957
rect 44836 13864 44864 13960
rect 46216 13929 46244 13960
rect 45649 13923 45707 13929
rect 45649 13889 45661 13923
rect 45695 13920 45707 13923
rect 46201 13923 46259 13929
rect 45695 13892 46060 13920
rect 45695 13889 45707 13892
rect 45649 13883 45707 13889
rect 40865 13855 40923 13861
rect 40865 13852 40877 13855
rect 39908 13824 40877 13852
rect 39908 13812 39914 13824
rect 40865 13821 40877 13824
rect 40911 13821 40923 13855
rect 40865 13815 40923 13821
rect 42429 13855 42487 13861
rect 42429 13821 42441 13855
rect 42475 13821 42487 13855
rect 42429 13815 42487 13821
rect 36906 13744 36912 13796
rect 36964 13744 36970 13796
rect 38746 13716 38752 13728
rect 36832 13688 38752 13716
rect 38746 13676 38752 13688
rect 38804 13716 38810 13728
rect 40770 13716 40776 13728
rect 38804 13688 40776 13716
rect 38804 13676 38810 13688
rect 40770 13676 40776 13688
rect 40828 13676 40834 13728
rect 42444 13716 42472 13815
rect 44818 13812 44824 13864
rect 44876 13812 44882 13864
rect 46032 13861 46060 13892
rect 46201 13889 46213 13923
rect 46247 13920 46259 13923
rect 46477 13923 46535 13929
rect 46477 13920 46489 13923
rect 46247 13892 46489 13920
rect 46247 13889 46259 13892
rect 46201 13883 46259 13889
rect 46477 13889 46489 13892
rect 46523 13889 46535 13923
rect 46477 13883 46535 13889
rect 46661 13923 46719 13929
rect 46661 13889 46673 13923
rect 46707 13920 46719 13923
rect 47210 13920 47216 13932
rect 46707 13892 47216 13920
rect 46707 13889 46719 13892
rect 46661 13883 46719 13889
rect 45005 13855 45063 13861
rect 45005 13821 45017 13855
rect 45051 13821 45063 13855
rect 45005 13815 45063 13821
rect 45833 13855 45891 13861
rect 45833 13821 45845 13855
rect 45879 13821 45891 13855
rect 45833 13815 45891 13821
rect 46017 13855 46075 13861
rect 46017 13821 46029 13855
rect 46063 13852 46075 13855
rect 46676 13852 46704 13883
rect 47210 13880 47216 13892
rect 47268 13880 47274 13932
rect 48056 13929 48084 14028
rect 49602 14016 49608 14028
rect 49660 14016 49666 14068
rect 49694 14016 49700 14068
rect 49752 14056 49758 14068
rect 50709 14059 50767 14065
rect 50709 14056 50721 14059
rect 49752 14028 50721 14056
rect 49752 14016 49758 14028
rect 50709 14025 50721 14028
rect 50755 14025 50767 14059
rect 50709 14019 50767 14025
rect 50798 14016 50804 14068
rect 50856 14056 50862 14068
rect 51905 14059 51963 14065
rect 51905 14056 51917 14059
rect 50856 14028 51917 14056
rect 50856 14016 50862 14028
rect 51905 14025 51917 14028
rect 51951 14025 51963 14059
rect 52365 14059 52423 14065
rect 52365 14056 52377 14059
rect 51905 14019 51963 14025
rect 52012 14028 52377 14056
rect 49786 13988 49792 14000
rect 48240 13960 49792 13988
rect 48240 13929 48268 13960
rect 49786 13948 49792 13960
rect 49844 13948 49850 14000
rect 51258 13988 51264 14000
rect 50080 13960 51264 13988
rect 48041 13923 48099 13929
rect 48041 13889 48053 13923
rect 48087 13889 48099 13923
rect 48041 13883 48099 13889
rect 48225 13923 48283 13929
rect 48225 13889 48237 13923
rect 48271 13889 48283 13923
rect 48225 13883 48283 13889
rect 48317 13923 48375 13929
rect 48317 13889 48329 13923
rect 48363 13920 48375 13923
rect 48406 13920 48412 13932
rect 48363 13892 48412 13920
rect 48363 13889 48375 13892
rect 48317 13883 48375 13889
rect 48406 13880 48412 13892
rect 48464 13880 48470 13932
rect 48501 13923 48559 13929
rect 48501 13889 48513 13923
rect 48547 13889 48559 13923
rect 48501 13883 48559 13889
rect 46063 13824 46704 13852
rect 46063 13821 46075 13824
rect 46017 13815 46075 13821
rect 43806 13744 43812 13796
rect 43864 13784 43870 13796
rect 44542 13784 44548 13796
rect 43864 13756 44548 13784
rect 43864 13744 43870 13756
rect 44542 13744 44548 13756
rect 44600 13784 44606 13796
rect 45020 13784 45048 13815
rect 45848 13784 45876 13815
rect 48130 13812 48136 13864
rect 48188 13812 48194 13864
rect 48516 13784 48544 13883
rect 48682 13880 48688 13932
rect 48740 13920 48746 13932
rect 48777 13923 48835 13929
rect 48777 13920 48789 13923
rect 48740 13892 48789 13920
rect 48740 13880 48746 13892
rect 48777 13889 48789 13892
rect 48823 13889 48835 13923
rect 48777 13883 48835 13889
rect 48866 13880 48872 13932
rect 48924 13880 48930 13932
rect 49053 13923 49111 13929
rect 49053 13889 49065 13923
rect 49099 13920 49111 13923
rect 49142 13920 49148 13932
rect 49099 13892 49148 13920
rect 49099 13889 49111 13892
rect 49053 13883 49111 13889
rect 49142 13880 49148 13892
rect 49200 13880 49206 13932
rect 49234 13880 49240 13932
rect 49292 13880 49298 13932
rect 50080 13929 50108 13960
rect 51258 13948 51264 13960
rect 51316 13948 51322 14000
rect 52012 13988 52040 14028
rect 52365 14025 52377 14028
rect 52411 14025 52423 14059
rect 52365 14019 52423 14025
rect 51476 13960 52040 13988
rect 52104 13960 52592 13988
rect 49697 13923 49755 13929
rect 49697 13889 49709 13923
rect 49743 13889 49755 13923
rect 49697 13883 49755 13889
rect 50065 13923 50123 13929
rect 50065 13889 50077 13923
rect 50111 13889 50123 13923
rect 50065 13883 50123 13889
rect 50157 13923 50215 13929
rect 50157 13889 50169 13923
rect 50203 13920 50215 13923
rect 50246 13920 50252 13932
rect 50203 13892 50252 13920
rect 50203 13889 50215 13892
rect 50157 13883 50215 13889
rect 48593 13855 48651 13861
rect 48593 13821 48605 13855
rect 48639 13852 48651 13855
rect 48884 13852 48912 13880
rect 48639 13824 48912 13852
rect 48961 13855 49019 13861
rect 48639 13821 48651 13824
rect 48593 13815 48651 13821
rect 48961 13821 48973 13855
rect 49007 13852 49019 13855
rect 49418 13852 49424 13864
rect 49007 13824 49424 13852
rect 49007 13821 49019 13824
rect 48961 13815 49019 13821
rect 44600 13756 48544 13784
rect 44600 13744 44606 13756
rect 42794 13716 42800 13728
rect 42444 13688 42800 13716
rect 42794 13676 42800 13688
rect 42852 13676 42858 13728
rect 44358 13676 44364 13728
rect 44416 13676 44422 13728
rect 45186 13676 45192 13728
rect 45244 13676 45250 13728
rect 46382 13676 46388 13728
rect 46440 13676 46446 13728
rect 46474 13676 46480 13728
rect 46532 13676 46538 13728
rect 47026 13676 47032 13728
rect 47084 13716 47090 13728
rect 47857 13719 47915 13725
rect 47857 13716 47869 13719
rect 47084 13688 47869 13716
rect 47084 13676 47090 13688
rect 47857 13685 47869 13688
rect 47903 13685 47915 13719
rect 47857 13679 47915 13685
rect 47946 13676 47952 13728
rect 48004 13716 48010 13728
rect 48608 13716 48636 13815
rect 49418 13812 49424 13824
rect 49476 13812 49482 13864
rect 49712 13852 49740 13883
rect 50246 13880 50252 13892
rect 50304 13880 50310 13932
rect 51077 13923 51135 13929
rect 51077 13889 51089 13923
rect 51123 13920 51135 13923
rect 51476 13920 51504 13960
rect 51123 13892 51504 13920
rect 51537 13923 51595 13929
rect 51123 13889 51135 13892
rect 51077 13883 51135 13889
rect 51537 13889 51549 13923
rect 51583 13889 51595 13923
rect 51537 13883 51595 13889
rect 51721 13923 51779 13929
rect 51721 13889 51733 13923
rect 51767 13920 51779 13923
rect 52104 13920 52132 13960
rect 52564 13932 52592 13960
rect 51767 13892 52132 13920
rect 52181 13923 52239 13929
rect 51767 13889 51779 13892
rect 51721 13883 51779 13889
rect 52181 13889 52193 13923
rect 52227 13889 52239 13923
rect 52181 13883 52239 13889
rect 50706 13852 50712 13864
rect 49712 13824 50712 13852
rect 50706 13812 50712 13824
rect 50764 13852 50770 13864
rect 50764 13824 51120 13852
rect 50764 13812 50770 13824
rect 50154 13744 50160 13796
rect 50212 13784 50218 13796
rect 50341 13787 50399 13793
rect 50341 13784 50353 13787
rect 50212 13756 50353 13784
rect 50212 13744 50218 13756
rect 50341 13753 50353 13756
rect 50387 13753 50399 13787
rect 51092 13784 51120 13824
rect 51166 13812 51172 13864
rect 51224 13812 51230 13864
rect 51261 13855 51319 13861
rect 51261 13821 51273 13855
rect 51307 13852 51319 13855
rect 51552 13852 51580 13883
rect 51307 13824 51580 13852
rect 51307 13821 51319 13824
rect 51261 13815 51319 13821
rect 51276 13784 51304 13815
rect 51810 13812 51816 13864
rect 51868 13852 51874 13864
rect 51997 13855 52055 13861
rect 51997 13852 52009 13855
rect 51868 13824 52009 13852
rect 51868 13812 51874 13824
rect 51997 13821 52009 13824
rect 52043 13821 52055 13855
rect 51997 13815 52055 13821
rect 51092 13756 51304 13784
rect 50341 13747 50399 13753
rect 51718 13744 51724 13796
rect 51776 13784 51782 13796
rect 52196 13784 52224 13883
rect 52546 13880 52552 13932
rect 52604 13880 52610 13932
rect 51776 13756 52224 13784
rect 51776 13744 51782 13756
rect 48004 13688 48636 13716
rect 48004 13676 48010 13688
rect 48774 13676 48780 13728
rect 48832 13716 48838 13728
rect 49421 13719 49479 13725
rect 49421 13716 49433 13719
rect 48832 13688 49433 13716
rect 48832 13676 48838 13688
rect 49421 13685 49433 13688
rect 49467 13716 49479 13719
rect 49789 13719 49847 13725
rect 49789 13716 49801 13719
rect 49467 13688 49801 13716
rect 49467 13685 49479 13688
rect 49421 13679 49479 13685
rect 49789 13685 49801 13688
rect 49835 13685 49847 13719
rect 49789 13679 49847 13685
rect 51350 13676 51356 13728
rect 51408 13716 51414 13728
rect 51537 13719 51595 13725
rect 51537 13716 51549 13719
rect 51408 13688 51549 13716
rect 51408 13676 51414 13688
rect 51537 13685 51549 13688
rect 51583 13685 51595 13719
rect 51537 13679 51595 13685
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 23198 13472 23204 13524
rect 23256 13512 23262 13524
rect 23385 13515 23443 13521
rect 23385 13512 23397 13515
rect 23256 13484 23397 13512
rect 23256 13472 23262 13484
rect 23385 13481 23397 13484
rect 23431 13481 23443 13515
rect 23385 13475 23443 13481
rect 23934 13472 23940 13524
rect 23992 13472 23998 13524
rect 29641 13515 29699 13521
rect 29641 13481 29653 13515
rect 29687 13512 29699 13515
rect 29730 13512 29736 13524
rect 29687 13484 29736 13512
rect 29687 13481 29699 13484
rect 29641 13475 29699 13481
rect 29730 13472 29736 13484
rect 29788 13472 29794 13524
rect 31941 13515 31999 13521
rect 31941 13481 31953 13515
rect 31987 13512 31999 13515
rect 33318 13512 33324 13524
rect 31987 13484 33324 13512
rect 31987 13481 31999 13484
rect 31941 13475 31999 13481
rect 33318 13472 33324 13484
rect 33376 13472 33382 13524
rect 39206 13472 39212 13524
rect 39264 13472 39270 13524
rect 39393 13515 39451 13521
rect 39393 13481 39405 13515
rect 39439 13512 39451 13515
rect 39574 13512 39580 13524
rect 39439 13484 39580 13512
rect 39439 13481 39451 13484
rect 39393 13475 39451 13481
rect 39574 13472 39580 13484
rect 39632 13472 39638 13524
rect 39666 13472 39672 13524
rect 39724 13472 39730 13524
rect 40494 13512 40500 13524
rect 39868 13484 40500 13512
rect 24946 13404 24952 13456
rect 25004 13404 25010 13456
rect 32033 13447 32091 13453
rect 32033 13444 32045 13447
rect 30944 13416 32045 13444
rect 25501 13379 25559 13385
rect 25501 13376 25513 13379
rect 22388 13348 25513 13376
rect 22388 13320 22416 13348
rect 25501 13345 25513 13348
rect 25547 13376 25559 13379
rect 27062 13376 27068 13388
rect 25547 13348 27068 13376
rect 25547 13345 25559 13348
rect 25501 13339 25559 13345
rect 27062 13336 27068 13348
rect 27120 13336 27126 13388
rect 30098 13376 30104 13388
rect 29840 13348 30104 13376
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 992 13280 1593 13308
rect 992 13268 998 13280
rect 1581 13277 1593 13280
rect 1627 13277 1639 13311
rect 1581 13271 1639 13277
rect 22370 13268 22376 13320
rect 22428 13268 22434 13320
rect 23566 13268 23572 13320
rect 23624 13268 23630 13320
rect 23842 13268 23848 13320
rect 23900 13268 23906 13320
rect 29840 13317 29868 13348
rect 30098 13336 30104 13348
rect 30156 13336 30162 13388
rect 30944 13385 30972 13416
rect 32033 13413 32045 13416
rect 32079 13413 32091 13447
rect 32033 13407 32091 13413
rect 39485 13447 39543 13453
rect 39485 13413 39497 13447
rect 39531 13444 39543 13447
rect 39684 13444 39712 13472
rect 39531 13416 39712 13444
rect 39531 13413 39543 13416
rect 39485 13407 39543 13413
rect 30929 13379 30987 13385
rect 30929 13345 30941 13379
rect 30975 13345 30987 13379
rect 30929 13339 30987 13345
rect 31478 13336 31484 13388
rect 31536 13336 31542 13388
rect 31573 13379 31631 13385
rect 31573 13345 31585 13379
rect 31619 13376 31631 13379
rect 31662 13376 31668 13388
rect 31619 13348 31668 13376
rect 31619 13345 31631 13348
rect 31573 13339 31631 13345
rect 31662 13336 31668 13348
rect 31720 13336 31726 13388
rect 31938 13376 31944 13388
rect 31772 13348 31944 13376
rect 25133 13311 25191 13317
rect 25133 13277 25145 13311
rect 25179 13277 25191 13311
rect 25133 13271 25191 13277
rect 29641 13311 29699 13317
rect 29641 13277 29653 13311
rect 29687 13277 29699 13311
rect 29641 13271 29699 13277
rect 29825 13311 29883 13317
rect 29825 13277 29837 13311
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 24854 13200 24860 13252
rect 24912 13240 24918 13252
rect 24912 13212 24992 13240
rect 24912 13200 24918 13212
rect 24964 13172 24992 13212
rect 25038 13200 25044 13252
rect 25096 13200 25102 13252
rect 25148 13240 25176 13271
rect 25314 13240 25320 13252
rect 25148 13212 25320 13240
rect 25314 13200 25320 13212
rect 25372 13200 25378 13252
rect 25774 13200 25780 13252
rect 25832 13200 25838 13252
rect 26510 13200 26516 13252
rect 26568 13200 26574 13252
rect 27525 13243 27583 13249
rect 27525 13209 27537 13243
rect 27571 13209 27583 13243
rect 29656 13240 29684 13271
rect 30006 13268 30012 13320
rect 30064 13268 30070 13320
rect 30116 13308 30144 13336
rect 31496 13308 31524 13336
rect 31772 13317 31800 13348
rect 31938 13336 31944 13348
rect 31996 13336 32002 13388
rect 32324 13348 32904 13376
rect 30116 13280 31524 13308
rect 31757 13311 31815 13317
rect 31757 13277 31769 13311
rect 31803 13277 31815 13311
rect 31757 13271 31815 13277
rect 32214 13268 32220 13320
rect 32272 13268 32278 13320
rect 32324 13317 32352 13348
rect 32309 13311 32367 13317
rect 32309 13277 32321 13311
rect 32355 13277 32367 13311
rect 32309 13271 32367 13277
rect 32398 13268 32404 13320
rect 32456 13268 32462 13320
rect 32490 13268 32496 13320
rect 32548 13268 32554 13320
rect 31481 13243 31539 13249
rect 31481 13240 31493 13243
rect 29656 13212 31493 13240
rect 27525 13203 27583 13209
rect 31481 13209 31493 13212
rect 31527 13209 31539 13243
rect 31481 13203 31539 13209
rect 32033 13243 32091 13249
rect 32033 13209 32045 13243
rect 32079 13240 32091 13243
rect 32508 13240 32536 13268
rect 32876 13252 32904 13348
rect 38838 13336 38844 13388
rect 38896 13376 38902 13388
rect 39577 13379 39635 13385
rect 38896 13348 39528 13376
rect 38896 13336 38902 13348
rect 33042 13268 33048 13320
rect 33100 13308 33106 13320
rect 33137 13311 33195 13317
rect 33137 13308 33149 13311
rect 33100 13280 33149 13308
rect 33100 13268 33106 13280
rect 33137 13277 33149 13280
rect 33183 13308 33195 13311
rect 35069 13311 35127 13317
rect 35069 13308 35081 13311
rect 33183 13280 35081 13308
rect 33183 13277 33195 13280
rect 33137 13271 33195 13277
rect 35069 13277 35081 13280
rect 35115 13308 35127 13311
rect 37093 13311 37151 13317
rect 37093 13308 37105 13311
rect 35115 13280 37105 13308
rect 35115 13277 35127 13280
rect 35069 13271 35127 13277
rect 37093 13277 37105 13280
rect 37139 13277 37151 13311
rect 37093 13271 37151 13277
rect 38657 13311 38715 13317
rect 38657 13277 38669 13311
rect 38703 13308 38715 13311
rect 39301 13311 39359 13317
rect 39301 13308 39313 13311
rect 38703 13280 39313 13308
rect 38703 13277 38715 13280
rect 38657 13271 38715 13277
rect 39301 13277 39313 13280
rect 39347 13277 39359 13311
rect 39500 13308 39528 13348
rect 39577 13345 39589 13379
rect 39623 13376 39635 13379
rect 39868 13376 39896 13484
rect 40494 13472 40500 13484
rect 40552 13512 40558 13524
rect 44818 13521 44824 13524
rect 41969 13515 42027 13521
rect 41969 13512 41981 13515
rect 40552 13484 41981 13512
rect 40552 13472 40558 13484
rect 41969 13481 41981 13484
rect 42015 13481 42027 13515
rect 41969 13475 42027 13481
rect 44775 13515 44824 13521
rect 44775 13481 44787 13515
rect 44821 13481 44824 13515
rect 44775 13475 44824 13481
rect 44818 13472 44824 13475
rect 44876 13472 44882 13524
rect 48222 13512 48228 13524
rect 45388 13484 48228 13512
rect 40862 13404 40868 13456
rect 40920 13444 40926 13456
rect 40920 13416 41414 13444
rect 40920 13404 40926 13416
rect 39623 13348 39896 13376
rect 39623 13345 39635 13348
rect 39577 13339 39635 13345
rect 39850 13308 39856 13320
rect 39500 13280 39856 13308
rect 39301 13271 39359 13277
rect 32079 13212 32536 13240
rect 32079 13209 32091 13212
rect 32033 13203 32091 13209
rect 25498 13172 25504 13184
rect 24964 13144 25504 13172
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 26694 13132 26700 13184
rect 26752 13172 26758 13184
rect 27540 13172 27568 13203
rect 32858 13200 32864 13252
rect 32916 13200 32922 13252
rect 33404 13243 33462 13249
rect 33404 13209 33416 13243
rect 33450 13240 33462 13243
rect 34054 13240 34060 13252
rect 33450 13212 34060 13240
rect 33450 13209 33462 13212
rect 33404 13203 33462 13209
rect 34054 13200 34060 13212
rect 34112 13200 34118 13252
rect 35336 13243 35394 13249
rect 35336 13209 35348 13243
rect 35382 13240 35394 13243
rect 36262 13240 36268 13252
rect 35382 13212 36268 13240
rect 35382 13209 35394 13212
rect 35336 13203 35394 13209
rect 36262 13200 36268 13212
rect 36320 13200 36326 13252
rect 37360 13243 37418 13249
rect 37360 13209 37372 13243
rect 37406 13240 37418 13243
rect 37642 13240 37648 13252
rect 37406 13212 37648 13240
rect 37406 13209 37418 13212
rect 37360 13203 37418 13209
rect 37642 13200 37648 13212
rect 37700 13200 37706 13252
rect 26752 13144 27568 13172
rect 26752 13132 26758 13144
rect 30558 13132 30564 13184
rect 30616 13132 30622 13184
rect 32122 13132 32128 13184
rect 32180 13172 32186 13184
rect 33045 13175 33103 13181
rect 33045 13172 33057 13175
rect 32180 13144 33057 13172
rect 32180 13132 32186 13144
rect 33045 13141 33057 13144
rect 33091 13141 33103 13175
rect 33045 13135 33103 13141
rect 34422 13132 34428 13184
rect 34480 13172 34486 13184
rect 34517 13175 34575 13181
rect 34517 13172 34529 13175
rect 34480 13144 34529 13172
rect 34480 13132 34486 13144
rect 34517 13141 34529 13144
rect 34563 13141 34575 13175
rect 34517 13135 34575 13141
rect 36446 13132 36452 13184
rect 36504 13132 36510 13184
rect 38473 13175 38531 13181
rect 38473 13141 38485 13175
rect 38519 13172 38531 13175
rect 38672 13172 38700 13271
rect 39850 13268 39856 13280
rect 39908 13268 39914 13320
rect 40120 13243 40178 13249
rect 40120 13209 40132 13243
rect 40166 13240 40178 13243
rect 41046 13240 41052 13252
rect 40166 13212 41052 13240
rect 40166 13209 40178 13212
rect 40120 13203 40178 13209
rect 41046 13200 41052 13212
rect 41104 13200 41110 13252
rect 41386 13240 41414 13416
rect 42518 13376 42524 13388
rect 41984 13348 42524 13376
rect 41984 13317 42012 13348
rect 42518 13336 42524 13348
rect 42576 13376 42582 13388
rect 42889 13379 42947 13385
rect 42889 13376 42901 13379
rect 42576 13348 42901 13376
rect 42576 13336 42582 13348
rect 42889 13345 42901 13348
rect 42935 13345 42947 13379
rect 42889 13339 42947 13345
rect 43349 13379 43407 13385
rect 43349 13345 43361 13379
rect 43395 13376 43407 13379
rect 45388 13376 45416 13484
rect 48222 13472 48228 13484
rect 48280 13472 48286 13524
rect 48317 13515 48375 13521
rect 48317 13481 48329 13515
rect 48363 13481 48375 13515
rect 48317 13475 48375 13481
rect 47210 13404 47216 13456
rect 47268 13444 47274 13456
rect 47946 13444 47952 13456
rect 47268 13416 47952 13444
rect 47268 13404 47274 13416
rect 47946 13404 47952 13416
rect 48004 13404 48010 13456
rect 48130 13404 48136 13456
rect 48188 13444 48194 13456
rect 48332 13444 48360 13475
rect 48774 13472 48780 13524
rect 48832 13472 48838 13524
rect 49786 13472 49792 13524
rect 49844 13472 49850 13524
rect 51261 13515 51319 13521
rect 51261 13481 51273 13515
rect 51307 13512 51319 13515
rect 51442 13512 51448 13524
rect 51307 13484 51448 13512
rect 51307 13481 51319 13484
rect 51261 13475 51319 13481
rect 51442 13472 51448 13484
rect 51500 13512 51506 13524
rect 51718 13512 51724 13524
rect 51500 13484 51724 13512
rect 51500 13472 51506 13484
rect 51718 13472 51724 13484
rect 51776 13472 51782 13524
rect 48188 13416 48360 13444
rect 48188 13404 48194 13416
rect 49142 13404 49148 13456
rect 49200 13404 49206 13456
rect 50982 13444 50988 13456
rect 49436 13416 50988 13444
rect 43395 13348 45416 13376
rect 45465 13379 45523 13385
rect 43395 13345 43407 13348
rect 43349 13339 43407 13345
rect 45465 13345 45477 13379
rect 45511 13376 45523 13379
rect 46106 13376 46112 13388
rect 45511 13348 46112 13376
rect 45511 13345 45523 13348
rect 45465 13339 45523 13345
rect 46106 13336 46112 13348
rect 46164 13336 46170 13388
rect 49160 13376 49188 13404
rect 47780 13348 48544 13376
rect 41969 13311 42027 13317
rect 41969 13277 41981 13311
rect 42015 13277 42027 13311
rect 41969 13271 42027 13277
rect 42153 13311 42211 13317
rect 42153 13277 42165 13311
rect 42199 13308 42211 13311
rect 42242 13308 42248 13320
rect 42199 13280 42248 13308
rect 42199 13277 42211 13280
rect 42153 13271 42211 13277
rect 42168 13240 42196 13271
rect 42242 13268 42248 13280
rect 42300 13268 42306 13320
rect 42334 13268 42340 13320
rect 42392 13268 42398 13320
rect 42978 13268 42984 13320
rect 43036 13268 43042 13320
rect 46750 13268 46756 13320
rect 46808 13308 46814 13320
rect 47780 13317 47808 13348
rect 47765 13311 47823 13317
rect 46808 13280 46874 13308
rect 46808 13268 46814 13280
rect 47765 13277 47777 13311
rect 47811 13277 47823 13311
rect 47765 13271 47823 13277
rect 47946 13268 47952 13320
rect 48004 13268 48010 13320
rect 48222 13268 48228 13320
rect 48280 13268 48286 13320
rect 48516 13317 48544 13348
rect 48976 13348 49188 13376
rect 48501 13311 48559 13317
rect 48501 13277 48513 13311
rect 48547 13277 48559 13311
rect 48501 13271 48559 13277
rect 44542 13240 44548 13252
rect 41386 13212 42196 13240
rect 44390 13212 44548 13240
rect 44542 13200 44548 13212
rect 44600 13200 44606 13252
rect 45738 13200 45744 13252
rect 45796 13200 45802 13252
rect 47857 13243 47915 13249
rect 47857 13209 47869 13243
rect 47903 13209 47915 13243
rect 47857 13203 47915 13209
rect 48087 13243 48145 13249
rect 48087 13209 48099 13243
rect 48133 13240 48145 13243
rect 48314 13240 48320 13252
rect 48133 13212 48320 13240
rect 48133 13209 48145 13212
rect 48087 13203 48145 13209
rect 38519 13144 38700 13172
rect 38519 13141 38531 13144
rect 38473 13135 38531 13141
rect 39942 13132 39948 13184
rect 40000 13172 40006 13184
rect 41233 13175 41291 13181
rect 41233 13172 41245 13175
rect 40000 13144 41245 13172
rect 40000 13132 40006 13144
rect 41233 13141 41245 13144
rect 41279 13172 41291 13175
rect 42426 13172 42432 13184
rect 41279 13144 42432 13172
rect 41279 13141 41291 13144
rect 41233 13135 41291 13141
rect 42426 13132 42432 13144
rect 42484 13132 42490 13184
rect 47302 13132 47308 13184
rect 47360 13172 47366 13184
rect 47581 13175 47639 13181
rect 47581 13172 47593 13175
rect 47360 13144 47593 13172
rect 47360 13132 47366 13144
rect 47581 13141 47593 13144
rect 47627 13141 47639 13175
rect 47872 13172 47900 13203
rect 48314 13200 48320 13212
rect 48372 13200 48378 13252
rect 48516 13240 48544 13271
rect 48590 13268 48596 13320
rect 48648 13268 48654 13320
rect 48866 13268 48872 13320
rect 48924 13268 48930 13320
rect 48976 13317 49004 13348
rect 48961 13311 49019 13317
rect 48961 13277 48973 13311
rect 49007 13277 49019 13311
rect 48961 13271 49019 13277
rect 49145 13311 49203 13317
rect 49145 13277 49157 13311
rect 49191 13308 49203 13311
rect 49234 13308 49240 13320
rect 49191 13280 49240 13308
rect 49191 13277 49203 13280
rect 49145 13271 49203 13277
rect 49053 13243 49111 13249
rect 49053 13240 49065 13243
rect 48516 13212 49065 13240
rect 49053 13209 49065 13212
rect 49099 13209 49111 13243
rect 49053 13203 49111 13209
rect 48774 13172 48780 13184
rect 47872 13144 48780 13172
rect 47581 13135 47639 13141
rect 48774 13132 48780 13144
rect 48832 13132 48838 13184
rect 48958 13132 48964 13184
rect 49016 13172 49022 13184
rect 49160 13172 49188 13271
rect 49234 13268 49240 13280
rect 49292 13268 49298 13320
rect 49326 13268 49332 13320
rect 49384 13308 49390 13320
rect 49436 13317 49464 13416
rect 50982 13404 50988 13416
rect 51040 13404 51046 13456
rect 51626 13404 51632 13456
rect 51684 13404 51690 13456
rect 50614 13376 50620 13388
rect 49528 13348 50620 13376
rect 49528 13317 49556 13348
rect 50614 13336 50620 13348
rect 50672 13376 50678 13388
rect 50890 13376 50896 13388
rect 50672 13348 50896 13376
rect 50672 13336 50678 13348
rect 50890 13336 50896 13348
rect 50948 13336 50954 13388
rect 51184 13348 51580 13376
rect 51184 13320 51212 13348
rect 51552 13320 51580 13348
rect 49421 13311 49479 13317
rect 49421 13308 49433 13311
rect 49384 13280 49433 13308
rect 49384 13268 49390 13280
rect 49421 13277 49433 13280
rect 49467 13277 49479 13311
rect 49421 13271 49479 13277
rect 49513 13311 49571 13317
rect 49513 13277 49525 13311
rect 49559 13277 49571 13311
rect 49513 13271 49571 13277
rect 49605 13311 49663 13317
rect 49605 13277 49617 13311
rect 49651 13308 49663 13311
rect 50246 13308 50252 13320
rect 49651 13280 50252 13308
rect 49651 13277 49663 13280
rect 49605 13271 49663 13277
rect 49528 13240 49556 13271
rect 49694 13240 49700 13252
rect 49528 13212 49700 13240
rect 49694 13200 49700 13212
rect 49752 13200 49758 13252
rect 50080 13184 50108 13280
rect 50246 13268 50252 13280
rect 50304 13268 50310 13320
rect 51077 13311 51135 13317
rect 51077 13277 51089 13311
rect 51123 13277 51135 13311
rect 51077 13271 51135 13277
rect 51092 13240 51120 13271
rect 51166 13268 51172 13320
rect 51224 13268 51230 13320
rect 51350 13268 51356 13320
rect 51408 13268 51414 13320
rect 51534 13268 51540 13320
rect 51592 13268 51598 13320
rect 51644 13308 51672 13404
rect 51721 13311 51779 13317
rect 51721 13308 51733 13311
rect 51644 13280 51733 13308
rect 51721 13277 51733 13280
rect 51767 13277 51779 13311
rect 51721 13271 51779 13277
rect 51994 13268 52000 13320
rect 52052 13268 52058 13320
rect 51442 13240 51448 13252
rect 51092 13212 51448 13240
rect 51442 13200 51448 13212
rect 51500 13200 51506 13252
rect 51629 13243 51687 13249
rect 51629 13209 51641 13243
rect 51675 13209 51687 13243
rect 52273 13243 52331 13249
rect 52273 13240 52285 13243
rect 51629 13203 51687 13209
rect 51920 13212 52285 13240
rect 49970 13172 49976 13184
rect 49016 13144 49976 13172
rect 49016 13132 49022 13144
rect 49970 13132 49976 13144
rect 50028 13132 50034 13184
rect 50062 13132 50068 13184
rect 50120 13132 50126 13184
rect 51460 13172 51488 13200
rect 51644 13172 51672 13203
rect 51920 13181 51948 13212
rect 52273 13209 52285 13212
rect 52319 13209 52331 13243
rect 53558 13240 53564 13252
rect 53498 13212 53564 13240
rect 52273 13203 52331 13209
rect 53558 13200 53564 13212
rect 53616 13200 53622 13252
rect 51460 13144 51672 13172
rect 51905 13175 51963 13181
rect 51905 13141 51917 13175
rect 51951 13141 51963 13175
rect 51905 13135 51963 13141
rect 53742 13132 53748 13184
rect 53800 13132 53806 13184
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 23566 12928 23572 12980
rect 23624 12968 23630 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 23624 12940 24777 12968
rect 23624 12928 23630 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 25038 12928 25044 12980
rect 25096 12968 25102 12980
rect 26694 12968 26700 12980
rect 25096 12940 26700 12968
rect 25096 12928 25102 12940
rect 26694 12928 26700 12940
rect 26752 12928 26758 12980
rect 30006 12928 30012 12980
rect 30064 12968 30070 12980
rect 30469 12971 30527 12977
rect 30469 12968 30481 12971
rect 30064 12940 30481 12968
rect 30064 12928 30070 12940
rect 30469 12937 30481 12940
rect 30515 12937 30527 12971
rect 30469 12931 30527 12937
rect 30558 12928 30564 12980
rect 30616 12928 30622 12980
rect 30926 12968 30932 12980
rect 30668 12940 30932 12968
rect 23658 12860 23664 12912
rect 23716 12860 23722 12912
rect 24673 12903 24731 12909
rect 24673 12869 24685 12903
rect 24719 12900 24731 12903
rect 29264 12903 29322 12909
rect 24719 12872 25360 12900
rect 24719 12869 24731 12872
rect 24673 12863 24731 12869
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 25133 12835 25191 12841
rect 25133 12832 25145 12835
rect 24912 12804 25145 12832
rect 24912 12792 24918 12804
rect 25133 12801 25145 12804
rect 25179 12801 25191 12835
rect 25133 12795 25191 12801
rect 25332 12832 25360 12872
rect 27540 12872 29040 12900
rect 25593 12835 25651 12841
rect 25593 12832 25605 12835
rect 25332 12804 25605 12832
rect 25332 12776 25360 12804
rect 25593 12801 25605 12804
rect 25639 12832 25651 12835
rect 26513 12835 26571 12841
rect 26513 12832 26525 12835
rect 25639 12804 26525 12832
rect 25639 12801 25651 12804
rect 25593 12795 25651 12801
rect 26513 12801 26525 12804
rect 26559 12801 26571 12835
rect 26513 12795 26571 12801
rect 26789 12835 26847 12841
rect 26789 12801 26801 12835
rect 26835 12832 26847 12835
rect 26973 12835 27031 12841
rect 26973 12832 26985 12835
rect 26835 12804 26985 12832
rect 26835 12801 26847 12804
rect 26789 12795 26847 12801
rect 22370 12724 22376 12776
rect 22428 12764 22434 12776
rect 22649 12767 22707 12773
rect 22649 12764 22661 12767
rect 22428 12736 22661 12764
rect 22428 12724 22434 12736
rect 22649 12733 22661 12736
rect 22695 12733 22707 12767
rect 22649 12727 22707 12733
rect 22925 12767 22983 12773
rect 22925 12733 22937 12767
rect 22971 12764 22983 12767
rect 24486 12764 24492 12776
rect 22971 12736 24492 12764
rect 22971 12733 22983 12736
rect 22925 12727 22983 12733
rect 24486 12724 24492 12736
rect 24544 12724 24550 12776
rect 25222 12724 25228 12776
rect 25280 12724 25286 12776
rect 25314 12724 25320 12776
rect 25372 12724 25378 12776
rect 25409 12767 25467 12773
rect 25409 12733 25421 12767
rect 25455 12733 25467 12767
rect 25409 12727 25467 12733
rect 25424 12696 25452 12727
rect 26896 12708 26924 12804
rect 26973 12801 26985 12804
rect 27019 12801 27031 12835
rect 26973 12795 27031 12801
rect 27062 12792 27068 12844
rect 27120 12832 27126 12844
rect 27540 12841 27568 12872
rect 29012 12844 29040 12872
rect 29264 12869 29276 12903
rect 29310 12900 29322 12903
rect 30576 12900 30604 12928
rect 29310 12872 30604 12900
rect 29310 12869 29322 12872
rect 29264 12863 29322 12869
rect 27798 12841 27804 12844
rect 27525 12835 27583 12841
rect 27525 12832 27537 12835
rect 27120 12804 27537 12832
rect 27120 12792 27126 12804
rect 27525 12801 27537 12804
rect 27571 12801 27583 12835
rect 27792 12832 27804 12841
rect 27759 12804 27804 12832
rect 27525 12795 27583 12801
rect 27792 12795 27804 12804
rect 27798 12792 27804 12795
rect 27856 12792 27862 12844
rect 28994 12792 29000 12844
rect 29052 12792 29058 12844
rect 30668 12841 30696 12940
rect 30926 12928 30932 12940
rect 30984 12928 30990 12980
rect 31202 12928 31208 12980
rect 31260 12968 31266 12980
rect 31260 12940 32168 12968
rect 31260 12928 31266 12940
rect 32030 12900 32036 12912
rect 30852 12872 32036 12900
rect 30653 12835 30711 12841
rect 30653 12801 30665 12835
rect 30699 12801 30711 12835
rect 30653 12795 30711 12801
rect 25498 12696 25504 12708
rect 25424 12668 25504 12696
rect 25498 12656 25504 12668
rect 25556 12696 25562 12708
rect 26878 12696 26884 12708
rect 25556 12668 26884 12696
rect 25556 12656 25562 12668
rect 26878 12656 26884 12668
rect 26936 12656 26942 12708
rect 30377 12699 30435 12705
rect 30377 12665 30389 12699
rect 30423 12696 30435 12699
rect 30466 12696 30472 12708
rect 30423 12668 30472 12696
rect 30423 12665 30435 12668
rect 30377 12659 30435 12665
rect 30466 12656 30472 12668
rect 30524 12696 30530 12708
rect 30852 12705 30880 12872
rect 30929 12835 30987 12841
rect 30929 12801 30941 12835
rect 30975 12801 30987 12835
rect 30929 12795 30987 12801
rect 30944 12764 30972 12795
rect 31110 12792 31116 12844
rect 31168 12792 31174 12844
rect 31220 12841 31248 12872
rect 32030 12860 32036 12872
rect 32088 12860 32094 12912
rect 32140 12841 32168 12940
rect 32398 12928 32404 12980
rect 32456 12928 32462 12980
rect 32858 12928 32864 12980
rect 32916 12968 32922 12980
rect 33962 12968 33968 12980
rect 32916 12940 33968 12968
rect 32916 12928 32922 12940
rect 33962 12928 33968 12940
rect 34020 12928 34026 12980
rect 34054 12928 34060 12980
rect 34112 12928 34118 12980
rect 34146 12928 34152 12980
rect 34204 12968 34210 12980
rect 34204 12940 36216 12968
rect 34204 12928 34210 12940
rect 31205 12835 31263 12841
rect 31205 12801 31217 12835
rect 31251 12801 31263 12835
rect 31205 12795 31263 12801
rect 31757 12835 31815 12841
rect 31757 12801 31769 12835
rect 31803 12801 31815 12835
rect 31757 12795 31815 12801
rect 32125 12835 32183 12841
rect 32125 12801 32137 12835
rect 32171 12801 32183 12835
rect 32416 12832 32444 12928
rect 34422 12900 34428 12912
rect 32876 12872 34428 12900
rect 32876 12841 32904 12872
rect 34422 12860 34428 12872
rect 34480 12860 34486 12912
rect 34606 12860 34612 12912
rect 34664 12909 34670 12912
rect 34664 12903 34693 12909
rect 34681 12869 34693 12903
rect 34664 12863 34693 12869
rect 34664 12860 34670 12863
rect 34790 12860 34796 12912
rect 34848 12860 34854 12912
rect 36188 12900 36216 12940
rect 36262 12928 36268 12980
rect 36320 12928 36326 12980
rect 36372 12940 37596 12968
rect 36372 12900 36400 12940
rect 36188 12872 36400 12900
rect 36446 12860 36452 12912
rect 36504 12900 36510 12912
rect 36633 12903 36691 12909
rect 36633 12900 36645 12903
rect 36504 12872 36645 12900
rect 36504 12860 36510 12872
rect 36633 12869 36645 12872
rect 36679 12869 36691 12903
rect 36633 12863 36691 12869
rect 36814 12860 36820 12912
rect 36872 12909 36878 12912
rect 36872 12903 36901 12909
rect 36889 12869 36901 12903
rect 37568 12900 37596 12940
rect 37642 12928 37648 12980
rect 37700 12928 37706 12980
rect 38654 12928 38660 12980
rect 38712 12968 38718 12980
rect 39025 12971 39083 12977
rect 39025 12968 39037 12971
rect 38712 12940 39037 12968
rect 38712 12928 38718 12940
rect 39025 12937 39037 12940
rect 39071 12937 39083 12971
rect 40218 12968 40224 12980
rect 39025 12931 39083 12937
rect 39868 12940 40224 12968
rect 38473 12903 38531 12909
rect 38473 12900 38485 12903
rect 37568 12872 38485 12900
rect 36872 12863 36901 12869
rect 36872 12860 36878 12863
rect 32861 12835 32919 12841
rect 32861 12832 32873 12835
rect 32416 12804 32873 12832
rect 32125 12795 32183 12801
rect 32861 12801 32873 12804
rect 32907 12801 32919 12835
rect 32861 12795 32919 12801
rect 33045 12835 33103 12841
rect 33045 12801 33057 12835
rect 33091 12832 33103 12835
rect 33870 12832 33876 12844
rect 33091 12804 33876 12832
rect 33091 12801 33103 12804
rect 33045 12795 33103 12801
rect 31386 12764 31392 12776
rect 30944 12736 31392 12764
rect 31386 12724 31392 12736
rect 31444 12724 31450 12776
rect 31481 12767 31539 12773
rect 31481 12733 31493 12767
rect 31527 12764 31539 12767
rect 31573 12767 31631 12773
rect 31573 12764 31585 12767
rect 31527 12736 31585 12764
rect 31527 12733 31539 12736
rect 31481 12727 31539 12733
rect 31573 12733 31585 12736
rect 31619 12764 31631 12767
rect 31662 12764 31668 12776
rect 31619 12736 31668 12764
rect 31619 12733 31631 12736
rect 31573 12727 31631 12733
rect 31662 12724 31668 12736
rect 31720 12724 31726 12776
rect 31772 12764 31800 12795
rect 31938 12764 31944 12776
rect 31772 12736 31944 12764
rect 31938 12724 31944 12736
rect 31996 12764 32002 12776
rect 33060 12764 33088 12795
rect 33870 12792 33876 12804
rect 33928 12792 33934 12844
rect 33962 12792 33968 12844
rect 34020 12832 34026 12844
rect 34333 12835 34391 12841
rect 34333 12832 34345 12835
rect 34020 12804 34345 12832
rect 34020 12792 34026 12804
rect 34333 12801 34345 12804
rect 34379 12801 34391 12835
rect 34333 12795 34391 12801
rect 34517 12835 34575 12841
rect 34517 12801 34529 12835
rect 34563 12832 34575 12835
rect 34808 12832 34836 12860
rect 36541 12835 36599 12841
rect 34563 12804 36492 12832
rect 34563 12801 34575 12804
rect 34517 12795 34575 12801
rect 31996 12736 33088 12764
rect 33505 12767 33563 12773
rect 31996 12724 32002 12736
rect 33505 12733 33517 12767
rect 33551 12764 33563 12767
rect 34149 12767 34207 12773
rect 34149 12764 34161 12767
rect 33551 12736 34161 12764
rect 33551 12733 33563 12736
rect 33505 12727 33563 12733
rect 34149 12733 34161 12736
rect 34195 12733 34207 12767
rect 34793 12767 34851 12773
rect 34793 12764 34805 12767
rect 34149 12727 34207 12733
rect 34532 12736 34805 12764
rect 34532 12708 34560 12736
rect 34793 12733 34805 12736
rect 34839 12733 34851 12767
rect 34793 12727 34851 12733
rect 35713 12767 35771 12773
rect 35713 12733 35725 12767
rect 35759 12764 35771 12767
rect 36357 12767 36415 12773
rect 36357 12764 36369 12767
rect 35759 12736 36369 12764
rect 35759 12733 35771 12736
rect 35713 12727 35771 12733
rect 36357 12733 36369 12736
rect 36403 12733 36415 12767
rect 36357 12727 36415 12733
rect 30745 12699 30803 12705
rect 30745 12696 30757 12699
rect 30524 12668 30757 12696
rect 30524 12656 30530 12668
rect 30745 12665 30757 12668
rect 30791 12665 30803 12699
rect 30745 12659 30803 12665
rect 30837 12699 30895 12705
rect 30837 12665 30849 12699
rect 30883 12665 30895 12699
rect 30837 12659 30895 12665
rect 31297 12699 31355 12705
rect 31297 12665 31309 12699
rect 31343 12696 31355 12699
rect 33778 12696 33784 12708
rect 31343 12668 31616 12696
rect 31343 12665 31355 12668
rect 31297 12659 31355 12665
rect 31588 12640 31616 12668
rect 31956 12668 33784 12696
rect 26234 12588 26240 12640
rect 26292 12588 26298 12640
rect 26326 12588 26332 12640
rect 26384 12588 26390 12640
rect 26694 12588 26700 12640
rect 26752 12628 26758 12640
rect 27065 12631 27123 12637
rect 27065 12628 27077 12631
rect 26752 12600 27077 12628
rect 26752 12588 26758 12600
rect 27065 12597 27077 12600
rect 27111 12597 27123 12631
rect 27065 12591 27123 12597
rect 27430 12588 27436 12640
rect 27488 12588 27494 12640
rect 28905 12631 28963 12637
rect 28905 12597 28917 12631
rect 28951 12628 28963 12631
rect 29270 12628 29276 12640
rect 28951 12600 29276 12628
rect 28951 12597 28963 12600
rect 28905 12591 28963 12597
rect 29270 12588 29276 12600
rect 29328 12588 29334 12640
rect 31570 12588 31576 12640
rect 31628 12588 31634 12640
rect 31956 12637 31984 12668
rect 33778 12656 33784 12668
rect 33836 12656 33842 12708
rect 34514 12656 34520 12708
rect 34572 12656 34578 12708
rect 36464 12696 36492 12804
rect 36541 12801 36553 12835
rect 36587 12801 36599 12835
rect 36541 12795 36599 12801
rect 36556 12764 36584 12795
rect 36722 12792 36728 12844
rect 36780 12792 36786 12844
rect 36998 12792 37004 12844
rect 37056 12792 37062 12844
rect 37274 12792 37280 12844
rect 37332 12792 37338 12844
rect 37458 12792 37464 12844
rect 37516 12792 37522 12844
rect 37553 12835 37611 12841
rect 37553 12801 37565 12835
rect 37599 12801 37611 12835
rect 37553 12795 37611 12801
rect 37568 12764 37596 12795
rect 37826 12792 37832 12844
rect 37884 12792 37890 12844
rect 37918 12792 37924 12844
rect 37976 12832 37982 12844
rect 38120 12841 38148 12872
rect 38473 12869 38485 12872
rect 38519 12900 38531 12903
rect 38519 12872 38654 12900
rect 38519 12869 38531 12872
rect 38473 12863 38531 12869
rect 38105 12835 38163 12841
rect 37976 12804 38056 12832
rect 37976 12792 37982 12804
rect 38028 12764 38056 12804
rect 38105 12801 38117 12835
rect 38151 12801 38163 12835
rect 38105 12795 38163 12801
rect 36556 12736 38056 12764
rect 38626 12764 38654 12872
rect 38746 12860 38752 12912
rect 38804 12900 38810 12912
rect 38841 12903 38899 12909
rect 38841 12900 38853 12903
rect 38804 12872 38853 12900
rect 38804 12860 38810 12872
rect 38841 12869 38853 12872
rect 38887 12900 38899 12903
rect 38887 12872 39160 12900
rect 38887 12869 38899 12872
rect 38841 12863 38899 12869
rect 39132 12841 39160 12872
rect 38933 12835 38991 12841
rect 38933 12801 38945 12835
rect 38979 12801 38991 12835
rect 38933 12795 38991 12801
rect 39117 12835 39175 12841
rect 39117 12801 39129 12835
rect 39163 12801 39175 12835
rect 39117 12795 39175 12801
rect 38948 12764 38976 12795
rect 39206 12792 39212 12844
rect 39264 12792 39270 12844
rect 39868 12841 39896 12940
rect 40218 12928 40224 12940
rect 40276 12928 40282 12980
rect 41046 12928 41052 12980
rect 41104 12928 41110 12980
rect 41233 12971 41291 12977
rect 41233 12937 41245 12971
rect 41279 12968 41291 12971
rect 41279 12940 41414 12968
rect 41279 12937 41291 12940
rect 41233 12931 41291 12937
rect 39942 12860 39948 12912
rect 40000 12860 40006 12912
rect 41386 12900 41414 12940
rect 42334 12928 42340 12980
rect 42392 12968 42398 12980
rect 43809 12971 43867 12977
rect 43809 12968 43821 12971
rect 42392 12940 43821 12968
rect 42392 12928 42398 12940
rect 43809 12937 43821 12940
rect 43855 12937 43867 12971
rect 43809 12931 43867 12937
rect 44542 12928 44548 12980
rect 44600 12928 44606 12980
rect 45557 12971 45615 12977
rect 45557 12937 45569 12971
rect 45603 12968 45615 12971
rect 45738 12968 45744 12980
rect 45603 12940 45744 12968
rect 45603 12937 45615 12940
rect 45557 12931 45615 12937
rect 45738 12928 45744 12940
rect 45796 12928 45802 12980
rect 48222 12928 48228 12980
rect 48280 12968 48286 12980
rect 48777 12971 48835 12977
rect 48777 12968 48789 12971
rect 48280 12940 48789 12968
rect 48280 12928 48286 12940
rect 48777 12937 48789 12940
rect 48823 12937 48835 12971
rect 48777 12931 48835 12937
rect 51350 12928 51356 12980
rect 51408 12968 51414 12980
rect 53377 12971 53435 12977
rect 53377 12968 53389 12971
rect 51408 12940 53389 12968
rect 51408 12928 51414 12940
rect 53377 12937 53389 12940
rect 53423 12937 53435 12971
rect 53377 12931 53435 12937
rect 53558 12928 53564 12980
rect 53616 12928 53622 12980
rect 53742 12928 53748 12980
rect 53800 12928 53806 12980
rect 42674 12903 42732 12909
rect 42674 12900 42686 12903
rect 41386 12872 42686 12900
rect 42674 12869 42686 12872
rect 42720 12869 42732 12903
rect 42674 12863 42732 12869
rect 44174 12860 44180 12912
rect 44232 12900 44238 12912
rect 44910 12900 44916 12912
rect 44232 12872 44916 12900
rect 44232 12860 44238 12872
rect 44910 12860 44916 12872
rect 44968 12860 44974 12912
rect 48406 12860 48412 12912
rect 48464 12900 48470 12912
rect 49053 12903 49111 12909
rect 49053 12900 49065 12903
rect 48464 12872 49065 12900
rect 48464 12860 48470 12872
rect 49053 12869 49065 12872
rect 49099 12869 49111 12903
rect 49053 12863 49111 12869
rect 51626 12860 51632 12912
rect 51684 12900 51690 12912
rect 51905 12903 51963 12909
rect 51905 12900 51917 12903
rect 51684 12872 51917 12900
rect 51684 12860 51690 12872
rect 51905 12869 51917 12872
rect 51951 12869 51963 12903
rect 53760 12900 53788 12928
rect 51905 12863 51963 12869
rect 52012 12872 53788 12900
rect 39853 12835 39911 12841
rect 39853 12801 39865 12835
rect 39899 12801 39911 12835
rect 40034 12832 40040 12844
rect 39853 12795 39911 12801
rect 39960 12804 40040 12832
rect 39224 12764 39252 12792
rect 39960 12764 39988 12804
rect 40034 12792 40040 12804
rect 40092 12792 40098 12844
rect 40126 12792 40132 12844
rect 40184 12841 40190 12844
rect 40184 12835 40213 12841
rect 40201 12801 40213 12835
rect 40184 12795 40213 12801
rect 40313 12835 40371 12841
rect 40313 12801 40325 12835
rect 40359 12832 40371 12835
rect 41230 12832 41236 12844
rect 40359 12804 41236 12832
rect 40359 12801 40371 12804
rect 40313 12795 40371 12801
rect 40184 12792 40190 12795
rect 41230 12792 41236 12804
rect 41288 12792 41294 12844
rect 41417 12835 41475 12841
rect 41417 12801 41429 12835
rect 41463 12832 41475 12835
rect 42150 12832 42156 12844
rect 41463 12804 42156 12832
rect 41463 12801 41475 12804
rect 41417 12795 41475 12801
rect 42150 12792 42156 12804
rect 42208 12792 42214 12844
rect 42242 12792 42248 12844
rect 42300 12832 42306 12844
rect 43901 12835 43959 12841
rect 43901 12832 43913 12835
rect 42300 12804 43913 12832
rect 42300 12792 42306 12804
rect 43901 12801 43913 12804
rect 43947 12801 43959 12835
rect 43901 12795 43959 12801
rect 44453 12835 44511 12841
rect 44453 12801 44465 12835
rect 44499 12832 44511 12835
rect 44726 12832 44732 12844
rect 44499 12804 44732 12832
rect 44499 12801 44511 12804
rect 44453 12795 44511 12801
rect 44726 12792 44732 12804
rect 44784 12792 44790 12844
rect 45741 12835 45799 12841
rect 45741 12801 45753 12835
rect 45787 12832 45799 12835
rect 45830 12832 45836 12844
rect 45787 12804 45836 12832
rect 45787 12801 45799 12804
rect 45741 12795 45799 12801
rect 45830 12792 45836 12804
rect 45888 12792 45894 12844
rect 46017 12835 46075 12841
rect 46017 12801 46029 12835
rect 46063 12832 46075 12835
rect 46474 12832 46480 12844
rect 46063 12804 46480 12832
rect 46063 12801 46075 12804
rect 46017 12795 46075 12801
rect 46474 12792 46480 12804
rect 46532 12792 46538 12844
rect 49142 12792 49148 12844
rect 49200 12832 49206 12844
rect 49605 12835 49663 12841
rect 49605 12832 49617 12835
rect 49200 12804 49617 12832
rect 49200 12792 49206 12804
rect 49605 12801 49617 12804
rect 49651 12801 49663 12835
rect 49605 12795 49663 12801
rect 49789 12835 49847 12841
rect 49789 12801 49801 12835
rect 49835 12801 49847 12835
rect 49789 12795 49847 12801
rect 38626 12736 38884 12764
rect 38948 12736 39252 12764
rect 39592 12736 39988 12764
rect 40405 12767 40463 12773
rect 36722 12696 36728 12708
rect 36464 12668 36728 12696
rect 36722 12656 36728 12668
rect 36780 12656 36786 12708
rect 38654 12696 38660 12708
rect 37200 12668 38660 12696
rect 31941 12631 31999 12637
rect 31941 12597 31953 12631
rect 31987 12597 31999 12631
rect 31941 12591 31999 12597
rect 32766 12588 32772 12640
rect 32824 12588 32830 12640
rect 33226 12588 33232 12640
rect 33284 12588 33290 12640
rect 35894 12588 35900 12640
rect 35952 12628 35958 12640
rect 37200 12628 37228 12668
rect 38654 12656 38660 12668
rect 38712 12656 38718 12708
rect 35952 12600 37228 12628
rect 35952 12588 35958 12600
rect 37274 12588 37280 12640
rect 37332 12588 37338 12640
rect 37921 12631 37979 12637
rect 37921 12597 37933 12631
rect 37967 12628 37979 12631
rect 38286 12628 38292 12640
rect 37967 12600 38292 12628
rect 37967 12597 37979 12600
rect 37921 12591 37979 12597
rect 38286 12588 38292 12600
rect 38344 12588 38350 12640
rect 38856 12628 38884 12736
rect 38930 12656 38936 12708
rect 38988 12696 38994 12708
rect 39592 12696 39620 12736
rect 40405 12733 40417 12767
rect 40451 12733 40463 12767
rect 40405 12727 40463 12733
rect 42429 12767 42487 12773
rect 42429 12733 42441 12767
rect 42475 12733 42487 12767
rect 42429 12727 42487 12733
rect 45925 12767 45983 12773
rect 45925 12733 45937 12767
rect 45971 12764 45983 12767
rect 46382 12764 46388 12776
rect 45971 12736 46388 12764
rect 45971 12733 45983 12736
rect 45925 12727 45983 12733
rect 38988 12668 39620 12696
rect 39669 12699 39727 12705
rect 38988 12656 38994 12668
rect 39669 12665 39681 12699
rect 39715 12696 39727 12699
rect 40420 12696 40448 12727
rect 39715 12668 40448 12696
rect 39715 12665 39727 12668
rect 39669 12659 39727 12665
rect 39758 12628 39764 12640
rect 38856 12600 39764 12628
rect 39758 12588 39764 12600
rect 39816 12628 39822 12640
rect 40770 12628 40776 12640
rect 39816 12600 40776 12628
rect 39816 12588 39822 12600
rect 40770 12588 40776 12600
rect 40828 12588 40834 12640
rect 42444 12628 42472 12727
rect 46382 12724 46388 12736
rect 46440 12724 46446 12776
rect 48222 12724 48228 12776
rect 48280 12764 48286 12776
rect 48958 12764 48964 12776
rect 48280 12736 48964 12764
rect 48280 12724 48286 12736
rect 48958 12724 48964 12736
rect 49016 12724 49022 12776
rect 49326 12724 49332 12776
rect 49384 12724 49390 12776
rect 49421 12767 49479 12773
rect 49421 12733 49433 12767
rect 49467 12764 49479 12767
rect 49694 12764 49700 12776
rect 49467 12736 49700 12764
rect 49467 12733 49479 12736
rect 49421 12727 49479 12733
rect 49694 12724 49700 12736
rect 49752 12724 49758 12776
rect 46106 12696 46112 12708
rect 43364 12668 46112 12696
rect 42794 12628 42800 12640
rect 42444 12600 42800 12628
rect 42794 12588 42800 12600
rect 42852 12628 42858 12640
rect 43364 12628 43392 12668
rect 46106 12656 46112 12668
rect 46164 12656 46170 12708
rect 49804 12696 49832 12795
rect 50062 12792 50068 12844
rect 50120 12832 50126 12844
rect 50522 12832 50528 12844
rect 50120 12804 50528 12832
rect 50120 12792 50126 12804
rect 50522 12792 50528 12804
rect 50580 12792 50586 12844
rect 50890 12792 50896 12844
rect 50948 12832 50954 12844
rect 52012 12832 52040 12872
rect 50948 12804 52040 12832
rect 52089 12835 52147 12841
rect 50948 12792 50954 12804
rect 52089 12801 52101 12835
rect 52135 12832 52147 12835
rect 52178 12832 52184 12844
rect 52135 12804 52184 12832
rect 52135 12801 52147 12804
rect 52089 12795 52147 12801
rect 52178 12792 52184 12804
rect 52236 12792 52242 12844
rect 52840 12841 52868 12872
rect 52825 12835 52883 12841
rect 52825 12801 52837 12835
rect 52871 12801 52883 12835
rect 52825 12795 52883 12801
rect 53466 12792 53472 12844
rect 53524 12792 53530 12844
rect 49970 12724 49976 12776
rect 50028 12724 50034 12776
rect 51258 12724 51264 12776
rect 51316 12724 51322 12776
rect 51534 12724 51540 12776
rect 51592 12764 51598 12776
rect 52273 12767 52331 12773
rect 52273 12764 52285 12767
rect 51592 12736 52285 12764
rect 51592 12724 51598 12736
rect 52273 12733 52285 12736
rect 52319 12733 52331 12767
rect 52273 12727 52331 12733
rect 50433 12699 50491 12705
rect 50433 12696 50445 12699
rect 49804 12668 50445 12696
rect 50433 12665 50445 12668
rect 50479 12665 50491 12699
rect 50433 12659 50491 12665
rect 42852 12600 43392 12628
rect 49513 12631 49571 12637
rect 42852 12588 42858 12600
rect 49513 12597 49525 12631
rect 49559 12628 49571 12631
rect 49602 12628 49608 12640
rect 49559 12600 49608 12628
rect 49559 12597 49571 12600
rect 49513 12591 49571 12597
rect 49602 12588 49608 12600
rect 49660 12588 49666 12640
rect 51810 12588 51816 12640
rect 51868 12588 51874 12640
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 23658 12384 23664 12436
rect 23716 12384 23722 12436
rect 24486 12384 24492 12436
rect 24544 12384 24550 12436
rect 26510 12384 26516 12436
rect 26568 12424 26574 12436
rect 26605 12427 26663 12433
rect 26605 12424 26617 12427
rect 26568 12396 26617 12424
rect 26568 12384 26574 12396
rect 26605 12393 26617 12396
rect 26651 12393 26663 12427
rect 26605 12387 26663 12393
rect 29362 12384 29368 12436
rect 29420 12424 29426 12436
rect 32306 12424 32312 12436
rect 29420 12396 32312 12424
rect 29420 12384 29426 12396
rect 26326 12356 26332 12368
rect 24688 12328 26332 12356
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12220 23627 12223
rect 23842 12220 23848 12232
rect 23615 12192 23848 12220
rect 23615 12189 23627 12192
rect 23569 12183 23627 12189
rect 23584 12096 23612 12183
rect 23842 12180 23848 12192
rect 23900 12180 23906 12232
rect 24688 12229 24716 12328
rect 26326 12316 26332 12328
rect 26384 12356 26390 12368
rect 26384 12328 27016 12356
rect 26384 12316 26390 12328
rect 24946 12248 24952 12300
rect 25004 12248 25010 12300
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12288 25191 12291
rect 26234 12288 26240 12300
rect 25179 12260 26240 12288
rect 25179 12257 25191 12260
rect 25133 12251 25191 12257
rect 26234 12248 26240 12260
rect 26292 12248 26298 12300
rect 26988 12297 27016 12328
rect 26973 12291 27031 12297
rect 26973 12257 26985 12291
rect 27019 12257 27031 12291
rect 26973 12251 27031 12257
rect 29270 12248 29276 12300
rect 29328 12288 29334 12300
rect 29549 12291 29607 12297
rect 29549 12288 29561 12291
rect 29328 12260 29561 12288
rect 29328 12248 29334 12260
rect 29549 12257 29561 12260
rect 29595 12257 29607 12291
rect 29549 12251 29607 12257
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12220 24823 12223
rect 24964 12220 24992 12248
rect 24811 12192 24992 12220
rect 24811 12189 24823 12192
rect 24765 12183 24823 12189
rect 25222 12180 25228 12232
rect 25280 12180 25286 12232
rect 26513 12223 26571 12229
rect 26513 12220 26525 12223
rect 25332 12192 26525 12220
rect 24854 12112 24860 12164
rect 24912 12112 24918 12164
rect 24995 12155 25053 12161
rect 24995 12121 25007 12155
rect 25041 12152 25053 12155
rect 25240 12152 25268 12180
rect 25041 12124 25268 12152
rect 25041 12121 25053 12124
rect 24995 12115 25053 12121
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 25332 12084 25360 12192
rect 26513 12189 26525 12192
rect 26559 12189 26571 12223
rect 26513 12183 26571 12189
rect 27430 12180 27436 12232
rect 27488 12180 27494 12232
rect 29181 12223 29239 12229
rect 29181 12189 29193 12223
rect 29227 12189 29239 12223
rect 29181 12183 29239 12189
rect 29365 12223 29423 12229
rect 29365 12189 29377 12223
rect 29411 12220 29423 12223
rect 29656 12220 29684 12396
rect 32306 12384 32312 12396
rect 32364 12384 32370 12436
rect 32674 12384 32680 12436
rect 32732 12424 32738 12436
rect 32950 12424 32956 12436
rect 32732 12396 32956 12424
rect 32732 12384 32738 12396
rect 32950 12384 32956 12396
rect 33008 12424 33014 12436
rect 34606 12424 34612 12436
rect 33008 12396 34612 12424
rect 33008 12384 33014 12396
rect 34606 12384 34612 12396
rect 34664 12384 34670 12436
rect 37366 12384 37372 12436
rect 37424 12424 37430 12436
rect 38381 12427 38439 12433
rect 38381 12424 38393 12427
rect 37424 12396 38393 12424
rect 37424 12384 37430 12396
rect 38381 12393 38393 12396
rect 38427 12393 38439 12427
rect 38381 12387 38439 12393
rect 38654 12384 38660 12436
rect 38712 12424 38718 12436
rect 38841 12427 38899 12433
rect 38841 12424 38853 12427
rect 38712 12396 38853 12424
rect 38712 12384 38718 12396
rect 38841 12393 38853 12396
rect 38887 12424 38899 12427
rect 47949 12427 48007 12433
rect 38887 12396 39436 12424
rect 38887 12393 38899 12396
rect 38841 12387 38899 12393
rect 31478 12316 31484 12368
rect 31536 12356 31542 12368
rect 31536 12328 33272 12356
rect 31536 12316 31542 12328
rect 30926 12248 30932 12300
rect 30984 12288 30990 12300
rect 31662 12288 31668 12300
rect 30984 12260 31668 12288
rect 30984 12248 30990 12260
rect 31662 12248 31668 12260
rect 31720 12288 31726 12300
rect 32585 12291 32643 12297
rect 31720 12248 31754 12288
rect 32585 12257 32597 12291
rect 32631 12288 32643 12291
rect 33045 12291 33103 12297
rect 33045 12288 33057 12291
rect 32631 12260 33057 12288
rect 32631 12257 32643 12260
rect 32585 12251 32643 12257
rect 33045 12257 33057 12260
rect 33091 12257 33103 12291
rect 33045 12251 33103 12257
rect 33134 12248 33140 12300
rect 33192 12248 33198 12300
rect 33244 12288 33272 12328
rect 36998 12316 37004 12368
rect 37056 12356 37062 12368
rect 38930 12356 38936 12368
rect 37056 12328 38936 12356
rect 37056 12316 37062 12328
rect 38930 12316 38936 12328
rect 38988 12316 38994 12368
rect 39408 12300 39436 12396
rect 47949 12393 47961 12427
rect 47995 12424 48007 12427
rect 48222 12424 48228 12436
rect 47995 12396 48228 12424
rect 47995 12393 48007 12396
rect 47949 12387 48007 12393
rect 48222 12384 48228 12396
rect 48280 12384 48286 12436
rect 51258 12384 51264 12436
rect 51316 12384 51322 12436
rect 51442 12384 51448 12436
rect 51500 12384 51506 12436
rect 40586 12316 40592 12368
rect 40644 12356 40650 12368
rect 40644 12328 41000 12356
rect 40644 12316 40650 12328
rect 37093 12291 37151 12297
rect 33244 12260 33824 12288
rect 29411 12192 29684 12220
rect 29411 12189 29423 12192
rect 29365 12183 29423 12189
rect 28626 12152 28632 12164
rect 27264 12124 28632 12152
rect 27264 12093 27292 12124
rect 28626 12112 28632 12124
rect 28684 12112 28690 12164
rect 29196 12152 29224 12183
rect 30374 12180 30380 12232
rect 30432 12180 30438 12232
rect 30834 12180 30840 12232
rect 30892 12220 30898 12232
rect 31021 12223 31079 12229
rect 31021 12220 31033 12223
rect 30892 12192 31033 12220
rect 30892 12180 30898 12192
rect 31021 12189 31033 12192
rect 31067 12189 31079 12223
rect 31726 12220 31754 12248
rect 32033 12223 32091 12229
rect 32033 12220 32045 12223
rect 31726 12192 32045 12220
rect 31021 12183 31079 12189
rect 32033 12189 32045 12192
rect 32079 12189 32091 12223
rect 32033 12183 32091 12189
rect 30929 12155 30987 12161
rect 30929 12152 30941 12155
rect 29196 12124 30941 12152
rect 30929 12121 30941 12124
rect 30975 12121 30987 12155
rect 32048 12152 32076 12183
rect 32398 12180 32404 12232
rect 32456 12220 32462 12232
rect 32858 12220 32864 12232
rect 32456 12192 32864 12220
rect 32456 12180 32462 12192
rect 32858 12180 32864 12192
rect 32916 12180 32922 12232
rect 32950 12180 32956 12232
rect 33008 12180 33014 12232
rect 33594 12180 33600 12232
rect 33652 12180 33658 12232
rect 33796 12229 33824 12260
rect 37093 12257 37105 12291
rect 37139 12288 37151 12291
rect 37274 12288 37280 12300
rect 37139 12260 37280 12288
rect 37139 12257 37151 12260
rect 37093 12251 37151 12257
rect 37274 12248 37280 12260
rect 37332 12248 37338 12300
rect 37458 12248 37464 12300
rect 37516 12248 37522 12300
rect 39390 12248 39396 12300
rect 39448 12248 39454 12300
rect 40972 12297 41000 12328
rect 40957 12291 41015 12297
rect 40957 12257 40969 12291
rect 41003 12257 41015 12291
rect 40957 12251 41015 12257
rect 43070 12248 43076 12300
rect 43128 12248 43134 12300
rect 46106 12248 46112 12300
rect 46164 12288 46170 12300
rect 46201 12291 46259 12297
rect 46201 12288 46213 12291
rect 46164 12260 46213 12288
rect 46164 12248 46170 12260
rect 46201 12257 46213 12260
rect 46247 12257 46259 12291
rect 46201 12251 46259 12257
rect 46477 12291 46535 12297
rect 46477 12257 46489 12291
rect 46523 12288 46535 12291
rect 47118 12288 47124 12300
rect 46523 12260 47124 12288
rect 46523 12257 46535 12260
rect 46477 12251 46535 12257
rect 47118 12248 47124 12260
rect 47176 12248 47182 12300
rect 50433 12291 50491 12297
rect 50433 12288 50445 12291
rect 49988 12260 50445 12288
rect 33781 12223 33839 12229
rect 33781 12189 33793 12223
rect 33827 12189 33839 12223
rect 33781 12183 33839 12189
rect 34701 12223 34759 12229
rect 34701 12189 34713 12223
rect 34747 12220 34759 12223
rect 34790 12220 34796 12232
rect 34747 12192 34796 12220
rect 34747 12189 34759 12192
rect 34701 12183 34759 12189
rect 32048 12124 32904 12152
rect 30929 12115 30987 12121
rect 32876 12096 32904 12124
rect 23624 12056 25360 12084
rect 27249 12087 27307 12093
rect 23624 12044 23630 12056
rect 27249 12053 27261 12087
rect 27295 12053 27307 12087
rect 27249 12047 27307 12053
rect 27341 12087 27399 12093
rect 27341 12053 27353 12087
rect 27387 12084 27399 12087
rect 27430 12084 27436 12096
rect 27387 12056 27436 12084
rect 27387 12053 27399 12056
rect 27341 12047 27399 12053
rect 27430 12044 27436 12056
rect 27488 12044 27494 12096
rect 29270 12044 29276 12096
rect 29328 12044 29334 12096
rect 30190 12044 30196 12096
rect 30248 12044 30254 12096
rect 31662 12044 31668 12096
rect 31720 12044 31726 12096
rect 32674 12044 32680 12096
rect 32732 12044 32738 12096
rect 32858 12044 32864 12096
rect 32916 12044 32922 12096
rect 33686 12044 33692 12096
rect 33744 12044 33750 12096
rect 33796 12084 33824 12183
rect 34790 12180 34796 12192
rect 34848 12180 34854 12232
rect 36265 12223 36323 12229
rect 36265 12189 36277 12223
rect 36311 12220 36323 12223
rect 37476 12220 37504 12248
rect 49988 12232 50016 12260
rect 50433 12257 50445 12260
rect 50479 12257 50491 12291
rect 50433 12251 50491 12257
rect 50522 12248 50528 12300
rect 50580 12288 50586 12300
rect 51276 12288 51304 12384
rect 50580 12260 51304 12288
rect 50580 12248 50586 12260
rect 51442 12248 51448 12300
rect 51500 12288 51506 12300
rect 51500 12260 51580 12288
rect 51500 12248 51506 12260
rect 36311 12192 37504 12220
rect 36311 12189 36323 12192
rect 36265 12183 36323 12189
rect 34968 12155 35026 12161
rect 34968 12121 34980 12155
rect 35014 12152 35026 12155
rect 35066 12152 35072 12164
rect 35014 12124 35072 12152
rect 35014 12121 35026 12124
rect 34968 12115 35026 12121
rect 35066 12112 35072 12124
rect 35124 12112 35130 12164
rect 35158 12084 35164 12096
rect 33796 12056 35164 12084
rect 35158 12044 35164 12056
rect 35216 12084 35222 12096
rect 35894 12084 35900 12096
rect 35216 12056 35900 12084
rect 35216 12044 35222 12056
rect 35894 12044 35900 12056
rect 35952 12044 35958 12096
rect 36081 12087 36139 12093
rect 36081 12053 36093 12087
rect 36127 12084 36139 12087
rect 36280 12084 36308 12183
rect 37826 12180 37832 12232
rect 37884 12180 37890 12232
rect 38838 12220 38844 12232
rect 38580 12192 38844 12220
rect 36354 12112 36360 12164
rect 36412 12152 36418 12164
rect 37645 12155 37703 12161
rect 37645 12152 37657 12155
rect 36412 12124 37657 12152
rect 36412 12112 36418 12124
rect 37645 12121 37657 12124
rect 37691 12121 37703 12155
rect 37645 12115 37703 12121
rect 38010 12112 38016 12164
rect 38068 12152 38074 12164
rect 38580 12161 38608 12192
rect 38838 12180 38844 12192
rect 38896 12180 38902 12232
rect 38930 12180 38936 12232
rect 38988 12220 38994 12232
rect 39209 12223 39267 12229
rect 39209 12220 39221 12223
rect 38988 12192 39221 12220
rect 38988 12180 38994 12192
rect 39209 12189 39221 12192
rect 39255 12189 39267 12223
rect 39209 12183 39267 12189
rect 40218 12180 40224 12232
rect 40276 12220 40282 12232
rect 40589 12223 40647 12229
rect 40589 12220 40601 12223
rect 40276 12192 40601 12220
rect 40276 12180 40282 12192
rect 40589 12189 40601 12192
rect 40635 12220 40647 12223
rect 40678 12220 40684 12232
rect 40635 12192 40684 12220
rect 40635 12189 40647 12192
rect 40589 12183 40647 12189
rect 40678 12180 40684 12192
rect 40736 12180 40742 12232
rect 40862 12180 40868 12232
rect 40920 12180 40926 12232
rect 41230 12180 41236 12232
rect 41288 12220 41294 12232
rect 41693 12223 41751 12229
rect 41693 12220 41705 12223
rect 41288 12192 41705 12220
rect 41288 12180 41294 12192
rect 41693 12189 41705 12192
rect 41739 12189 41751 12223
rect 41693 12183 41751 12189
rect 42242 12180 42248 12232
rect 42300 12220 42306 12232
rect 42521 12223 42579 12229
rect 42521 12220 42533 12223
rect 42300 12192 42533 12220
rect 42300 12180 42306 12192
rect 42521 12189 42533 12192
rect 42567 12189 42579 12223
rect 42521 12183 42579 12189
rect 44910 12180 44916 12232
rect 44968 12220 44974 12232
rect 45005 12223 45063 12229
rect 45005 12220 45017 12223
rect 44968 12192 45017 12220
rect 44968 12180 44974 12192
rect 45005 12189 45017 12192
rect 45051 12189 45063 12223
rect 45005 12183 45063 12189
rect 49970 12180 49976 12232
rect 50028 12180 50034 12232
rect 51552 12229 51580 12260
rect 50341 12223 50399 12229
rect 50341 12189 50353 12223
rect 50387 12189 50399 12223
rect 50341 12183 50399 12189
rect 50617 12223 50675 12229
rect 50617 12189 50629 12223
rect 50663 12189 50675 12223
rect 50617 12183 50675 12189
rect 51537 12223 51595 12229
rect 51537 12189 51549 12223
rect 51583 12189 51595 12223
rect 51537 12183 51595 12189
rect 38565 12155 38623 12161
rect 38565 12152 38577 12155
rect 38068 12124 38577 12152
rect 38068 12112 38074 12124
rect 38565 12121 38577 12124
rect 38611 12121 38623 12155
rect 38565 12115 38623 12121
rect 40313 12155 40371 12161
rect 40313 12121 40325 12155
rect 40359 12152 40371 12155
rect 42337 12155 42395 12161
rect 42337 12152 42349 12155
rect 40359 12124 42349 12152
rect 40359 12121 40371 12124
rect 40313 12115 40371 12121
rect 42337 12121 42349 12124
rect 42383 12121 42395 12155
rect 42337 12115 42395 12121
rect 42797 12155 42855 12161
rect 42797 12121 42809 12155
rect 42843 12121 42855 12155
rect 42797 12115 42855 12121
rect 36127 12056 36308 12084
rect 36127 12053 36139 12056
rect 36081 12047 36139 12053
rect 36906 12044 36912 12096
rect 36964 12044 36970 12096
rect 38746 12044 38752 12096
rect 38804 12084 38810 12096
rect 39025 12087 39083 12093
rect 39025 12084 39037 12087
rect 38804 12056 39037 12084
rect 38804 12044 38810 12056
rect 39025 12053 39037 12056
rect 39071 12053 39083 12087
rect 40402 12084 40408 12096
rect 40460 12093 40466 12096
rect 40369 12056 40408 12084
rect 39025 12047 39083 12053
rect 40402 12044 40408 12056
rect 40460 12047 40469 12093
rect 40497 12087 40555 12093
rect 40497 12053 40509 12087
rect 40543 12084 40555 12087
rect 40586 12084 40592 12096
rect 40543 12056 40592 12084
rect 40543 12053 40555 12056
rect 40497 12047 40555 12053
rect 40460 12044 40466 12047
rect 40586 12044 40592 12056
rect 40644 12044 40650 12096
rect 40770 12044 40776 12096
rect 40828 12044 40834 12096
rect 41598 12044 41604 12096
rect 41656 12044 41662 12096
rect 42812 12084 42840 12115
rect 43346 12112 43352 12164
rect 43404 12112 43410 12164
rect 45097 12155 45155 12161
rect 45097 12152 45109 12155
rect 44574 12124 45109 12152
rect 45097 12121 45109 12124
rect 45143 12121 45155 12155
rect 45097 12115 45155 12121
rect 47118 12112 47124 12164
rect 47176 12112 47182 12164
rect 49326 12112 49332 12164
rect 49384 12152 49390 12164
rect 50356 12152 50384 12183
rect 49384 12124 50384 12152
rect 50632 12152 50660 12183
rect 50982 12152 50988 12164
rect 50632 12124 50988 12152
rect 49384 12112 49390 12124
rect 50982 12112 50988 12124
rect 51040 12152 51046 12164
rect 51077 12155 51135 12161
rect 51077 12152 51089 12155
rect 51040 12124 51089 12152
rect 51040 12112 51046 12124
rect 51077 12121 51089 12124
rect 51123 12121 51135 12155
rect 52086 12152 52092 12164
rect 51077 12115 51135 12121
rect 51368 12124 52092 12152
rect 44726 12084 44732 12096
rect 42812 12056 44732 12084
rect 44726 12044 44732 12056
rect 44784 12044 44790 12096
rect 44818 12044 44824 12096
rect 44876 12044 44882 12096
rect 50154 12044 50160 12096
rect 50212 12044 50218 12096
rect 50614 12044 50620 12096
rect 50672 12084 50678 12096
rect 51277 12087 51335 12093
rect 51277 12084 51289 12087
rect 50672 12056 51289 12084
rect 50672 12044 50678 12056
rect 51277 12053 51289 12056
rect 51323 12084 51335 12087
rect 51368 12084 51396 12124
rect 52086 12112 52092 12124
rect 52144 12112 52150 12164
rect 51323 12056 51396 12084
rect 51323 12053 51335 12056
rect 51277 12047 51335 12053
rect 51442 12044 51448 12096
rect 51500 12084 51506 12096
rect 51629 12087 51687 12093
rect 51629 12084 51641 12087
rect 51500 12056 51641 12084
rect 51500 12044 51506 12056
rect 51629 12053 51641 12056
rect 51675 12053 51687 12087
rect 51629 12047 51687 12053
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 25774 11840 25780 11892
rect 25832 11880 25838 11892
rect 25961 11883 26019 11889
rect 25961 11880 25973 11883
rect 25832 11852 25973 11880
rect 25832 11840 25838 11852
rect 25961 11849 25973 11852
rect 26007 11849 26019 11883
rect 27154 11880 27160 11892
rect 25961 11843 26019 11849
rect 26252 11852 27160 11880
rect 26252 11821 26280 11852
rect 27154 11840 27160 11852
rect 27212 11880 27218 11892
rect 27341 11883 27399 11889
rect 27341 11880 27353 11883
rect 27212 11852 27353 11880
rect 27212 11840 27218 11852
rect 27341 11849 27353 11852
rect 27387 11849 27399 11883
rect 27341 11843 27399 11849
rect 29270 11840 29276 11892
rect 29328 11840 29334 11892
rect 30374 11840 30380 11892
rect 30432 11880 30438 11892
rect 31027 11883 31085 11889
rect 31027 11880 31039 11883
rect 30432 11852 31039 11880
rect 30432 11840 30438 11852
rect 31027 11849 31039 11852
rect 31073 11849 31085 11883
rect 31027 11843 31085 11849
rect 31113 11883 31171 11889
rect 31113 11849 31125 11883
rect 31159 11880 31171 11883
rect 31662 11880 31668 11892
rect 31159 11852 31668 11880
rect 31159 11849 31171 11852
rect 31113 11843 31171 11849
rect 31662 11840 31668 11852
rect 31720 11840 31726 11892
rect 32306 11840 32312 11892
rect 32364 11840 32370 11892
rect 33686 11840 33692 11892
rect 33744 11840 33750 11892
rect 35066 11840 35072 11892
rect 35124 11880 35130 11892
rect 35161 11883 35219 11889
rect 35161 11880 35173 11883
rect 35124 11852 35173 11880
rect 35124 11840 35130 11852
rect 35161 11849 35173 11852
rect 35207 11849 35219 11883
rect 36354 11880 36360 11892
rect 35161 11843 35219 11849
rect 35268 11852 36360 11880
rect 26237 11815 26295 11821
rect 26237 11781 26249 11815
rect 26283 11781 26295 11815
rect 26237 11775 26295 11781
rect 26329 11815 26387 11821
rect 26329 11781 26341 11815
rect 26375 11781 26387 11815
rect 26329 11775 26387 11781
rect 24765 11747 24823 11753
rect 24765 11713 24777 11747
rect 24811 11744 24823 11747
rect 25682 11744 25688 11756
rect 24811 11716 25688 11744
rect 24811 11713 24823 11716
rect 24765 11707 24823 11713
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 26145 11747 26203 11753
rect 26145 11713 26157 11747
rect 26191 11742 26203 11747
rect 26191 11714 26280 11742
rect 26191 11713 26203 11714
rect 26145 11707 26203 11713
rect 26252 11608 26280 11714
rect 26344 11676 26372 11775
rect 26694 11772 26700 11824
rect 26752 11772 26758 11824
rect 26878 11772 26884 11824
rect 26936 11812 26942 11824
rect 26973 11815 27031 11821
rect 26973 11812 26985 11815
rect 26936 11784 26985 11812
rect 26936 11772 26942 11784
rect 26973 11781 26985 11784
rect 27019 11781 27031 11815
rect 29288 11812 29316 11840
rect 29702 11815 29760 11821
rect 29702 11812 29714 11815
rect 29288 11784 29714 11812
rect 26973 11775 27031 11781
rect 29702 11781 29714 11784
rect 29748 11781 29760 11815
rect 29702 11775 29760 11781
rect 30926 11772 30932 11824
rect 30984 11772 30990 11824
rect 31386 11772 31392 11824
rect 31444 11812 31450 11824
rect 32324 11812 32352 11840
rect 33312 11815 33370 11821
rect 31444 11784 31708 11812
rect 32324 11784 33272 11812
rect 31444 11772 31450 11784
rect 26418 11704 26424 11756
rect 26476 11753 26482 11756
rect 26476 11747 26505 11753
rect 26493 11713 26505 11747
rect 26476 11707 26505 11713
rect 26605 11747 26663 11753
rect 26605 11713 26617 11747
rect 26651 11744 26663 11747
rect 26712 11744 26740 11772
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 26651 11716 27169 11744
rect 26651 11713 26663 11716
rect 26605 11707 26663 11713
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 26476 11704 26482 11707
rect 28074 11704 28080 11756
rect 28132 11704 28138 11756
rect 31202 11704 31208 11756
rect 31260 11704 31266 11756
rect 31297 11747 31355 11753
rect 31297 11713 31309 11747
rect 31343 11713 31355 11747
rect 31297 11707 31355 11713
rect 26344 11648 28948 11676
rect 28920 11608 28948 11648
rect 28994 11636 29000 11688
rect 29052 11676 29058 11688
rect 29457 11679 29515 11685
rect 29457 11676 29469 11679
rect 29052 11648 29469 11676
rect 29052 11636 29058 11648
rect 29457 11645 29469 11648
rect 29503 11645 29515 11679
rect 29457 11639 29515 11645
rect 31312 11608 31340 11707
rect 31478 11704 31484 11756
rect 31536 11704 31542 11756
rect 31680 11753 31708 11784
rect 31573 11747 31631 11753
rect 31573 11713 31585 11747
rect 31619 11713 31631 11747
rect 31573 11707 31631 11713
rect 31665 11747 31723 11753
rect 31665 11713 31677 11747
rect 31711 11713 31723 11747
rect 31665 11707 31723 11713
rect 32401 11747 32459 11753
rect 32401 11713 32413 11747
rect 32447 11744 32459 11747
rect 32674 11744 32680 11756
rect 32447 11716 32680 11744
rect 32447 11713 32459 11716
rect 32401 11707 32459 11713
rect 31588 11676 31616 11707
rect 32674 11704 32680 11716
rect 32732 11704 32738 11756
rect 33244 11744 33272 11784
rect 33312 11781 33324 11815
rect 33358 11812 33370 11815
rect 33704 11812 33732 11840
rect 35268 11812 35296 11852
rect 36354 11840 36360 11852
rect 36412 11840 36418 11892
rect 36906 11840 36912 11892
rect 36964 11840 36970 11892
rect 37734 11880 37740 11892
rect 37016 11852 37740 11880
rect 36924 11812 36952 11840
rect 33358 11784 33732 11812
rect 35084 11784 35296 11812
rect 36004 11784 36952 11812
rect 33358 11781 33370 11784
rect 33312 11775 33370 11781
rect 34606 11744 34612 11756
rect 33244 11716 34612 11744
rect 34606 11704 34612 11716
rect 34664 11704 34670 11756
rect 35084 11753 35112 11784
rect 35069 11747 35127 11753
rect 35069 11713 35081 11747
rect 35115 11713 35127 11747
rect 35069 11707 35127 11713
rect 35158 11704 35164 11756
rect 35216 11744 35222 11756
rect 35253 11747 35311 11753
rect 35253 11744 35265 11747
rect 35216 11716 35265 11744
rect 35216 11704 35222 11716
rect 35253 11713 35265 11716
rect 35299 11713 35311 11747
rect 35253 11707 35311 11713
rect 35621 11747 35679 11753
rect 35621 11713 35633 11747
rect 35667 11744 35679 11747
rect 35802 11744 35808 11756
rect 35667 11716 35808 11744
rect 35667 11713 35679 11716
rect 35621 11707 35679 11713
rect 35802 11704 35808 11716
rect 35860 11704 35866 11756
rect 35897 11747 35955 11753
rect 35897 11713 35909 11747
rect 35943 11744 35955 11747
rect 36004 11744 36032 11784
rect 35943 11716 36032 11744
rect 35943 11713 35955 11716
rect 35897 11707 35955 11713
rect 36078 11704 36084 11756
rect 36136 11704 36142 11756
rect 36265 11747 36323 11753
rect 36265 11713 36277 11747
rect 36311 11744 36323 11747
rect 37016 11744 37044 11852
rect 37734 11840 37740 11852
rect 37792 11840 37798 11892
rect 37826 11840 37832 11892
rect 37884 11880 37890 11892
rect 38657 11883 38715 11889
rect 38657 11880 38669 11883
rect 37884 11852 38669 11880
rect 37884 11840 37890 11852
rect 38657 11849 38669 11852
rect 38703 11849 38715 11883
rect 38657 11843 38715 11849
rect 40221 11883 40279 11889
rect 40221 11849 40233 11883
rect 40267 11849 40279 11883
rect 40221 11843 40279 11849
rect 40236 11812 40264 11843
rect 41598 11840 41604 11892
rect 41656 11840 41662 11892
rect 42150 11840 42156 11892
rect 42208 11840 42214 11892
rect 43346 11840 43352 11892
rect 43404 11880 43410 11892
rect 44177 11883 44235 11889
rect 44177 11880 44189 11883
rect 43404 11852 44189 11880
rect 43404 11840 43410 11852
rect 44177 11849 44189 11852
rect 44223 11849 44235 11883
rect 44177 11843 44235 11849
rect 47118 11840 47124 11892
rect 47176 11840 47182 11892
rect 49326 11840 49332 11892
rect 49384 11840 49390 11892
rect 50154 11880 50160 11892
rect 49804 11852 50160 11880
rect 40586 11812 40592 11824
rect 37292 11784 38884 11812
rect 40236 11784 40592 11812
rect 37292 11753 37320 11784
rect 38856 11756 38884 11784
rect 40586 11772 40592 11784
rect 40644 11812 40650 11824
rect 40644 11784 41092 11812
rect 40644 11772 40650 11784
rect 36311 11716 37044 11744
rect 37277 11747 37335 11753
rect 36311 11713 36323 11716
rect 36265 11707 36323 11713
rect 37277 11713 37289 11747
rect 37323 11713 37335 11747
rect 37277 11707 37335 11713
rect 37544 11747 37602 11753
rect 37544 11713 37556 11747
rect 37590 11744 37602 11747
rect 38746 11744 38752 11756
rect 37590 11716 38752 11744
rect 37590 11713 37602 11716
rect 37544 11707 37602 11713
rect 38746 11704 38752 11716
rect 38804 11704 38810 11756
rect 38838 11704 38844 11756
rect 38896 11704 38902 11756
rect 39114 11753 39120 11756
rect 39108 11707 39120 11753
rect 39114 11704 39120 11707
rect 39172 11704 39178 11756
rect 40402 11704 40408 11756
rect 40460 11704 40466 11756
rect 41064 11753 41092 11784
rect 41049 11747 41107 11753
rect 41049 11713 41061 11747
rect 41095 11713 41107 11747
rect 41616 11744 41644 11840
rect 44726 11772 44732 11824
rect 44784 11812 44790 11824
rect 44784 11784 47072 11812
rect 44784 11772 44790 11784
rect 41785 11747 41843 11753
rect 41785 11744 41797 11747
rect 41616 11716 41797 11744
rect 41049 11707 41107 11713
rect 41785 11713 41797 11716
rect 41831 11713 41843 11747
rect 41785 11707 41843 11713
rect 41969 11747 42027 11753
rect 41969 11713 41981 11747
rect 42015 11713 42027 11747
rect 41969 11707 42027 11713
rect 44361 11747 44419 11753
rect 44361 11713 44373 11747
rect 44407 11744 44419 11747
rect 44450 11744 44456 11756
rect 44407 11716 44456 11744
rect 44407 11713 44419 11716
rect 44361 11707 44419 11713
rect 32214 11676 32220 11688
rect 31588 11648 32220 11676
rect 32214 11636 32220 11648
rect 32272 11636 32278 11688
rect 32582 11636 32588 11688
rect 32640 11676 32646 11688
rect 33042 11676 33048 11688
rect 32640 11648 33048 11676
rect 32640 11636 32646 11648
rect 33042 11636 33048 11648
rect 33100 11636 33106 11688
rect 35437 11679 35495 11685
rect 35437 11645 35449 11679
rect 35483 11676 35495 11679
rect 35483 11648 36032 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 32766 11608 32772 11620
rect 26252 11580 26648 11608
rect 28920 11580 29500 11608
rect 31312 11580 32772 11608
rect 26620 11552 26648 11580
rect 24854 11500 24860 11552
rect 24912 11500 24918 11552
rect 25222 11500 25228 11552
rect 25280 11540 25286 11552
rect 26418 11540 26424 11552
rect 25280 11512 26424 11540
rect 25280 11500 25286 11512
rect 26418 11500 26424 11512
rect 26476 11500 26482 11552
rect 26602 11500 26608 11552
rect 26660 11500 26666 11552
rect 28261 11543 28319 11549
rect 28261 11509 28273 11543
rect 28307 11540 28319 11543
rect 28902 11540 28908 11552
rect 28307 11512 28908 11540
rect 28307 11509 28319 11512
rect 28261 11503 28319 11509
rect 28902 11500 28908 11512
rect 28960 11500 28966 11552
rect 29472 11540 29500 11580
rect 32766 11568 32772 11580
rect 32824 11568 32830 11620
rect 30558 11540 30564 11552
rect 29472 11512 30564 11540
rect 30558 11500 30564 11512
rect 30616 11500 30622 11552
rect 30834 11500 30840 11552
rect 30892 11500 30898 11552
rect 31294 11500 31300 11552
rect 31352 11500 31358 11552
rect 32674 11500 32680 11552
rect 32732 11540 32738 11552
rect 32953 11543 33011 11549
rect 32953 11540 32965 11543
rect 32732 11512 32965 11540
rect 32732 11500 32738 11512
rect 32953 11509 32965 11512
rect 32999 11509 33011 11543
rect 32953 11503 33011 11509
rect 33962 11500 33968 11552
rect 34020 11540 34026 11552
rect 34425 11543 34483 11549
rect 34425 11540 34437 11543
rect 34020 11512 34437 11540
rect 34020 11500 34026 11512
rect 34425 11509 34437 11512
rect 34471 11509 34483 11543
rect 34425 11503 34483 11509
rect 35802 11500 35808 11552
rect 35860 11500 35866 11552
rect 36004 11540 36032 11648
rect 36096 11608 36124 11704
rect 36446 11636 36452 11688
rect 36504 11636 36510 11688
rect 40770 11636 40776 11688
rect 40828 11676 40834 11688
rect 41138 11676 41144 11688
rect 40828 11648 41144 11676
rect 40828 11636 40834 11648
rect 41138 11636 41144 11648
rect 41196 11676 41202 11688
rect 41984 11676 42012 11707
rect 44450 11704 44456 11716
rect 44508 11704 44514 11756
rect 44910 11704 44916 11756
rect 44968 11744 44974 11756
rect 45189 11747 45247 11753
rect 45189 11744 45201 11747
rect 44968 11716 45201 11744
rect 44968 11704 44974 11716
rect 45189 11713 45201 11716
rect 45235 11713 45247 11747
rect 45189 11707 45247 11713
rect 45373 11747 45431 11753
rect 45373 11713 45385 11747
rect 45419 11713 45431 11747
rect 45373 11707 45431 11713
rect 41196 11648 42012 11676
rect 41196 11636 41202 11648
rect 42426 11636 42432 11688
rect 42484 11636 42490 11688
rect 44637 11679 44695 11685
rect 44637 11645 44649 11679
rect 44683 11645 44695 11679
rect 44637 11639 44695 11645
rect 44729 11679 44787 11685
rect 44729 11645 44741 11679
rect 44775 11676 44787 11679
rect 44818 11676 44824 11688
rect 44775 11648 44824 11676
rect 44775 11645 44787 11648
rect 44729 11639 44787 11645
rect 40957 11611 41015 11617
rect 40957 11608 40969 11611
rect 36096 11580 37136 11608
rect 36446 11540 36452 11552
rect 36004 11512 36452 11540
rect 36446 11500 36452 11512
rect 36504 11500 36510 11552
rect 36998 11500 37004 11552
rect 37056 11500 37062 11552
rect 37108 11540 37136 11580
rect 39776 11580 40969 11608
rect 38286 11540 38292 11552
rect 37108 11512 38292 11540
rect 38286 11500 38292 11512
rect 38344 11500 38350 11552
rect 39206 11500 39212 11552
rect 39264 11540 39270 11552
rect 39776 11540 39804 11580
rect 40957 11577 40969 11580
rect 41003 11577 41015 11611
rect 44652 11608 44680 11639
rect 44818 11636 44824 11648
rect 44876 11676 44882 11688
rect 45094 11676 45100 11688
rect 44876 11648 45100 11676
rect 44876 11636 44882 11648
rect 45094 11636 45100 11648
rect 45152 11676 45158 11688
rect 45388 11676 45416 11707
rect 46106 11704 46112 11756
rect 46164 11704 46170 11756
rect 47044 11753 47072 11784
rect 47762 11772 47768 11824
rect 47820 11812 47826 11824
rect 49804 11812 49832 11852
rect 50154 11840 50160 11852
rect 50212 11840 50218 11892
rect 51442 11880 51448 11892
rect 51276 11852 51448 11880
rect 47820 11784 48346 11812
rect 49712 11784 49832 11812
rect 47820 11772 47826 11784
rect 47029 11747 47087 11753
rect 47029 11713 47041 11747
rect 47075 11744 47087 11747
rect 47210 11744 47216 11756
rect 47075 11716 47216 11744
rect 47075 11713 47087 11716
rect 47029 11707 47087 11713
rect 47210 11704 47216 11716
rect 47268 11704 47274 11756
rect 49712 11753 49740 11784
rect 49878 11772 49884 11824
rect 49936 11772 49942 11824
rect 50019 11815 50077 11821
rect 50019 11781 50031 11815
rect 50065 11812 50077 11815
rect 50338 11812 50344 11824
rect 50065 11784 50344 11812
rect 50065 11781 50077 11784
rect 50019 11775 50077 11781
rect 50338 11772 50344 11784
rect 50396 11772 50402 11824
rect 50522 11772 50528 11824
rect 50580 11812 50586 11824
rect 50982 11812 50988 11824
rect 50580 11784 50988 11812
rect 50580 11772 50586 11784
rect 50982 11772 50988 11784
rect 51040 11772 51046 11824
rect 49697 11747 49755 11753
rect 49697 11713 49709 11747
rect 49743 11713 49755 11747
rect 49697 11707 49755 11713
rect 49789 11747 49847 11753
rect 49789 11713 49801 11747
rect 49835 11713 49847 11747
rect 49789 11707 49847 11713
rect 50157 11747 50215 11753
rect 50157 11713 50169 11747
rect 50203 11744 50215 11747
rect 51169 11747 51227 11753
rect 51169 11744 51181 11747
rect 50203 11742 51028 11744
rect 51092 11742 51181 11744
rect 50203 11716 51181 11742
rect 50203 11713 50215 11716
rect 51000 11714 51120 11716
rect 50157 11707 50215 11713
rect 51169 11713 51181 11716
rect 51215 11713 51227 11747
rect 51169 11707 51227 11713
rect 45152 11648 45416 11676
rect 46124 11676 46152 11704
rect 47578 11676 47584 11688
rect 46124 11648 47584 11676
rect 45152 11636 45158 11648
rect 47578 11636 47584 11648
rect 47636 11636 47642 11688
rect 47854 11636 47860 11688
rect 47912 11636 47918 11688
rect 45189 11611 45247 11617
rect 45189 11608 45201 11611
rect 44652 11580 45201 11608
rect 40957 11571 41015 11577
rect 45189 11577 45201 11580
rect 45235 11577 45247 11611
rect 45189 11571 45247 11577
rect 49602 11568 49608 11620
rect 49660 11568 49666 11620
rect 49804 11608 49832 11707
rect 50430 11636 50436 11688
rect 50488 11676 50494 11688
rect 50525 11679 50583 11685
rect 50525 11676 50537 11679
rect 50488 11648 50537 11676
rect 50488 11636 50494 11648
rect 50525 11645 50537 11648
rect 50571 11645 50583 11679
rect 51276 11676 51304 11852
rect 51442 11840 51448 11852
rect 51500 11840 51506 11892
rect 52178 11880 52184 11892
rect 51762 11852 52184 11880
rect 51762 11821 51790 11852
rect 52178 11840 52184 11852
rect 52236 11840 52242 11892
rect 51629 11815 51687 11821
rect 51629 11812 51641 11815
rect 50525 11639 50583 11645
rect 50632 11648 51304 11676
rect 51368 11784 51641 11812
rect 50632 11608 50660 11648
rect 51368 11608 51396 11784
rect 51629 11781 51641 11784
rect 51675 11781 51687 11815
rect 51629 11775 51687 11781
rect 51747 11815 51805 11821
rect 51747 11781 51759 11815
rect 51793 11781 51805 11815
rect 51747 11775 51805 11781
rect 51997 11815 52055 11821
rect 51997 11781 52009 11815
rect 52043 11812 52055 11815
rect 52086 11812 52092 11824
rect 52043 11784 52092 11812
rect 52043 11781 52055 11784
rect 51997 11775 52055 11781
rect 52086 11772 52092 11784
rect 52144 11812 52150 11824
rect 52144 11784 52776 11812
rect 52144 11772 52150 11784
rect 51445 11747 51503 11753
rect 51445 11713 51457 11747
rect 51491 11713 51503 11747
rect 51445 11707 51503 11713
rect 51460 11676 51488 11707
rect 51534 11704 51540 11756
rect 51592 11704 51598 11756
rect 51902 11704 51908 11756
rect 51960 11704 51966 11756
rect 52181 11747 52239 11753
rect 52181 11713 52193 11747
rect 52227 11744 52239 11747
rect 52270 11744 52276 11756
rect 52227 11716 52276 11744
rect 52227 11713 52239 11716
rect 52181 11707 52239 11713
rect 52270 11704 52276 11716
rect 52328 11744 52334 11756
rect 52748 11753 52776 11784
rect 52733 11747 52791 11753
rect 52328 11716 52592 11744
rect 52328 11704 52334 11716
rect 52365 11679 52423 11685
rect 52365 11676 52377 11679
rect 51460 11648 52377 11676
rect 52365 11645 52377 11648
rect 52411 11645 52423 11679
rect 52564 11676 52592 11716
rect 52733 11713 52745 11747
rect 52779 11713 52791 11747
rect 52733 11707 52791 11713
rect 52917 11747 52975 11753
rect 52917 11713 52929 11747
rect 52963 11713 52975 11747
rect 52917 11707 52975 11713
rect 52932 11676 52960 11707
rect 52564 11648 52960 11676
rect 52365 11639 52423 11645
rect 49804 11580 50660 11608
rect 51046 11580 51396 11608
rect 39264 11512 39804 11540
rect 39264 11500 39270 11512
rect 41690 11500 41696 11552
rect 41748 11500 41754 11552
rect 41874 11500 41880 11552
rect 41932 11540 41938 11552
rect 43073 11543 43131 11549
rect 43073 11540 43085 11543
rect 41932 11512 43085 11540
rect 41932 11500 41938 11512
rect 43073 11509 43085 11512
rect 43119 11509 43131 11543
rect 43073 11503 43131 11509
rect 44545 11543 44603 11549
rect 44545 11509 44557 11543
rect 44591 11540 44603 11543
rect 45097 11543 45155 11549
rect 45097 11540 45109 11543
rect 44591 11512 45109 11540
rect 44591 11509 44603 11512
rect 44545 11503 44603 11509
rect 45097 11509 45109 11512
rect 45143 11509 45155 11543
rect 45097 11503 45155 11509
rect 49510 11500 49516 11552
rect 49568 11500 49574 11552
rect 49620 11540 49648 11568
rect 51046 11540 51074 11580
rect 49620 11512 51074 11540
rect 51258 11500 51264 11552
rect 51316 11500 51322 11552
rect 51368 11540 51396 11580
rect 51718 11568 51724 11620
rect 51776 11608 51782 11620
rect 52825 11611 52883 11617
rect 52825 11608 52837 11611
rect 51776 11580 52837 11608
rect 51776 11568 51782 11580
rect 52825 11577 52837 11580
rect 52871 11577 52883 11611
rect 52825 11571 52883 11577
rect 68462 11568 68468 11620
rect 68520 11568 68526 11620
rect 51810 11540 51816 11552
rect 51368 11512 51816 11540
rect 51810 11500 51816 11512
rect 51868 11500 51874 11552
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 26510 11336 26516 11348
rect 26160 11308 26516 11336
rect 22370 11160 22376 11212
rect 22428 11160 22434 11212
rect 22649 11203 22707 11209
rect 22649 11169 22661 11203
rect 22695 11200 22707 11203
rect 24394 11200 24400 11212
rect 22695 11172 24400 11200
rect 22695 11169 22707 11172
rect 22649 11163 22707 11169
rect 24394 11160 24400 11172
rect 24452 11160 24458 11212
rect 25498 11160 25504 11212
rect 25556 11200 25562 11212
rect 25593 11203 25651 11209
rect 25593 11200 25605 11203
rect 25556 11172 25605 11200
rect 25556 11160 25562 11172
rect 25593 11169 25605 11172
rect 25639 11169 25651 11203
rect 25593 11163 25651 11169
rect 25685 11203 25743 11209
rect 25685 11169 25697 11203
rect 25731 11200 25743 11203
rect 25958 11200 25964 11212
rect 25731 11172 25964 11200
rect 25731 11169 25743 11172
rect 25685 11163 25743 11169
rect 25958 11160 25964 11172
rect 26016 11200 26022 11212
rect 26160 11200 26188 11308
rect 26510 11296 26516 11308
rect 26568 11296 26574 11348
rect 26602 11296 26608 11348
rect 26660 11296 26666 11348
rect 27154 11296 27160 11348
rect 27212 11296 27218 11348
rect 27617 11339 27675 11345
rect 27617 11305 27629 11339
rect 27663 11336 27675 11339
rect 28074 11336 28080 11348
rect 27663 11308 28080 11336
rect 27663 11305 27675 11308
rect 27617 11299 27675 11305
rect 28074 11296 28080 11308
rect 28132 11296 28138 11348
rect 28350 11296 28356 11348
rect 28408 11296 28414 11348
rect 28626 11296 28632 11348
rect 28684 11336 28690 11348
rect 28684 11308 30144 11336
rect 28684 11296 28690 11308
rect 26421 11271 26479 11277
rect 26421 11237 26433 11271
rect 26467 11268 26479 11271
rect 28721 11271 28779 11277
rect 26467 11240 28672 11268
rect 26467 11237 26479 11240
rect 26421 11231 26479 11237
rect 26016 11172 26188 11200
rect 26016 11160 26022 11172
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11132 24823 11135
rect 25130 11132 25136 11144
rect 24811 11104 25136 11132
rect 24811 11101 24823 11104
rect 24765 11095 24823 11101
rect 23658 11024 23664 11076
rect 23716 11024 23722 11076
rect 24121 10999 24179 11005
rect 24121 10965 24133 10999
rect 24167 10996 24179 10999
rect 24780 10996 24808 11095
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 25314 11092 25320 11144
rect 25372 11132 25378 11144
rect 25774 11132 25780 11144
rect 25372 11104 25780 11132
rect 25372 11092 25378 11104
rect 25774 11092 25780 11104
rect 25832 11092 25838 11144
rect 25866 11092 25872 11144
rect 25924 11092 25930 11144
rect 26050 11092 26056 11144
rect 26108 11092 26114 11144
rect 26160 11141 26188 11172
rect 26234 11160 26240 11212
rect 26292 11160 26298 11212
rect 26896 11172 27476 11200
rect 26145 11135 26203 11141
rect 26145 11101 26157 11135
rect 26191 11132 26203 11135
rect 26191 11104 26225 11132
rect 26191 11101 26203 11104
rect 26145 11095 26203 11101
rect 26418 11092 26424 11144
rect 26476 11092 26482 11144
rect 26513 11135 26571 11141
rect 26513 11101 26525 11135
rect 26559 11101 26571 11135
rect 26513 11095 26571 11101
rect 26688 11135 26746 11141
rect 26688 11101 26700 11135
rect 26734 11110 26746 11135
rect 26734 11101 26748 11110
rect 26688 11095 26748 11101
rect 25498 11024 25504 11076
rect 25556 11064 25562 11076
rect 26528 11064 26556 11095
rect 26712 11082 26748 11095
rect 25556 11036 26556 11064
rect 26720 11064 26748 11082
rect 26786 11064 26792 11076
rect 26720 11036 26792 11064
rect 25556 11024 25562 11036
rect 26786 11024 26792 11036
rect 26844 11024 26850 11076
rect 24167 10968 24808 10996
rect 24167 10965 24179 10968
rect 24121 10959 24179 10965
rect 25038 10956 25044 11008
rect 25096 10996 25102 11008
rect 25317 10999 25375 11005
rect 25317 10996 25329 10999
rect 25096 10968 25329 10996
rect 25096 10956 25102 10968
rect 25317 10965 25329 10968
rect 25363 10965 25375 10999
rect 25317 10959 25375 10965
rect 25406 10956 25412 11008
rect 25464 10956 25470 11008
rect 25774 10956 25780 11008
rect 25832 10996 25838 11008
rect 26234 10996 26240 11008
rect 25832 10968 26240 10996
rect 25832 10956 25838 10968
rect 26234 10956 26240 10968
rect 26292 10996 26298 11008
rect 26896 10996 26924 11172
rect 27448 11144 27476 11172
rect 27338 11092 27344 11144
rect 27396 11092 27402 11144
rect 27430 11092 27436 11144
rect 27488 11092 27494 11144
rect 27893 11135 27951 11141
rect 27893 11101 27905 11135
rect 27939 11132 27951 11135
rect 28074 11132 28080 11144
rect 27939 11104 28080 11132
rect 27939 11101 27951 11104
rect 27893 11095 27951 11101
rect 28074 11092 28080 11104
rect 28132 11092 28138 11144
rect 28169 11135 28227 11141
rect 28169 11101 28181 11135
rect 28215 11132 28227 11135
rect 28350 11132 28356 11144
rect 28215 11104 28356 11132
rect 28215 11101 28227 11104
rect 28169 11095 28227 11101
rect 28350 11092 28356 11104
rect 28408 11092 28414 11144
rect 28445 11135 28503 11141
rect 28445 11101 28457 11135
rect 28491 11101 28503 11135
rect 28445 11095 28503 11101
rect 27157 11067 27215 11073
rect 27157 11033 27169 11067
rect 27203 11064 27215 11067
rect 27709 11067 27767 11073
rect 27709 11064 27721 11067
rect 27203 11036 27721 11064
rect 27203 11033 27215 11036
rect 27157 11027 27215 11033
rect 27709 11033 27721 11036
rect 27755 11033 27767 11067
rect 28092 11064 28120 11092
rect 28261 11067 28319 11073
rect 28261 11064 28273 11067
rect 28092 11036 28273 11064
rect 27709 11027 27767 11033
rect 28261 11033 28273 11036
rect 28307 11033 28319 11067
rect 28460 11064 28488 11095
rect 28534 11092 28540 11144
rect 28592 11092 28598 11144
rect 28644 11132 28672 11240
rect 28721 11237 28733 11271
rect 28767 11268 28779 11271
rect 30009 11271 30067 11277
rect 30009 11268 30021 11271
rect 28767 11240 30021 11268
rect 28767 11237 28779 11240
rect 28721 11231 28779 11237
rect 30009 11237 30021 11240
rect 30055 11237 30067 11271
rect 30009 11231 30067 11237
rect 30116 11209 30144 11308
rect 30392 11308 32904 11336
rect 29733 11203 29791 11209
rect 29733 11169 29745 11203
rect 29779 11200 29791 11203
rect 30101 11203 30159 11209
rect 29779 11172 30052 11200
rect 29779 11169 29791 11172
rect 29733 11163 29791 11169
rect 30024 11144 30052 11172
rect 30101 11169 30113 11203
rect 30147 11169 30159 11203
rect 30101 11163 30159 11169
rect 30193 11203 30251 11209
rect 30193 11169 30205 11203
rect 30239 11169 30251 11203
rect 30193 11163 30251 11169
rect 29917 11135 29975 11141
rect 29917 11132 29929 11135
rect 28644 11104 29929 11132
rect 29917 11101 29929 11104
rect 29963 11101 29975 11135
rect 29917 11095 29975 11101
rect 30006 11092 30012 11144
rect 30064 11092 30070 11144
rect 30208 11064 30236 11163
rect 30392 11141 30420 11308
rect 30558 11228 30564 11280
rect 30616 11268 30622 11280
rect 31113 11271 31171 11277
rect 31113 11268 31125 11271
rect 30616 11240 31125 11268
rect 30616 11228 30622 11240
rect 31113 11237 31125 11240
rect 31159 11237 31171 11271
rect 31113 11231 31171 11237
rect 32674 11228 32680 11280
rect 32732 11228 32738 11280
rect 30377 11135 30435 11141
rect 30377 11101 30389 11135
rect 30423 11101 30435 11135
rect 30377 11095 30435 11101
rect 30558 11092 30564 11144
rect 30616 11092 30622 11144
rect 31386 11092 31392 11144
rect 31444 11132 31450 11144
rect 31573 11135 31631 11141
rect 31573 11132 31585 11135
rect 31444 11104 31585 11132
rect 31444 11092 31450 11104
rect 31573 11101 31585 11104
rect 31619 11132 31631 11135
rect 32582 11132 32588 11144
rect 31619 11104 32588 11132
rect 31619 11101 31631 11104
rect 31573 11095 31631 11101
rect 32582 11092 32588 11104
rect 32640 11092 32646 11144
rect 30650 11064 30656 11076
rect 28460 11036 30144 11064
rect 30208 11036 30656 11064
rect 28261 11027 28319 11033
rect 26292 10968 26924 10996
rect 28077 10999 28135 11005
rect 26292 10956 26298 10968
rect 28077 10965 28089 10999
rect 28123 10996 28135 10999
rect 28166 10996 28172 11008
rect 28123 10968 28172 10996
rect 28123 10965 28135 10968
rect 28077 10959 28135 10965
rect 28166 10956 28172 10968
rect 28224 10956 28230 11008
rect 30116 10996 30144 11036
rect 30650 11024 30656 11036
rect 30708 11024 30714 11076
rect 30742 11024 30748 11076
rect 30800 11064 30806 11076
rect 31840 11067 31898 11073
rect 30800 11036 31754 11064
rect 30800 11024 30806 11036
rect 30760 10996 30788 11024
rect 30116 10968 30788 10996
rect 31726 10996 31754 11036
rect 31840 11033 31852 11067
rect 31886 11064 31898 11067
rect 32692 11064 32720 11228
rect 32876 11200 32904 11308
rect 35802 11296 35808 11348
rect 35860 11296 35866 11348
rect 35894 11296 35900 11348
rect 35952 11336 35958 11348
rect 36173 11339 36231 11345
rect 36173 11336 36185 11339
rect 35952 11308 36185 11336
rect 35952 11296 35958 11308
rect 36173 11305 36185 11308
rect 36219 11336 36231 11339
rect 38749 11339 38807 11345
rect 36219 11308 38424 11336
rect 36219 11305 36231 11308
rect 36173 11299 36231 11305
rect 35820 11268 35848 11296
rect 35820 11240 38240 11268
rect 38212 11209 38240 11240
rect 38396 11209 38424 11308
rect 38749 11305 38761 11339
rect 38795 11336 38807 11339
rect 38930 11336 38936 11348
rect 38795 11308 38936 11336
rect 38795 11305 38807 11308
rect 38749 11299 38807 11305
rect 38930 11296 38936 11308
rect 38988 11296 38994 11348
rect 39114 11296 39120 11348
rect 39172 11336 39178 11348
rect 39209 11339 39267 11345
rect 39209 11336 39221 11339
rect 39172 11308 39221 11336
rect 39172 11296 39178 11308
rect 39209 11305 39221 11308
rect 39255 11305 39267 11339
rect 39209 11299 39267 11305
rect 39758 11296 39764 11348
rect 39816 11336 39822 11348
rect 39816 11308 40816 11336
rect 39816 11296 39822 11308
rect 40788 11268 40816 11308
rect 41230 11296 41236 11348
rect 41288 11296 41294 11348
rect 45925 11339 45983 11345
rect 45925 11336 45937 11339
rect 41340 11308 45937 11336
rect 41340 11268 41368 11308
rect 45925 11305 45937 11308
rect 45971 11305 45983 11339
rect 45925 11299 45983 11305
rect 47305 11339 47363 11345
rect 47305 11305 47317 11339
rect 47351 11336 47363 11339
rect 47854 11336 47860 11348
rect 47351 11308 47860 11336
rect 47351 11305 47363 11308
rect 47305 11299 47363 11305
rect 47854 11296 47860 11308
rect 47912 11296 47918 11348
rect 49881 11339 49939 11345
rect 49881 11305 49893 11339
rect 49927 11336 49939 11339
rect 50614 11336 50620 11348
rect 49927 11308 50620 11336
rect 49927 11305 49939 11308
rect 49881 11299 49939 11305
rect 50614 11296 50620 11308
rect 50672 11296 50678 11348
rect 50788 11339 50846 11345
rect 50788 11305 50800 11339
rect 50834 11336 50846 11339
rect 51258 11336 51264 11348
rect 50834 11308 51264 11336
rect 50834 11305 50846 11308
rect 50788 11299 50846 11305
rect 51258 11296 51264 11308
rect 51316 11296 51322 11348
rect 51350 11296 51356 11348
rect 51408 11336 51414 11348
rect 51408 11308 52316 11336
rect 51408 11296 51414 11308
rect 40788 11240 41368 11268
rect 46201 11271 46259 11277
rect 46201 11237 46213 11271
rect 46247 11268 46259 11271
rect 47026 11268 47032 11280
rect 46247 11240 47032 11268
rect 46247 11237 46259 11240
rect 46201 11231 46259 11237
rect 47026 11228 47032 11240
rect 47084 11228 47090 11280
rect 47762 11228 47768 11280
rect 47820 11228 47826 11280
rect 47949 11271 48007 11277
rect 47949 11237 47961 11271
rect 47995 11237 48007 11271
rect 47949 11231 48007 11237
rect 36357 11203 36415 11209
rect 32876 11172 34928 11200
rect 34790 11092 34796 11144
rect 34848 11092 34854 11144
rect 34900 11132 34928 11172
rect 36357 11169 36369 11203
rect 36403 11200 36415 11203
rect 37737 11203 37795 11209
rect 37737 11200 37749 11203
rect 36403 11172 37749 11200
rect 36403 11169 36415 11172
rect 36357 11163 36415 11169
rect 37737 11169 37749 11172
rect 37783 11169 37795 11203
rect 37737 11163 37795 11169
rect 38197 11203 38255 11209
rect 38197 11169 38209 11203
rect 38243 11169 38255 11203
rect 38197 11163 38255 11169
rect 38381 11203 38439 11209
rect 38381 11169 38393 11203
rect 38427 11169 38439 11203
rect 38381 11163 38439 11169
rect 38838 11160 38844 11212
rect 38896 11200 38902 11212
rect 39850 11200 39856 11212
rect 38896 11172 39856 11200
rect 38896 11160 38902 11172
rect 39850 11160 39856 11172
rect 39908 11160 39914 11212
rect 41386 11172 41828 11200
rect 37093 11135 37151 11141
rect 34900 11104 37044 11132
rect 31886 11036 32720 11064
rect 35060 11067 35118 11073
rect 31886 11033 31898 11036
rect 31840 11027 31898 11033
rect 35060 11033 35072 11067
rect 35106 11064 35118 11067
rect 36909 11067 36967 11073
rect 36909 11064 36921 11067
rect 35106 11036 36921 11064
rect 35106 11033 35118 11036
rect 35060 11027 35118 11033
rect 36909 11033 36921 11036
rect 36955 11033 36967 11067
rect 37016 11064 37044 11104
rect 37093 11101 37105 11135
rect 37139 11132 37151 11135
rect 37458 11132 37464 11144
rect 37139 11104 37464 11132
rect 37139 11101 37151 11104
rect 37093 11095 37151 11101
rect 37458 11092 37464 11104
rect 37516 11092 37522 11144
rect 37918 11092 37924 11144
rect 37976 11092 37982 11144
rect 38013 11135 38071 11141
rect 38013 11101 38025 11135
rect 38059 11101 38071 11135
rect 38013 11095 38071 11101
rect 37366 11064 37372 11076
rect 37016 11036 37372 11064
rect 36909 11027 36967 11033
rect 37366 11024 37372 11036
rect 37424 11024 37430 11076
rect 38028 11064 38056 11095
rect 38102 11092 38108 11144
rect 38160 11092 38166 11144
rect 38286 11092 38292 11144
rect 38344 11132 38350 11144
rect 38565 11135 38623 11141
rect 38565 11132 38577 11135
rect 38344 11104 38577 11132
rect 38344 11092 38350 11104
rect 38565 11101 38577 11104
rect 38611 11101 38623 11135
rect 38565 11095 38623 11101
rect 39206 11092 39212 11144
rect 39264 11092 39270 11144
rect 39390 11092 39396 11144
rect 39448 11092 39454 11144
rect 39868 11132 39896 11160
rect 41386 11144 41414 11172
rect 41322 11132 41328 11144
rect 39868 11104 41328 11132
rect 41322 11092 41328 11104
rect 41380 11104 41414 11144
rect 41800 11141 41828 11172
rect 45554 11160 45560 11212
rect 45612 11160 45618 11212
rect 46014 11160 46020 11212
rect 46072 11200 46078 11212
rect 46293 11203 46351 11209
rect 46293 11200 46305 11203
rect 46072 11172 46305 11200
rect 46072 11160 46078 11172
rect 46293 11169 46305 11172
rect 46339 11169 46351 11203
rect 47964 11200 47992 11231
rect 52288 11212 52316 11308
rect 46293 11163 46351 11169
rect 47504 11172 47992 11200
rect 41509 11135 41567 11141
rect 41380 11092 41386 11104
rect 41509 11101 41521 11135
rect 41555 11132 41567 11135
rect 41785 11135 41843 11141
rect 41555 11104 41736 11132
rect 41555 11101 41567 11104
rect 41509 11095 41567 11101
rect 41708 11076 41736 11104
rect 41785 11101 41797 11135
rect 41831 11101 41843 11135
rect 45572 11132 45600 11160
rect 46109 11135 46167 11141
rect 46109 11132 46121 11135
rect 45572 11104 46121 11132
rect 41785 11095 41843 11101
rect 46109 11101 46121 11104
rect 46155 11101 46167 11135
rect 46109 11095 46167 11101
rect 46382 11092 46388 11144
rect 46440 11092 46446 11144
rect 47504 11141 47532 11172
rect 48314 11160 48320 11212
rect 48372 11200 48378 11212
rect 48409 11203 48467 11209
rect 48409 11200 48421 11203
rect 48372 11172 48421 11200
rect 48372 11160 48378 11172
rect 48409 11169 48421 11172
rect 48455 11169 48467 11203
rect 48409 11163 48467 11169
rect 48593 11203 48651 11209
rect 48593 11169 48605 11203
rect 48639 11169 48651 11203
rect 48593 11163 48651 11169
rect 49513 11203 49571 11209
rect 49513 11169 49525 11203
rect 49559 11200 49571 11203
rect 49970 11200 49976 11212
rect 49559 11172 49976 11200
rect 49559 11169 49571 11172
rect 49513 11163 49571 11169
rect 46569 11135 46627 11141
rect 46569 11101 46581 11135
rect 46615 11101 46627 11135
rect 46569 11095 46627 11101
rect 47489 11135 47547 11141
rect 47489 11101 47501 11135
rect 47535 11101 47547 11135
rect 47489 11095 47547 11101
rect 47673 11135 47731 11141
rect 47673 11101 47685 11135
rect 47719 11101 47731 11135
rect 48608 11132 48636 11163
rect 49970 11160 49976 11172
rect 50028 11160 50034 11212
rect 51994 11200 52000 11212
rect 50540 11172 52000 11200
rect 49326 11132 49332 11144
rect 48608 11104 49332 11132
rect 47673 11095 47731 11101
rect 40126 11073 40132 11076
rect 37476 11036 38056 11064
rect 32766 10996 32772 11008
rect 31726 10968 32772 10996
rect 32766 10956 32772 10968
rect 32824 10956 32830 11008
rect 32858 10956 32864 11008
rect 32916 10996 32922 11008
rect 32953 10999 33011 11005
rect 32953 10996 32965 10999
rect 32916 10968 32965 10996
rect 32916 10956 32922 10968
rect 32953 10965 32965 10968
rect 32999 10965 33011 10999
rect 32953 10959 33011 10965
rect 37090 10956 37096 11008
rect 37148 10996 37154 11008
rect 37476 10996 37504 11036
rect 40120 11027 40132 11073
rect 40126 11024 40132 11027
rect 40184 11024 40190 11076
rect 41690 11024 41696 11076
rect 41748 11024 41754 11076
rect 42052 11067 42110 11073
rect 42052 11033 42064 11067
rect 42098 11064 42110 11067
rect 43070 11064 43076 11076
rect 42098 11036 43076 11064
rect 42098 11033 42110 11036
rect 42052 11027 42110 11033
rect 43070 11024 43076 11036
rect 43128 11024 43134 11076
rect 45830 11024 45836 11076
rect 45888 11064 45894 11076
rect 46584 11064 46612 11095
rect 45888 11036 46612 11064
rect 45888 11024 45894 11036
rect 47210 11024 47216 11076
rect 47268 11064 47274 11076
rect 47688 11064 47716 11095
rect 49326 11092 49332 11104
rect 49384 11132 49390 11144
rect 50540 11141 50568 11172
rect 51994 11160 52000 11172
rect 52052 11160 52058 11212
rect 52270 11160 52276 11212
rect 52328 11200 52334 11212
rect 52549 11203 52607 11209
rect 52549 11200 52561 11203
rect 52328 11172 52561 11200
rect 52328 11160 52334 11172
rect 52549 11169 52561 11172
rect 52595 11169 52607 11203
rect 52549 11163 52607 11169
rect 49697 11135 49755 11141
rect 49697 11132 49709 11135
rect 49384 11104 49709 11132
rect 49384 11092 49390 11104
rect 49697 11101 49709 11104
rect 49743 11101 49755 11135
rect 50525 11135 50583 11141
rect 50525 11132 50537 11135
rect 49697 11095 49755 11101
rect 49804 11104 50537 11132
rect 47268 11036 47716 11064
rect 48317 11067 48375 11073
rect 47268 11024 47274 11036
rect 48317 11033 48329 11067
rect 48363 11064 48375 11067
rect 49602 11064 49608 11076
rect 48363 11036 49608 11064
rect 48363 11033 48375 11036
rect 48317 11027 48375 11033
rect 49602 11024 49608 11036
rect 49660 11024 49666 11076
rect 37148 10968 37504 10996
rect 37148 10956 37154 10968
rect 37642 10956 37648 11008
rect 37700 10956 37706 11008
rect 41601 10999 41659 11005
rect 41601 10965 41613 10999
rect 41647 10996 41659 10999
rect 42518 10996 42524 11008
rect 41647 10968 42524 10996
rect 41647 10965 41659 10968
rect 41601 10959 41659 10965
rect 42518 10956 42524 10968
rect 42576 10956 42582 11008
rect 43162 10956 43168 11008
rect 43220 10956 43226 11008
rect 49234 10956 49240 11008
rect 49292 10996 49298 11008
rect 49804 10996 49832 11104
rect 50525 11101 50537 11104
rect 50571 11101 50583 11135
rect 50525 11095 50583 11101
rect 51442 11024 51448 11076
rect 51500 11024 51506 11076
rect 49292 10968 49832 10996
rect 49292 10956 49298 10968
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 23569 10795 23627 10801
rect 23569 10761 23581 10795
rect 23615 10792 23627 10795
rect 23658 10792 23664 10804
rect 23615 10764 23664 10792
rect 23615 10761 23627 10764
rect 23569 10755 23627 10761
rect 23658 10752 23664 10764
rect 23716 10752 23722 10804
rect 24394 10752 24400 10804
rect 24452 10752 24458 10804
rect 24854 10752 24860 10804
rect 24912 10752 24918 10804
rect 25314 10752 25320 10804
rect 25372 10752 25378 10804
rect 25498 10752 25504 10804
rect 25556 10752 25562 10804
rect 25682 10752 25688 10804
rect 25740 10752 25746 10804
rect 25869 10795 25927 10801
rect 25869 10761 25881 10795
rect 25915 10792 25927 10795
rect 26418 10792 26424 10804
rect 25915 10764 26424 10792
rect 25915 10761 25927 10764
rect 25869 10755 25927 10761
rect 26418 10752 26424 10764
rect 26476 10752 26482 10804
rect 26786 10752 26792 10804
rect 26844 10752 26850 10804
rect 27338 10752 27344 10804
rect 27396 10752 27402 10804
rect 28442 10792 28448 10804
rect 27540 10764 28448 10792
rect 24673 10727 24731 10733
rect 24673 10693 24685 10727
rect 24719 10724 24731 10727
rect 24872 10724 24900 10752
rect 27540 10736 27568 10764
rect 28442 10752 28448 10764
rect 28500 10792 28506 10804
rect 33594 10792 33600 10804
rect 28500 10764 33600 10792
rect 28500 10752 28506 10764
rect 33594 10752 33600 10764
rect 33652 10792 33658 10804
rect 38562 10792 38568 10804
rect 33652 10764 38568 10792
rect 33652 10752 33658 10764
rect 38562 10752 38568 10764
rect 38620 10792 38626 10804
rect 38620 10764 40816 10792
rect 38620 10752 38626 10764
rect 40788 10736 40816 10764
rect 41138 10752 41144 10804
rect 41196 10792 41202 10804
rect 41196 10764 42012 10792
rect 41196 10752 41202 10764
rect 24719 10696 24900 10724
rect 24719 10693 24731 10696
rect 24673 10687 24731 10693
rect 25222 10684 25228 10736
rect 25280 10684 25286 10736
rect 25409 10727 25467 10733
rect 25409 10693 25421 10727
rect 25455 10724 25467 10727
rect 25958 10724 25964 10736
rect 25455 10696 25964 10724
rect 25455 10693 25467 10696
rect 25409 10687 25467 10693
rect 25958 10684 25964 10696
rect 26016 10684 26022 10736
rect 26050 10684 26056 10736
rect 26108 10724 26114 10736
rect 26326 10724 26332 10736
rect 26108 10696 26332 10724
rect 26108 10684 26114 10696
rect 26326 10684 26332 10696
rect 26384 10724 26390 10736
rect 26384 10696 26924 10724
rect 26384 10684 26390 10696
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10656 23535 10659
rect 23658 10656 23664 10668
rect 23523 10628 23664 10656
rect 23523 10625 23535 10628
rect 23477 10619 23535 10625
rect 23658 10616 23664 10628
rect 23716 10616 23722 10668
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 24627 10628 24716 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 992 10424 1593 10452
rect 992 10412 998 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 24688 10452 24716 10628
rect 24762 10616 24768 10668
rect 24820 10616 24826 10668
rect 24903 10659 24961 10665
rect 24903 10625 24915 10659
rect 24949 10656 24961 10659
rect 25240 10656 25268 10684
rect 24949 10628 25268 10656
rect 24949 10625 24961 10628
rect 24903 10619 24961 10625
rect 25774 10616 25780 10668
rect 25832 10616 25838 10668
rect 25866 10616 25872 10668
rect 25924 10656 25930 10668
rect 26605 10659 26663 10665
rect 25924 10628 26556 10656
rect 25924 10616 25930 10628
rect 25038 10548 25044 10600
rect 25096 10548 25102 10600
rect 25130 10548 25136 10600
rect 25188 10588 25194 10600
rect 25884 10588 25912 10616
rect 25188 10560 25912 10588
rect 26421 10591 26479 10597
rect 25188 10548 25194 10560
rect 26421 10557 26433 10591
rect 26467 10557 26479 10591
rect 26421 10551 26479 10557
rect 25406 10480 25412 10532
rect 25464 10480 25470 10532
rect 26436 10520 26464 10551
rect 25516 10492 26464 10520
rect 25424 10452 25452 10480
rect 25516 10464 25544 10492
rect 24688 10424 25452 10452
rect 1581 10415 1639 10421
rect 25498 10412 25504 10464
rect 25556 10412 25562 10464
rect 26528 10452 26556 10628
rect 26605 10625 26617 10659
rect 26651 10656 26663 10659
rect 26651 10628 26832 10656
rect 26651 10625 26663 10628
rect 26605 10619 26663 10625
rect 26804 10520 26832 10628
rect 26896 10588 26924 10696
rect 27522 10684 27528 10736
rect 27580 10684 27586 10736
rect 28166 10684 28172 10736
rect 28224 10684 28230 10736
rect 28353 10727 28411 10733
rect 28353 10693 28365 10727
rect 28399 10724 28411 10727
rect 28994 10724 29000 10736
rect 28399 10696 29000 10724
rect 28399 10693 28411 10696
rect 28353 10687 28411 10693
rect 28994 10684 29000 10696
rect 29052 10684 29058 10736
rect 29089 10727 29147 10733
rect 29089 10693 29101 10727
rect 29135 10724 29147 10727
rect 30190 10724 30196 10736
rect 29135 10696 30196 10724
rect 29135 10693 29147 10696
rect 29089 10687 29147 10693
rect 30190 10684 30196 10696
rect 30248 10684 30254 10736
rect 33965 10727 34023 10733
rect 33965 10724 33977 10727
rect 33336 10696 33977 10724
rect 26973 10659 27031 10665
rect 26973 10625 26985 10659
rect 27019 10656 27031 10659
rect 28184 10656 28212 10684
rect 27019 10654 27200 10656
rect 27264 10654 28212 10656
rect 27019 10628 28212 10654
rect 27019 10625 27031 10628
rect 27172 10626 27292 10628
rect 26973 10619 27031 10625
rect 28534 10616 28540 10668
rect 28592 10616 28598 10668
rect 29733 10659 29791 10665
rect 29733 10625 29745 10659
rect 29779 10625 29791 10659
rect 29733 10619 29791 10625
rect 27249 10591 27307 10597
rect 27249 10588 27261 10591
rect 26896 10560 27261 10588
rect 27249 10557 27261 10560
rect 27295 10557 27307 10591
rect 27249 10551 27307 10557
rect 27338 10548 27344 10600
rect 27396 10588 27402 10600
rect 28552 10588 28580 10616
rect 28902 10588 28908 10600
rect 27396 10560 28580 10588
rect 28644 10560 28908 10588
rect 27396 10548 27402 10560
rect 28644 10520 28672 10560
rect 28902 10548 28908 10560
rect 28960 10588 28966 10600
rect 29181 10591 29239 10597
rect 29181 10588 29193 10591
rect 28960 10560 29193 10588
rect 28960 10548 28966 10560
rect 29181 10557 29193 10560
rect 29227 10557 29239 10591
rect 29181 10551 29239 10557
rect 29270 10548 29276 10600
rect 29328 10548 29334 10600
rect 26804 10492 28672 10520
rect 28721 10523 28779 10529
rect 28721 10489 28733 10523
rect 28767 10520 28779 10523
rect 29748 10520 29776 10619
rect 33042 10616 33048 10668
rect 33100 10656 33106 10668
rect 33336 10665 33364 10696
rect 33965 10693 33977 10696
rect 34011 10693 34023 10727
rect 36998 10724 37004 10736
rect 33965 10687 34023 10693
rect 35360 10696 37004 10724
rect 33321 10659 33379 10665
rect 33321 10656 33333 10659
rect 33100 10628 33333 10656
rect 33100 10616 33106 10628
rect 33321 10625 33333 10628
rect 33367 10625 33379 10659
rect 33321 10619 33379 10625
rect 33505 10659 33563 10665
rect 33505 10625 33517 10659
rect 33551 10656 33563 10659
rect 34514 10656 34520 10668
rect 33551 10628 34520 10656
rect 33551 10625 33563 10628
rect 33505 10619 33563 10625
rect 30558 10548 30564 10600
rect 30616 10588 30622 10600
rect 32861 10591 32919 10597
rect 32861 10588 32873 10591
rect 30616 10560 32873 10588
rect 30616 10548 30622 10560
rect 32861 10557 32873 10560
rect 32907 10588 32919 10591
rect 33520 10588 33548 10619
rect 34514 10616 34520 10628
rect 34572 10616 34578 10668
rect 35360 10665 35388 10696
rect 36998 10684 37004 10696
rect 37056 10684 37062 10736
rect 38102 10724 38108 10736
rect 37200 10696 38108 10724
rect 35345 10659 35403 10665
rect 35345 10625 35357 10659
rect 35391 10625 35403 10659
rect 36357 10659 36415 10665
rect 35345 10619 35403 10625
rect 35544 10628 36308 10656
rect 32907 10560 33548 10588
rect 32907 10557 32919 10560
rect 32861 10551 32919 10557
rect 34054 10548 34060 10600
rect 34112 10548 34118 10600
rect 34241 10591 34299 10597
rect 34241 10557 34253 10591
rect 34287 10588 34299 10591
rect 35250 10588 35256 10600
rect 34287 10560 35256 10588
rect 34287 10557 34299 10560
rect 34241 10551 34299 10557
rect 28767 10492 29776 10520
rect 28767 10489 28779 10492
rect 28721 10483 28779 10489
rect 32766 10480 32772 10532
rect 32824 10520 32830 10532
rect 34256 10520 34284 10551
rect 35250 10548 35256 10560
rect 35308 10548 35314 10600
rect 35544 10588 35572 10628
rect 35360 10560 35572 10588
rect 35621 10591 35679 10597
rect 32824 10492 34284 10520
rect 32824 10480 32830 10492
rect 35360 10464 35388 10560
rect 35621 10557 35633 10591
rect 35667 10588 35679 10591
rect 35802 10588 35808 10600
rect 35667 10560 35808 10588
rect 35667 10557 35679 10560
rect 35621 10551 35679 10557
rect 35802 10548 35808 10560
rect 35860 10548 35866 10600
rect 36280 10588 36308 10628
rect 36357 10625 36369 10659
rect 36403 10656 36415 10659
rect 37200 10656 37228 10696
rect 38102 10684 38108 10696
rect 38160 10684 38166 10736
rect 40681 10727 40739 10733
rect 40681 10724 40693 10727
rect 40236 10696 40693 10724
rect 36403 10628 37228 10656
rect 36403 10625 36415 10628
rect 36357 10619 36415 10625
rect 37366 10616 37372 10668
rect 37424 10616 37430 10668
rect 37553 10659 37611 10665
rect 37553 10625 37565 10659
rect 37599 10625 37611 10659
rect 37553 10619 37611 10625
rect 37645 10659 37703 10665
rect 37645 10625 37657 10659
rect 37691 10656 37703 10659
rect 37734 10656 37740 10668
rect 37691 10628 37740 10656
rect 37691 10625 37703 10628
rect 37645 10619 37703 10625
rect 36449 10591 36507 10597
rect 36449 10588 36461 10591
rect 36280 10560 36461 10588
rect 36449 10557 36461 10560
rect 36495 10557 36507 10591
rect 37568 10588 37596 10619
rect 37734 10616 37740 10628
rect 37792 10616 37798 10668
rect 37826 10616 37832 10668
rect 37884 10656 37890 10668
rect 40236 10665 40264 10696
rect 40681 10693 40693 10696
rect 40727 10693 40739 10727
rect 40681 10687 40739 10693
rect 40770 10684 40776 10736
rect 40828 10684 40834 10736
rect 37921 10659 37979 10665
rect 37921 10656 37933 10659
rect 37884 10628 37933 10656
rect 37884 10616 37890 10628
rect 37921 10625 37933 10628
rect 37967 10625 37979 10659
rect 37921 10619 37979 10625
rect 40221 10659 40279 10665
rect 40221 10625 40233 10659
rect 40267 10625 40279 10659
rect 40221 10619 40279 10625
rect 40497 10659 40555 10665
rect 40497 10625 40509 10659
rect 40543 10656 40555 10659
rect 41156 10656 41184 10752
rect 41322 10684 41328 10736
rect 41380 10724 41386 10736
rect 41509 10727 41567 10733
rect 41509 10724 41521 10727
rect 41380 10696 41521 10724
rect 41380 10684 41386 10696
rect 41509 10693 41521 10696
rect 41555 10693 41567 10727
rect 41509 10687 41567 10693
rect 41984 10671 42012 10764
rect 43070 10752 43076 10804
rect 43128 10752 43134 10804
rect 44177 10795 44235 10801
rect 44177 10761 44189 10795
rect 44223 10792 44235 10795
rect 44358 10792 44364 10804
rect 44223 10764 44364 10792
rect 44223 10761 44235 10764
rect 44177 10755 44235 10761
rect 44358 10752 44364 10764
rect 44416 10752 44422 10804
rect 44910 10752 44916 10804
rect 44968 10752 44974 10804
rect 45005 10795 45063 10801
rect 45005 10761 45017 10795
rect 45051 10792 45063 10795
rect 45186 10792 45192 10804
rect 45051 10764 45192 10792
rect 45051 10761 45063 10764
rect 45005 10755 45063 10761
rect 45186 10752 45192 10764
rect 45244 10752 45250 10804
rect 50982 10752 50988 10804
rect 51040 10752 51046 10804
rect 51442 10752 51448 10804
rect 51500 10752 51506 10804
rect 44269 10727 44327 10733
rect 44269 10693 44281 10727
rect 44315 10724 44327 10727
rect 44928 10724 44956 10752
rect 44315 10696 44956 10724
rect 44315 10693 44327 10696
rect 44269 10687 44327 10693
rect 49510 10684 49516 10736
rect 49568 10684 49574 10736
rect 51169 10727 51227 10733
rect 51169 10724 51181 10727
rect 50738 10696 51181 10724
rect 51169 10693 51181 10696
rect 51215 10693 51227 10727
rect 51169 10687 51227 10693
rect 40543 10628 41184 10656
rect 40543 10625 40555 10628
rect 40497 10619 40555 10625
rect 41598 10616 41604 10668
rect 41656 10656 41662 10668
rect 41874 10656 41880 10668
rect 41656 10628 41880 10656
rect 41656 10616 41662 10628
rect 41874 10616 41880 10628
rect 41932 10616 41938 10668
rect 41969 10665 42027 10671
rect 41969 10631 41981 10665
rect 42015 10631 42027 10665
rect 41969 10625 42027 10631
rect 47578 10616 47584 10668
rect 47636 10656 47642 10668
rect 49234 10656 49240 10668
rect 47636 10628 49240 10656
rect 47636 10616 47642 10628
rect 49234 10616 49240 10628
rect 49292 10616 49298 10668
rect 51074 10616 51080 10668
rect 51132 10656 51138 10668
rect 51353 10659 51411 10665
rect 51353 10656 51365 10659
rect 51132 10628 51365 10656
rect 51132 10616 51138 10628
rect 51353 10625 51365 10628
rect 51399 10625 51411 10659
rect 51353 10619 51411 10625
rect 39758 10588 39764 10600
rect 37568 10560 39764 10588
rect 36449 10551 36507 10557
rect 39758 10548 39764 10560
rect 39816 10548 39822 10600
rect 40313 10591 40371 10597
rect 40313 10557 40325 10591
rect 40359 10588 40371 10591
rect 41322 10588 41328 10600
rect 40359 10560 41328 10588
rect 40359 10557 40371 10560
rect 40313 10551 40371 10557
rect 41322 10548 41328 10560
rect 41380 10548 41386 10600
rect 42242 10548 42248 10600
rect 42300 10588 42306 10600
rect 42429 10591 42487 10597
rect 42429 10588 42441 10591
rect 42300 10560 42441 10588
rect 42300 10548 42306 10560
rect 42429 10557 42441 10560
rect 42475 10557 42487 10591
rect 42429 10551 42487 10557
rect 44453 10591 44511 10597
rect 44453 10557 44465 10591
rect 44499 10588 44511 10591
rect 44499 10560 45048 10588
rect 44499 10557 44511 10560
rect 44453 10551 44511 10557
rect 35437 10523 35495 10529
rect 35437 10489 35449 10523
rect 35483 10520 35495 10523
rect 37642 10520 37648 10532
rect 35483 10492 37648 10520
rect 35483 10489 35495 10492
rect 35437 10483 35495 10489
rect 37642 10480 37648 10492
rect 37700 10480 37706 10532
rect 37734 10480 37740 10532
rect 37792 10520 37798 10532
rect 38286 10520 38292 10532
rect 37792 10492 38292 10520
rect 37792 10480 37798 10492
rect 38286 10480 38292 10492
rect 38344 10480 38350 10532
rect 40037 10523 40095 10529
rect 40037 10489 40049 10523
rect 40083 10520 40095 10523
rect 40126 10520 40132 10532
rect 40083 10492 40132 10520
rect 40083 10489 40095 10492
rect 40037 10483 40095 10489
rect 40126 10480 40132 10492
rect 40184 10480 40190 10532
rect 45020 10520 45048 10560
rect 45094 10548 45100 10600
rect 45152 10548 45158 10600
rect 45281 10591 45339 10597
rect 45281 10557 45293 10591
rect 45327 10588 45339 10591
rect 45554 10588 45560 10600
rect 45327 10560 45560 10588
rect 45327 10557 45339 10560
rect 45281 10551 45339 10557
rect 45296 10520 45324 10551
rect 45554 10548 45560 10560
rect 45612 10548 45618 10600
rect 45020 10492 45324 10520
rect 27065 10455 27123 10461
rect 27065 10452 27077 10455
rect 26528 10424 27077 10452
rect 27065 10421 27077 10424
rect 27111 10452 27123 10455
rect 28350 10452 28356 10464
rect 27111 10424 28356 10452
rect 27111 10421 27123 10424
rect 27065 10415 27123 10421
rect 28350 10412 28356 10424
rect 28408 10412 28414 10464
rect 29546 10412 29552 10464
rect 29604 10412 29610 10464
rect 33226 10412 33232 10464
rect 33284 10412 33290 10464
rect 33321 10455 33379 10461
rect 33321 10421 33333 10455
rect 33367 10452 33379 10455
rect 33502 10452 33508 10464
rect 33367 10424 33508 10452
rect 33367 10421 33379 10424
rect 33321 10415 33379 10421
rect 33502 10412 33508 10424
rect 33560 10412 33566 10464
rect 33597 10455 33655 10461
rect 33597 10421 33609 10455
rect 33643 10452 33655 10455
rect 33686 10452 33692 10464
rect 33643 10424 33692 10452
rect 33643 10421 33655 10424
rect 33597 10415 33655 10421
rect 33686 10412 33692 10424
rect 33744 10412 33750 10464
rect 35342 10412 35348 10464
rect 35400 10412 35406 10464
rect 36630 10412 36636 10464
rect 36688 10452 36694 10464
rect 37093 10455 37151 10461
rect 37093 10452 37105 10455
rect 36688 10424 37105 10452
rect 36688 10412 36694 10424
rect 37093 10421 37105 10424
rect 37139 10421 37151 10455
rect 37093 10415 37151 10421
rect 37829 10455 37887 10461
rect 37829 10421 37841 10455
rect 37875 10452 37887 10455
rect 38838 10452 38844 10464
rect 37875 10424 38844 10452
rect 37875 10421 37887 10424
rect 37829 10415 37887 10421
rect 38838 10412 38844 10424
rect 38896 10412 38902 10464
rect 42150 10412 42156 10464
rect 42208 10412 42214 10464
rect 43806 10412 43812 10464
rect 43864 10412 43870 10464
rect 44634 10412 44640 10464
rect 44692 10412 44698 10464
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 25685 10251 25743 10257
rect 25685 10217 25697 10251
rect 25731 10248 25743 10251
rect 26418 10248 26424 10260
rect 25731 10220 26424 10248
rect 25731 10217 25743 10220
rect 25685 10211 25743 10217
rect 26418 10208 26424 10220
rect 26476 10208 26482 10260
rect 27338 10248 27344 10260
rect 26528 10220 27344 10248
rect 25869 10183 25927 10189
rect 25869 10180 25881 10183
rect 23952 10152 25881 10180
rect 23952 10053 23980 10152
rect 25869 10149 25881 10152
rect 25915 10149 25927 10183
rect 25869 10143 25927 10149
rect 24673 10115 24731 10121
rect 24673 10081 24685 10115
rect 24719 10112 24731 10115
rect 25774 10112 25780 10124
rect 24719 10084 25780 10112
rect 24719 10081 24731 10084
rect 24673 10075 24731 10081
rect 25774 10072 25780 10084
rect 25832 10072 25838 10124
rect 25884 10084 26188 10112
rect 23937 10047 23995 10053
rect 23937 10013 23949 10047
rect 23983 10013 23995 10047
rect 23937 10007 23995 10013
rect 24213 10047 24271 10053
rect 24213 10013 24225 10047
rect 24259 10013 24271 10047
rect 24213 10007 24271 10013
rect 24228 9976 24256 10007
rect 25590 10004 25596 10056
rect 25648 10044 25654 10056
rect 25884 10044 25912 10084
rect 25648 10016 25912 10044
rect 25961 10047 26019 10053
rect 25648 10004 25654 10016
rect 25961 10013 25973 10047
rect 26007 10044 26019 10047
rect 26050 10044 26056 10056
rect 26007 10016 26056 10044
rect 26007 10013 26019 10016
rect 25961 10007 26019 10013
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 26160 10053 26188 10084
rect 26145 10047 26203 10053
rect 26145 10013 26157 10047
rect 26191 10044 26203 10047
rect 26528 10044 26556 10220
rect 27338 10208 27344 10220
rect 27396 10208 27402 10260
rect 32907 10251 32965 10257
rect 32907 10217 32919 10251
rect 32953 10248 32965 10251
rect 33042 10248 33048 10260
rect 32953 10220 33048 10248
rect 32953 10217 32965 10220
rect 32907 10211 32965 10217
rect 33042 10208 33048 10220
rect 33100 10208 33106 10260
rect 33226 10208 33232 10260
rect 33284 10248 33290 10260
rect 33413 10251 33471 10257
rect 33413 10248 33425 10251
rect 33284 10220 33425 10248
rect 33284 10208 33290 10220
rect 33413 10217 33425 10220
rect 33459 10217 33471 10251
rect 33413 10211 33471 10217
rect 34054 10208 34060 10260
rect 34112 10248 34118 10260
rect 38657 10251 38715 10257
rect 38657 10248 38669 10251
rect 34112 10220 38669 10248
rect 34112 10208 34118 10220
rect 38657 10217 38669 10220
rect 38703 10217 38715 10251
rect 38657 10211 38715 10217
rect 42061 10251 42119 10257
rect 42061 10217 42073 10251
rect 42107 10248 42119 10251
rect 42242 10248 42248 10260
rect 42107 10220 42248 10248
rect 42107 10217 42119 10220
rect 42061 10211 42119 10217
rect 42242 10208 42248 10220
rect 42300 10208 42306 10260
rect 43162 10248 43168 10260
rect 42352 10220 43168 10248
rect 26786 10140 26792 10192
rect 26844 10140 26850 10192
rect 29270 10180 29276 10192
rect 26988 10152 29276 10180
rect 26191 10016 26556 10044
rect 26697 10047 26755 10053
rect 26191 10013 26203 10016
rect 26145 10007 26203 10013
rect 26697 10013 26709 10047
rect 26743 10044 26755 10047
rect 26804 10044 26832 10140
rect 26988 10121 27016 10152
rect 29270 10140 29276 10152
rect 29328 10180 29334 10192
rect 34701 10183 34759 10189
rect 29328 10152 30420 10180
rect 29328 10140 29334 10152
rect 30392 10121 30420 10152
rect 34701 10149 34713 10183
rect 34747 10180 34759 10183
rect 35618 10180 35624 10192
rect 34747 10152 35624 10180
rect 34747 10149 34759 10152
rect 34701 10143 34759 10149
rect 35618 10140 35624 10152
rect 35676 10140 35682 10192
rect 40586 10180 40592 10192
rect 38212 10152 40592 10180
rect 26973 10115 27031 10121
rect 26973 10081 26985 10115
rect 27019 10081 27031 10115
rect 30377 10115 30435 10121
rect 26973 10075 27031 10081
rect 27080 10084 28764 10112
rect 26743 10016 26832 10044
rect 26743 10013 26755 10016
rect 26697 10007 26755 10013
rect 26878 10004 26884 10056
rect 26936 10004 26942 10056
rect 24854 9976 24860 9988
rect 24228 9948 24860 9976
rect 24854 9936 24860 9948
rect 24912 9936 24918 9988
rect 25498 9936 25504 9988
rect 25556 9976 25562 9988
rect 27080 9976 27108 10084
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10044 27215 10047
rect 27203 10016 27476 10044
rect 27203 10013 27215 10016
rect 27157 10007 27215 10013
rect 25556 9948 27108 9976
rect 25556 9936 25562 9948
rect 27448 9920 27476 10016
rect 27522 10004 27528 10056
rect 27580 10004 27586 10056
rect 28736 10053 28764 10084
rect 30377 10081 30389 10115
rect 30423 10112 30435 10115
rect 30742 10112 30748 10124
rect 30423 10084 30748 10112
rect 30423 10081 30435 10084
rect 30377 10075 30435 10081
rect 30742 10072 30748 10084
rect 30800 10072 30806 10124
rect 30926 10072 30932 10124
rect 30984 10112 30990 10124
rect 31481 10115 31539 10121
rect 31481 10112 31493 10115
rect 30984 10084 31493 10112
rect 30984 10072 30990 10084
rect 31481 10081 31493 10084
rect 31527 10081 31539 10115
rect 34333 10115 34391 10121
rect 34333 10112 34345 10115
rect 31481 10075 31539 10081
rect 32784 10084 34345 10112
rect 32784 10056 32812 10084
rect 34333 10081 34345 10084
rect 34379 10081 34391 10115
rect 34333 10075 34391 10081
rect 35345 10115 35403 10121
rect 35345 10081 35357 10115
rect 35391 10112 35403 10115
rect 35434 10112 35440 10124
rect 35391 10084 35440 10112
rect 35391 10081 35403 10084
rect 35345 10075 35403 10081
rect 28537 10047 28595 10053
rect 28537 10013 28549 10047
rect 28583 10013 28595 10047
rect 28537 10007 28595 10013
rect 28721 10047 28779 10053
rect 28721 10013 28733 10047
rect 28767 10044 28779 10047
rect 30558 10044 30564 10056
rect 28767 10016 30564 10044
rect 28767 10013 28779 10016
rect 28721 10007 28779 10013
rect 28258 9936 28264 9988
rect 28316 9936 28322 9988
rect 28552 9976 28580 10007
rect 30558 10004 30564 10016
rect 30616 10004 30622 10056
rect 31113 10047 31171 10053
rect 31113 10013 31125 10047
rect 31159 10044 31171 10047
rect 31386 10044 31392 10056
rect 31159 10016 31392 10044
rect 31159 10013 31171 10016
rect 31113 10007 31171 10013
rect 31386 10004 31392 10016
rect 31444 10004 31450 10056
rect 32766 10004 32772 10056
rect 32824 10004 32830 10056
rect 33229 10047 33287 10053
rect 33229 10013 33241 10047
rect 33275 10013 33287 10047
rect 33229 10007 33287 10013
rect 28902 9976 28908 9988
rect 28552 9948 28908 9976
rect 28902 9936 28908 9948
rect 28960 9976 28966 9988
rect 28960 9948 31156 9976
rect 28960 9936 28966 9948
rect 31128 9920 31156 9948
rect 32214 9936 32220 9988
rect 32272 9936 32278 9988
rect 33244 9976 33272 10007
rect 33502 10004 33508 10056
rect 33560 10004 33566 10056
rect 33594 10004 33600 10056
rect 33652 10004 33658 10056
rect 34348 10044 34376 10075
rect 35434 10072 35440 10084
rect 35492 10072 35498 10124
rect 34790 10044 34796 10056
rect 34348 10016 34796 10044
rect 34790 10004 34796 10016
rect 34848 10044 34854 10056
rect 35805 10047 35863 10053
rect 35805 10044 35817 10047
rect 34848 10016 35817 10044
rect 34848 10004 34854 10016
rect 35805 10013 35817 10016
rect 35851 10013 35863 10047
rect 35805 10007 35863 10013
rect 37277 10047 37335 10053
rect 37277 10013 37289 10047
rect 37323 10044 37335 10047
rect 37642 10044 37648 10056
rect 37323 10016 37648 10044
rect 37323 10013 37335 10016
rect 37277 10007 37335 10013
rect 37642 10004 37648 10016
rect 37700 10004 37706 10056
rect 38212 10053 38240 10152
rect 40586 10140 40592 10152
rect 40644 10140 40650 10192
rect 42352 10189 42380 10220
rect 43162 10208 43168 10220
rect 43220 10248 43226 10260
rect 44775 10251 44833 10257
rect 43220 10220 44128 10248
rect 43220 10208 43226 10220
rect 42337 10183 42395 10189
rect 40880 10152 42288 10180
rect 38286 10072 38292 10124
rect 38344 10112 38350 10124
rect 38381 10115 38439 10121
rect 38381 10112 38393 10115
rect 38344 10084 38393 10112
rect 38344 10072 38350 10084
rect 38381 10081 38393 10084
rect 38427 10112 38439 10115
rect 39022 10112 39028 10124
rect 38427 10084 39028 10112
rect 38427 10081 38439 10084
rect 38381 10075 38439 10081
rect 39022 10072 39028 10084
rect 39080 10112 39086 10124
rect 39209 10115 39267 10121
rect 39209 10112 39221 10115
rect 39080 10084 39221 10112
rect 39080 10072 39086 10084
rect 39209 10081 39221 10084
rect 39255 10081 39267 10115
rect 39209 10075 39267 10081
rect 40034 10072 40040 10124
rect 40092 10112 40098 10124
rect 40880 10112 40908 10152
rect 40092 10084 40908 10112
rect 40092 10072 40098 10084
rect 38197 10047 38255 10053
rect 38197 10013 38209 10047
rect 38243 10013 38255 10047
rect 39574 10044 39580 10056
rect 38197 10007 38255 10013
rect 38948 10016 39580 10044
rect 32784 9948 33272 9976
rect 23474 9868 23480 9920
rect 23532 9908 23538 9920
rect 23753 9911 23811 9917
rect 23753 9908 23765 9911
rect 23532 9880 23765 9908
rect 23532 9868 23538 9880
rect 23753 9877 23765 9880
rect 23799 9877 23811 9911
rect 23753 9871 23811 9877
rect 24121 9911 24179 9917
rect 24121 9877 24133 9911
rect 24167 9908 24179 9911
rect 25225 9911 25283 9917
rect 25225 9908 25237 9911
rect 24167 9880 25237 9908
rect 24167 9877 24179 9880
rect 24121 9871 24179 9877
rect 25225 9877 25237 9880
rect 25271 9877 25283 9911
rect 25225 9871 25283 9877
rect 25682 9868 25688 9920
rect 25740 9917 25746 9920
rect 25740 9911 25759 9917
rect 25747 9877 25759 9911
rect 25740 9871 25759 9877
rect 26053 9911 26111 9917
rect 26053 9877 26065 9911
rect 26099 9908 26111 9911
rect 26142 9908 26148 9920
rect 26099 9880 26148 9908
rect 26099 9877 26111 9880
rect 26053 9871 26111 9877
rect 25740 9868 25746 9871
rect 26142 9868 26148 9880
rect 26200 9868 26206 9920
rect 26510 9868 26516 9920
rect 26568 9908 26574 9920
rect 27341 9911 27399 9917
rect 27341 9908 27353 9911
rect 26568 9880 27353 9908
rect 26568 9868 26574 9880
rect 27341 9877 27353 9880
rect 27387 9877 27399 9911
rect 27341 9871 27399 9877
rect 27430 9868 27436 9920
rect 27488 9908 27494 9920
rect 28629 9911 28687 9917
rect 28629 9908 28641 9911
rect 27488 9880 28641 9908
rect 27488 9868 27494 9880
rect 28629 9877 28641 9880
rect 28675 9877 28687 9911
rect 28629 9871 28687 9877
rect 31018 9868 31024 9920
rect 31076 9868 31082 9920
rect 31110 9868 31116 9920
rect 31168 9908 31174 9920
rect 32784 9908 32812 9948
rect 34514 9936 34520 9988
rect 34572 9976 34578 9988
rect 35069 9979 35127 9985
rect 35069 9976 35081 9979
rect 34572 9948 35081 9976
rect 34572 9936 34578 9948
rect 35069 9945 35081 9948
rect 35115 9945 35127 9979
rect 35069 9939 35127 9945
rect 36072 9979 36130 9985
rect 36072 9945 36084 9979
rect 36118 9976 36130 9979
rect 36722 9976 36728 9988
rect 36118 9948 36728 9976
rect 36118 9945 36130 9948
rect 36072 9939 36130 9945
rect 36722 9936 36728 9948
rect 36780 9936 36786 9988
rect 36832 9948 37872 9976
rect 31168 9880 32812 9908
rect 31168 9868 31174 9880
rect 33042 9868 33048 9920
rect 33100 9868 33106 9920
rect 35161 9911 35219 9917
rect 35161 9877 35173 9911
rect 35207 9908 35219 9911
rect 36832 9908 36860 9948
rect 35207 9880 36860 9908
rect 35207 9877 35219 9880
rect 35161 9871 35219 9877
rect 37182 9868 37188 9920
rect 37240 9868 37246 9920
rect 37366 9868 37372 9920
rect 37424 9868 37430 9920
rect 37844 9917 37872 9948
rect 38948 9920 38976 10016
rect 39574 10004 39580 10016
rect 39632 10004 39638 10056
rect 40678 10004 40684 10056
rect 40736 10044 40742 10056
rect 40880 10053 40908 10084
rect 41049 10115 41107 10121
rect 41049 10081 41061 10115
rect 41095 10112 41107 10115
rect 42058 10112 42064 10124
rect 41095 10084 42064 10112
rect 41095 10081 41107 10084
rect 41049 10075 41107 10081
rect 42058 10072 42064 10084
rect 42116 10072 42122 10124
rect 42260 10112 42288 10152
rect 42337 10149 42349 10183
rect 42383 10149 42395 10183
rect 42337 10143 42395 10149
rect 42426 10140 42432 10192
rect 42484 10140 42490 10192
rect 44100 10180 44128 10220
rect 44775 10217 44787 10251
rect 44821 10248 44833 10251
rect 44910 10248 44916 10260
rect 44821 10220 44916 10248
rect 44821 10217 44833 10220
rect 44775 10211 44833 10217
rect 44910 10208 44916 10220
rect 44968 10208 44974 10260
rect 45554 10208 45560 10260
rect 45612 10208 45618 10260
rect 46109 10251 46167 10257
rect 46109 10217 46121 10251
rect 46155 10217 46167 10251
rect 46109 10211 46167 10217
rect 46293 10251 46351 10257
rect 46293 10217 46305 10251
rect 46339 10248 46351 10251
rect 46382 10248 46388 10260
rect 46339 10220 46388 10248
rect 46339 10217 46351 10220
rect 46293 10211 46351 10217
rect 45572 10180 45600 10208
rect 46124 10180 46152 10211
rect 46382 10208 46388 10220
rect 46440 10208 46446 10260
rect 44100 10152 45232 10180
rect 45572 10152 45692 10180
rect 46124 10152 46520 10180
rect 42260 10084 42748 10112
rect 40773 10047 40831 10053
rect 40773 10044 40785 10047
rect 40736 10016 40785 10044
rect 40736 10004 40742 10016
rect 40773 10013 40785 10016
rect 40819 10013 40831 10047
rect 40773 10007 40831 10013
rect 40865 10047 40923 10053
rect 40865 10013 40877 10047
rect 40911 10013 40923 10047
rect 40865 10007 40923 10013
rect 40957 10047 41015 10053
rect 40957 10013 40969 10047
rect 41003 10013 41015 10047
rect 40957 10007 41015 10013
rect 40972 9976 41000 10007
rect 41322 10004 41328 10056
rect 41380 10004 41386 10056
rect 42242 10004 42248 10056
rect 42300 10004 42306 10056
rect 42518 10004 42524 10056
rect 42576 10004 42582 10056
rect 42720 10053 42748 10084
rect 42794 10072 42800 10124
rect 42852 10112 42858 10124
rect 42981 10115 43039 10121
rect 42981 10112 42993 10115
rect 42852 10084 42993 10112
rect 42852 10072 42858 10084
rect 42981 10081 42993 10084
rect 43027 10081 43039 10115
rect 43806 10112 43812 10124
rect 42981 10075 43039 10081
rect 43088 10084 43812 10112
rect 42705 10047 42763 10053
rect 42705 10013 42717 10047
rect 42751 10013 42763 10047
rect 42705 10007 42763 10013
rect 41969 9979 42027 9985
rect 41969 9976 41981 9979
rect 39040 9948 40724 9976
rect 40972 9948 41981 9976
rect 37829 9911 37887 9917
rect 37829 9877 37841 9911
rect 37875 9877 37887 9911
rect 37829 9871 37887 9877
rect 38289 9911 38347 9917
rect 38289 9877 38301 9911
rect 38335 9908 38347 9911
rect 38930 9908 38936 9920
rect 38335 9880 38936 9908
rect 38335 9877 38347 9880
rect 38289 9871 38347 9877
rect 38930 9868 38936 9880
rect 38988 9868 38994 9920
rect 39040 9917 39068 9948
rect 39025 9911 39083 9917
rect 39025 9877 39037 9911
rect 39071 9877 39083 9911
rect 39025 9871 39083 9877
rect 39114 9868 39120 9920
rect 39172 9868 39178 9920
rect 40586 9868 40592 9920
rect 40644 9868 40650 9920
rect 40696 9908 40724 9948
rect 41969 9945 41981 9948
rect 42015 9945 42027 9979
rect 41969 9939 42027 9945
rect 43088 9908 43116 10084
rect 43806 10072 43812 10084
rect 43864 10072 43870 10124
rect 43346 10004 43352 10056
rect 43404 10004 43410 10056
rect 45204 10053 45232 10152
rect 45281 10115 45339 10121
rect 45281 10081 45293 10115
rect 45327 10081 45339 10115
rect 45281 10075 45339 10081
rect 45189 10047 45247 10053
rect 45189 10013 45201 10047
rect 45235 10013 45247 10047
rect 45189 10007 45247 10013
rect 43898 9936 43904 9988
rect 43956 9936 43962 9988
rect 40696 9880 43116 9908
rect 45296 9908 45324 10075
rect 45554 10072 45560 10124
rect 45612 10072 45618 10124
rect 45664 10053 45692 10152
rect 45925 10115 45983 10121
rect 45925 10081 45937 10115
rect 45971 10112 45983 10115
rect 45971 10081 45984 10112
rect 45925 10075 45984 10081
rect 45649 10047 45707 10053
rect 45649 10013 45661 10047
rect 45695 10013 45707 10047
rect 45649 10007 45707 10013
rect 45956 9920 45984 10075
rect 46014 10004 46020 10056
rect 46072 10044 46078 10056
rect 46109 10047 46167 10053
rect 46109 10044 46121 10047
rect 46072 10016 46121 10044
rect 46072 10004 46078 10016
rect 46109 10013 46121 10016
rect 46155 10013 46167 10047
rect 46109 10007 46167 10013
rect 46492 9920 46520 10152
rect 47578 10072 47584 10124
rect 47636 10112 47642 10124
rect 47765 10115 47823 10121
rect 47765 10112 47777 10115
rect 47636 10084 47777 10112
rect 47636 10072 47642 10084
rect 47765 10081 47777 10084
rect 47811 10081 47823 10115
rect 47765 10075 47823 10081
rect 48225 10047 48283 10053
rect 48225 10013 48237 10047
rect 48271 10044 48283 10047
rect 50154 10044 50160 10056
rect 48271 10016 50160 10044
rect 48271 10013 48283 10016
rect 48225 10007 48283 10013
rect 50154 10004 50160 10016
rect 50212 10004 50218 10056
rect 46934 9936 46940 9988
rect 46992 9976 46998 9988
rect 47029 9979 47087 9985
rect 47029 9976 47041 9979
rect 46992 9948 47041 9976
rect 46992 9936 46998 9948
rect 47029 9945 47041 9948
rect 47075 9945 47087 9979
rect 47029 9939 47087 9945
rect 48038 9936 48044 9988
rect 48096 9936 48102 9988
rect 45922 9908 45928 9920
rect 45296 9880 45928 9908
rect 45922 9868 45928 9880
rect 45980 9868 45986 9920
rect 46474 9868 46480 9920
rect 46532 9908 46538 9920
rect 48409 9911 48467 9917
rect 48409 9908 48421 9911
rect 46532 9880 48421 9908
rect 46532 9868 46538 9880
rect 48409 9877 48421 9880
rect 48455 9877 48467 9911
rect 48409 9871 48467 9877
rect 50062 9868 50068 9920
rect 50120 9908 50126 9920
rect 50801 9911 50859 9917
rect 50801 9908 50813 9911
rect 50120 9880 50813 9908
rect 50120 9868 50126 9880
rect 50801 9877 50813 9880
rect 50847 9877 50859 9911
rect 50801 9871 50859 9877
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 24762 9704 24768 9716
rect 24504 9676 24768 9704
rect 23566 9596 23572 9648
rect 23624 9596 23630 9648
rect 24504 9577 24532 9676
rect 24762 9664 24768 9676
rect 24820 9664 24826 9716
rect 26142 9704 26148 9716
rect 25332 9676 26148 9704
rect 24673 9639 24731 9645
rect 24673 9605 24685 9639
rect 24719 9636 24731 9639
rect 25332 9636 25360 9676
rect 26142 9664 26148 9676
rect 26200 9664 26206 9716
rect 26326 9664 26332 9716
rect 26384 9664 26390 9716
rect 30742 9664 30748 9716
rect 30800 9664 30806 9716
rect 30926 9664 30932 9716
rect 30984 9664 30990 9716
rect 31018 9664 31024 9716
rect 31076 9664 31082 9716
rect 31386 9664 31392 9716
rect 31444 9704 31450 9716
rect 31444 9676 31754 9704
rect 31444 9664 31450 9676
rect 24719 9608 25360 9636
rect 24719 9605 24731 9608
rect 24673 9599 24731 9605
rect 25682 9596 25688 9648
rect 25740 9596 25746 9648
rect 25774 9596 25780 9648
rect 25832 9636 25838 9648
rect 25885 9639 25943 9645
rect 25885 9636 25897 9639
rect 25832 9608 25897 9636
rect 25832 9596 25838 9608
rect 25885 9605 25897 9608
rect 25931 9605 25943 9639
rect 25885 9599 25943 9605
rect 26050 9596 26056 9648
rect 26108 9636 26114 9648
rect 26237 9639 26295 9645
rect 26237 9636 26249 9639
rect 26108 9608 26249 9636
rect 26108 9596 26114 9608
rect 26237 9605 26249 9608
rect 26283 9605 26295 9639
rect 26237 9599 26295 9605
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9537 24547 9571
rect 24489 9531 24547 9537
rect 22557 9503 22615 9509
rect 22557 9469 22569 9503
rect 22603 9469 22615 9503
rect 22557 9463 22615 9469
rect 22833 9503 22891 9509
rect 22833 9469 22845 9503
rect 22879 9500 22891 9503
rect 23474 9500 23480 9512
rect 22879 9472 23480 9500
rect 22879 9469 22891 9472
rect 22833 9463 22891 9469
rect 22572 9364 22600 9463
rect 23474 9460 23480 9472
rect 23532 9460 23538 9512
rect 24504 9500 24532 9531
rect 24762 9528 24768 9580
rect 24820 9528 24826 9580
rect 24854 9528 24860 9580
rect 24912 9568 24918 9580
rect 25133 9571 25191 9577
rect 25133 9568 25145 9571
rect 24912 9540 25145 9568
rect 24912 9528 24918 9540
rect 25133 9537 25145 9540
rect 25179 9537 25191 9571
rect 25133 9531 25191 9537
rect 25222 9528 25228 9580
rect 25280 9568 25286 9580
rect 25317 9571 25375 9577
rect 25317 9568 25329 9571
rect 25280 9540 25329 9568
rect 25280 9528 25286 9540
rect 25317 9537 25329 9540
rect 25363 9537 25375 9571
rect 25317 9531 25375 9537
rect 25501 9571 25559 9577
rect 25501 9537 25513 9571
rect 25547 9537 25559 9571
rect 25501 9531 25559 9537
rect 25593 9571 25651 9577
rect 25593 9537 25605 9571
rect 25639 9568 25651 9571
rect 26068 9568 26096 9596
rect 26344 9577 26372 9664
rect 26602 9596 26608 9648
rect 26660 9636 26666 9648
rect 29273 9639 29331 9645
rect 26660 9608 27292 9636
rect 26660 9596 26666 9608
rect 25639 9540 26096 9568
rect 26145 9571 26203 9577
rect 25639 9537 25651 9540
rect 25593 9531 25651 9537
rect 26145 9537 26157 9571
rect 26191 9537 26203 9571
rect 26145 9531 26203 9537
rect 26329 9571 26387 9577
rect 26329 9537 26341 9571
rect 26375 9537 26387 9571
rect 26329 9531 26387 9537
rect 26513 9571 26571 9577
rect 26513 9537 26525 9571
rect 26559 9537 26571 9571
rect 26513 9531 26571 9537
rect 26697 9571 26755 9577
rect 26697 9537 26709 9571
rect 26743 9568 26755 9571
rect 26970 9568 26976 9580
rect 26743 9540 26976 9568
rect 26743 9537 26755 9540
rect 26697 9531 26755 9537
rect 24670 9500 24676 9512
rect 24504 9472 24676 9500
rect 24670 9460 24676 9472
rect 24728 9500 24734 9512
rect 25516 9500 25544 9531
rect 24728 9472 25544 9500
rect 24728 9460 24734 9472
rect 25774 9460 25780 9512
rect 25832 9500 25838 9512
rect 26160 9500 26188 9531
rect 25832 9472 26188 9500
rect 25832 9460 25838 9472
rect 25041 9435 25099 9441
rect 25041 9432 25053 9435
rect 23860 9404 25053 9432
rect 23198 9364 23204 9376
rect 22572 9336 23204 9364
rect 23198 9324 23204 9336
rect 23256 9324 23262 9376
rect 23474 9324 23480 9376
rect 23532 9364 23538 9376
rect 23860 9364 23888 9404
rect 25041 9401 25053 9404
rect 25087 9401 25099 9435
rect 25041 9395 25099 9401
rect 26050 9392 26056 9444
rect 26108 9432 26114 9444
rect 26528 9432 26556 9531
rect 26970 9528 26976 9540
rect 27028 9528 27034 9580
rect 27264 9577 27292 9608
rect 29273 9605 29285 9639
rect 29319 9636 29331 9639
rect 29546 9636 29552 9648
rect 29319 9608 29552 9636
rect 29319 9605 29331 9608
rect 29273 9599 29331 9605
rect 29546 9596 29552 9608
rect 29604 9596 29610 9648
rect 27249 9571 27307 9577
rect 27249 9537 27261 9571
rect 27295 9537 27307 9571
rect 27249 9531 27307 9537
rect 27430 9528 27436 9580
rect 27488 9528 27494 9580
rect 27893 9571 27951 9577
rect 27893 9568 27905 9571
rect 27540 9540 27905 9568
rect 26786 9460 26792 9512
rect 26844 9500 26850 9512
rect 27540 9500 27568 9540
rect 27893 9537 27905 9540
rect 27939 9537 27951 9571
rect 30837 9571 30895 9577
rect 27893 9531 27951 9537
rect 26844 9472 27568 9500
rect 26844 9460 26850 9472
rect 27614 9460 27620 9512
rect 27672 9500 27678 9512
rect 28258 9500 28264 9512
rect 27672 9472 28264 9500
rect 27672 9460 27678 9472
rect 28258 9460 28264 9472
rect 28316 9500 28322 9512
rect 28997 9503 29055 9509
rect 28997 9500 29009 9503
rect 28316 9472 29009 9500
rect 28316 9460 28322 9472
rect 28997 9469 29009 9472
rect 29043 9469 29055 9503
rect 30392 9500 30420 9554
rect 30837 9537 30849 9571
rect 30883 9568 30895 9571
rect 30926 9568 30932 9580
rect 30883 9540 30932 9568
rect 30883 9537 30895 9540
rect 30837 9531 30895 9537
rect 30926 9528 30932 9540
rect 30984 9528 30990 9580
rect 31036 9577 31064 9664
rect 31726 9636 31754 9676
rect 34514 9664 34520 9716
rect 34572 9664 34578 9716
rect 35802 9704 35808 9716
rect 35544 9676 35808 9704
rect 32674 9636 32680 9648
rect 31726 9608 32680 9636
rect 32674 9596 32680 9608
rect 32732 9596 32738 9648
rect 33042 9596 33048 9648
rect 33100 9596 33106 9648
rect 34422 9636 34428 9648
rect 34270 9608 34428 9636
rect 34422 9596 34428 9608
rect 34480 9596 34486 9648
rect 35544 9645 35572 9676
rect 35802 9664 35808 9676
rect 35860 9664 35866 9716
rect 36722 9664 36728 9716
rect 36780 9664 36786 9716
rect 38672 9676 39252 9704
rect 35526 9639 35584 9645
rect 35526 9605 35538 9639
rect 35572 9605 35584 9639
rect 35526 9599 35584 9605
rect 35636 9608 36952 9636
rect 31021 9571 31079 9577
rect 31021 9537 31033 9571
rect 31067 9537 31079 9571
rect 31021 9531 31079 9537
rect 31113 9571 31171 9577
rect 31113 9537 31125 9571
rect 31159 9568 31171 9571
rect 32125 9571 32183 9577
rect 31159 9540 31321 9568
rect 31159 9537 31171 9540
rect 31113 9531 31171 9537
rect 31205 9503 31263 9509
rect 31205 9500 31217 9503
rect 30392 9472 31217 9500
rect 28997 9463 29055 9469
rect 31205 9469 31217 9472
rect 31251 9469 31263 9503
rect 31205 9463 31263 9469
rect 26108 9404 26556 9432
rect 26108 9392 26114 9404
rect 23532 9336 23888 9364
rect 24305 9367 24363 9373
rect 23532 9324 23538 9336
rect 24305 9333 24317 9367
rect 24351 9364 24363 9367
rect 25869 9367 25927 9373
rect 25869 9364 25881 9367
rect 24351 9336 25881 9364
rect 24351 9333 24363 9336
rect 24305 9327 24363 9333
rect 25869 9333 25881 9336
rect 25915 9364 25927 9367
rect 26326 9364 26332 9376
rect 25915 9336 26332 9364
rect 25915 9333 25927 9336
rect 25869 9327 25927 9333
rect 26326 9324 26332 9336
rect 26384 9324 26390 9376
rect 27246 9324 27252 9376
rect 27304 9324 27310 9376
rect 27706 9324 27712 9376
rect 27764 9324 27770 9376
rect 30006 9324 30012 9376
rect 30064 9364 30070 9376
rect 31293 9364 31321 9540
rect 32125 9537 32137 9571
rect 32171 9537 32183 9571
rect 32125 9531 32183 9537
rect 31570 9460 31576 9512
rect 31628 9500 31634 9512
rect 32127 9500 32155 9531
rect 32214 9528 32220 9580
rect 32272 9528 32278 9580
rect 32490 9528 32496 9580
rect 32548 9528 32554 9580
rect 32508 9500 32536 9528
rect 31628 9472 32536 9500
rect 32692 9500 32720 9596
rect 34701 9571 34759 9577
rect 34701 9537 34713 9571
rect 34747 9568 34759 9571
rect 35636 9568 35664 9608
rect 34747 9566 35480 9568
rect 35544 9566 35664 9568
rect 34747 9540 35664 9566
rect 34747 9537 34759 9540
rect 35452 9538 35572 9540
rect 34701 9531 34759 9537
rect 35710 9528 35716 9580
rect 35768 9528 35774 9580
rect 35805 9574 35863 9577
rect 35894 9574 35900 9580
rect 35805 9571 35900 9574
rect 35805 9537 35817 9571
rect 35851 9546 35900 9571
rect 35851 9537 35863 9546
rect 35805 9531 35863 9537
rect 35894 9528 35900 9546
rect 35952 9528 35958 9580
rect 36924 9568 36952 9608
rect 37918 9596 37924 9648
rect 37976 9636 37982 9648
rect 38672 9636 38700 9676
rect 37976 9608 38700 9636
rect 38764 9608 39160 9636
rect 37976 9596 37982 9608
rect 38010 9568 38016 9580
rect 36924 9540 38016 9568
rect 38010 9528 38016 9540
rect 38068 9528 38074 9580
rect 38764 9577 38792 9608
rect 39132 9580 39160 9608
rect 38749 9571 38807 9577
rect 38749 9537 38761 9571
rect 38795 9537 38807 9571
rect 38749 9531 38807 9537
rect 38930 9528 38936 9580
rect 38988 9528 38994 9580
rect 39114 9528 39120 9580
rect 39172 9528 39178 9580
rect 39224 9577 39252 9676
rect 43346 9664 43352 9716
rect 43404 9664 43410 9716
rect 43898 9664 43904 9716
rect 43956 9664 43962 9716
rect 46014 9664 46020 9716
rect 46072 9704 46078 9716
rect 46072 9676 46888 9704
rect 46072 9664 46078 9676
rect 40488 9639 40546 9645
rect 39316 9608 39804 9636
rect 39316 9580 39344 9608
rect 39209 9571 39267 9577
rect 39209 9537 39221 9571
rect 39255 9537 39267 9571
rect 39209 9531 39267 9537
rect 39298 9528 39304 9580
rect 39356 9528 39362 9580
rect 39574 9528 39580 9580
rect 39632 9528 39638 9580
rect 39776 9577 39804 9608
rect 40488 9605 40500 9639
rect 40534 9636 40546 9639
rect 40586 9636 40592 9648
rect 40534 9608 40592 9636
rect 40534 9605 40546 9608
rect 40488 9599 40546 9605
rect 40586 9596 40592 9608
rect 40644 9596 40650 9648
rect 43916 9636 43944 9664
rect 43993 9639 44051 9645
rect 43993 9636 44005 9639
rect 41386 9608 43852 9636
rect 43916 9608 44005 9636
rect 39761 9571 39819 9577
rect 39761 9537 39773 9571
rect 39807 9537 39819 9571
rect 39761 9531 39819 9537
rect 32769 9503 32827 9509
rect 32769 9500 32781 9503
rect 32692 9472 32781 9500
rect 31628 9460 31634 9472
rect 32769 9469 32781 9472
rect 32815 9469 32827 9503
rect 32769 9463 32827 9469
rect 34977 9503 35035 9509
rect 34977 9469 34989 9503
rect 35023 9469 35035 9503
rect 34977 9463 35035 9469
rect 34790 9392 34796 9444
rect 34848 9432 34854 9444
rect 34992 9432 35020 9463
rect 36078 9460 36084 9512
rect 36136 9460 36142 9512
rect 38194 9460 38200 9512
rect 38252 9460 38258 9512
rect 38841 9503 38899 9509
rect 38841 9469 38853 9503
rect 38887 9500 38899 9503
rect 39485 9503 39543 9509
rect 39485 9500 39497 9503
rect 38887 9472 39497 9500
rect 38887 9469 38899 9472
rect 38841 9463 38899 9469
rect 39485 9469 39497 9472
rect 39531 9469 39543 9503
rect 39485 9463 39543 9469
rect 40126 9460 40132 9512
rect 40184 9500 40190 9512
rect 40221 9503 40279 9509
rect 40221 9500 40233 9503
rect 40184 9472 40233 9500
rect 40184 9460 40190 9472
rect 40221 9469 40233 9472
rect 40267 9469 40279 9503
rect 40221 9463 40279 9469
rect 34848 9404 40080 9432
rect 34848 9392 34854 9404
rect 40052 9376 40080 9404
rect 33502 9364 33508 9376
rect 30064 9336 33508 9364
rect 30064 9324 30070 9336
rect 33502 9324 33508 9336
rect 33560 9324 33566 9376
rect 35526 9324 35532 9376
rect 35584 9324 35590 9376
rect 39022 9324 39028 9376
rect 39080 9324 39086 9376
rect 39393 9367 39451 9373
rect 39393 9333 39405 9367
rect 39439 9364 39451 9367
rect 39945 9367 40003 9373
rect 39945 9364 39957 9367
rect 39439 9336 39957 9364
rect 39439 9333 39451 9336
rect 39393 9327 39451 9333
rect 39945 9333 39957 9336
rect 39991 9333 40003 9367
rect 39945 9327 40003 9333
rect 40034 9324 40040 9376
rect 40092 9364 40098 9376
rect 41386 9364 41414 9608
rect 41598 9528 41604 9580
rect 41656 9528 41662 9580
rect 41690 9528 41696 9580
rect 41748 9528 41754 9580
rect 41785 9571 41843 9577
rect 41785 9537 41797 9571
rect 41831 9537 41843 9571
rect 42429 9571 42487 9577
rect 42429 9568 42441 9571
rect 41785 9531 41843 9537
rect 41892 9540 42441 9568
rect 41616 9500 41644 9528
rect 41800 9500 41828 9531
rect 41892 9512 41920 9540
rect 42429 9537 42441 9540
rect 42475 9537 42487 9571
rect 42429 9531 42487 9537
rect 43257 9571 43315 9577
rect 43257 9537 43269 9571
rect 43303 9537 43315 9571
rect 43257 9531 43315 9537
rect 43441 9571 43499 9577
rect 43441 9537 43453 9571
rect 43487 9537 43499 9571
rect 43824 9568 43852 9608
rect 43993 9605 44005 9608
rect 44039 9605 44051 9639
rect 43993 9599 44051 9605
rect 45554 9596 45560 9648
rect 45612 9636 45618 9648
rect 46293 9639 46351 9645
rect 46293 9636 46305 9639
rect 45612 9608 46305 9636
rect 45612 9596 45618 9608
rect 46293 9605 46305 9608
rect 46339 9605 46351 9639
rect 46750 9636 46756 9648
rect 46293 9599 46351 9605
rect 46400 9608 46756 9636
rect 43898 9568 43904 9580
rect 43824 9540 43904 9568
rect 43441 9531 43499 9537
rect 41616 9472 41828 9500
rect 41874 9460 41880 9512
rect 41932 9460 41938 9512
rect 41969 9503 42027 9509
rect 41969 9469 41981 9503
rect 42015 9500 42027 9503
rect 42150 9500 42156 9512
rect 42015 9472 42156 9500
rect 42015 9469 42027 9472
rect 41969 9463 42027 9469
rect 41601 9435 41659 9441
rect 41601 9432 41613 9435
rect 41524 9404 41613 9432
rect 41524 9376 41552 9404
rect 41601 9401 41613 9404
rect 41647 9432 41659 9435
rect 41984 9432 42012 9463
rect 42150 9460 42156 9472
rect 42208 9460 42214 9512
rect 41647 9404 42012 9432
rect 41647 9401 41659 9404
rect 41601 9395 41659 9401
rect 43272 9376 43300 9531
rect 43456 9432 43484 9531
rect 43898 9528 43904 9540
rect 43956 9528 43962 9580
rect 44913 9571 44971 9577
rect 44913 9537 44925 9571
rect 44959 9537 44971 9571
rect 44913 9531 44971 9537
rect 44266 9460 44272 9512
rect 44324 9460 44330 9512
rect 44821 9435 44879 9441
rect 44821 9432 44833 9435
rect 43456 9404 44833 9432
rect 44821 9401 44833 9404
rect 44867 9401 44879 9435
rect 44821 9395 44879 9401
rect 40092 9336 41414 9364
rect 40092 9324 40098 9336
rect 41506 9324 41512 9376
rect 41564 9324 41570 9376
rect 41693 9367 41751 9373
rect 41693 9333 41705 9367
rect 41739 9364 41751 9367
rect 41782 9364 41788 9376
rect 41739 9336 41788 9364
rect 41739 9333 41751 9336
rect 41693 9327 41751 9333
rect 41782 9324 41788 9336
rect 41840 9324 41846 9376
rect 41874 9324 41880 9376
rect 41932 9364 41938 9376
rect 43073 9367 43131 9373
rect 43073 9364 43085 9367
rect 41932 9336 43085 9364
rect 41932 9324 41938 9336
rect 43073 9333 43085 9336
rect 43119 9333 43131 9367
rect 43073 9327 43131 9333
rect 43254 9324 43260 9376
rect 43312 9364 43318 9376
rect 44450 9364 44456 9376
rect 43312 9336 44456 9364
rect 43312 9324 43318 9336
rect 44450 9324 44456 9336
rect 44508 9364 44514 9376
rect 44928 9364 44956 9531
rect 45094 9528 45100 9580
rect 45152 9528 45158 9580
rect 45833 9571 45891 9577
rect 45833 9537 45845 9571
rect 45879 9568 45891 9571
rect 46400 9568 46428 9608
rect 46750 9596 46756 9608
rect 46808 9596 46814 9648
rect 46860 9636 46888 9676
rect 50154 9664 50160 9716
rect 50212 9704 50218 9716
rect 50985 9707 51043 9713
rect 50985 9704 50997 9707
rect 50212 9676 50997 9704
rect 50212 9664 50218 9676
rect 50985 9673 50997 9676
rect 51031 9673 51043 9707
rect 50985 9667 51043 9673
rect 48041 9639 48099 9645
rect 48041 9636 48053 9639
rect 46860 9608 48053 9636
rect 48041 9605 48053 9608
rect 48087 9605 48099 9639
rect 48041 9599 48099 9605
rect 48179 9639 48237 9645
rect 48179 9605 48191 9639
rect 48225 9636 48237 9639
rect 48958 9636 48964 9648
rect 48225 9608 48964 9636
rect 48225 9605 48237 9608
rect 48179 9599 48237 9605
rect 48958 9596 48964 9608
rect 49016 9596 49022 9648
rect 51169 9639 51227 9645
rect 51169 9636 51181 9639
rect 50738 9608 51181 9636
rect 51169 9605 51181 9608
rect 51215 9605 51227 9639
rect 51169 9599 51227 9605
rect 45879 9540 46428 9568
rect 45879 9537 45891 9540
rect 45833 9531 45891 9537
rect 46474 9528 46480 9580
rect 46532 9528 46538 9580
rect 46566 9528 46572 9580
rect 46624 9528 46630 9580
rect 47210 9528 47216 9580
rect 47268 9528 47274 9580
rect 47854 9528 47860 9580
rect 47912 9528 47918 9580
rect 47946 9528 47952 9580
rect 48004 9528 48010 9580
rect 48317 9571 48375 9577
rect 48317 9537 48329 9571
rect 48363 9568 48375 9571
rect 49053 9571 49111 9577
rect 49053 9568 49065 9571
rect 48363 9540 49065 9568
rect 48363 9537 48375 9540
rect 48317 9531 48375 9537
rect 49053 9537 49065 9540
rect 49099 9537 49111 9571
rect 49053 9531 49111 9537
rect 49234 9528 49240 9580
rect 49292 9528 49298 9580
rect 51074 9528 51080 9580
rect 51132 9568 51138 9580
rect 51132 9540 51157 9568
rect 51132 9528 51138 9540
rect 45281 9503 45339 9509
rect 45281 9469 45293 9503
rect 45327 9500 45339 9503
rect 45646 9500 45652 9512
rect 45327 9472 45652 9500
rect 45327 9469 45339 9472
rect 45281 9463 45339 9469
rect 45646 9460 45652 9472
rect 45704 9460 45710 9512
rect 47228 9500 47256 9528
rect 46400 9472 47256 9500
rect 45462 9392 45468 9444
rect 45520 9432 45526 9444
rect 46400 9432 46428 9472
rect 45520 9404 46428 9432
rect 45520 9392 45526 9404
rect 46750 9392 46756 9444
rect 46808 9392 46814 9444
rect 47228 9432 47256 9472
rect 48038 9460 48044 9512
rect 48096 9500 48102 9512
rect 48409 9503 48467 9509
rect 48409 9500 48421 9503
rect 48096 9472 48421 9500
rect 48096 9460 48102 9472
rect 48409 9469 48421 9472
rect 48455 9469 48467 9503
rect 51092 9500 51120 9528
rect 51442 9500 51448 9512
rect 48409 9463 48467 9469
rect 48516 9472 51448 9500
rect 48516 9432 48544 9472
rect 51442 9460 51448 9472
rect 51500 9460 51506 9512
rect 47228 9404 48544 9432
rect 45186 9364 45192 9376
rect 44508 9336 45192 9364
rect 44508 9324 44514 9336
rect 45186 9324 45192 9336
rect 45244 9364 45250 9376
rect 46017 9367 46075 9373
rect 46017 9364 46029 9367
rect 45244 9336 46029 9364
rect 45244 9324 45250 9336
rect 46017 9333 46029 9336
rect 46063 9333 46075 9367
rect 46017 9327 46075 9333
rect 46569 9367 46627 9373
rect 46569 9333 46581 9367
rect 46615 9364 46627 9367
rect 46658 9364 46664 9376
rect 46615 9336 46664 9364
rect 46615 9333 46627 9336
rect 46569 9327 46627 9333
rect 46658 9324 46664 9336
rect 46716 9324 46722 9376
rect 47302 9324 47308 9376
rect 47360 9324 47366 9376
rect 47670 9324 47676 9376
rect 47728 9324 47734 9376
rect 49142 9324 49148 9376
rect 49200 9364 49206 9376
rect 49494 9367 49552 9373
rect 49494 9364 49506 9367
rect 49200 9336 49506 9364
rect 49200 9324 49206 9336
rect 49494 9333 49506 9336
rect 49540 9333 49552 9367
rect 49494 9327 49552 9333
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 23566 9120 23572 9172
rect 23624 9160 23630 9172
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 23624 9132 23673 9160
rect 23624 9120 23630 9132
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 25501 9163 25559 9169
rect 25501 9160 25513 9163
rect 24820 9132 25513 9160
rect 24820 9120 24826 9132
rect 25501 9129 25513 9132
rect 25547 9129 25559 9163
rect 25501 9123 25559 9129
rect 25961 9163 26019 9169
rect 25961 9129 25973 9163
rect 26007 9160 26019 9163
rect 26050 9160 26056 9172
rect 26007 9132 26056 9160
rect 26007 9129 26019 9132
rect 25961 9123 26019 9129
rect 26050 9120 26056 9132
rect 26108 9120 26114 9172
rect 26142 9120 26148 9172
rect 26200 9120 26206 9172
rect 26602 9120 26608 9172
rect 26660 9120 26666 9172
rect 26786 9120 26792 9172
rect 26844 9120 26850 9172
rect 27246 9120 27252 9172
rect 27304 9120 27310 9172
rect 27706 9120 27712 9172
rect 27764 9120 27770 9172
rect 34422 9120 34428 9172
rect 34480 9120 34486 9172
rect 34790 9120 34796 9172
rect 34848 9120 34854 9172
rect 36078 9120 36084 9172
rect 36136 9120 36142 9172
rect 39022 9120 39028 9172
rect 39080 9160 39086 9172
rect 40110 9163 40168 9169
rect 40110 9160 40122 9163
rect 39080 9132 40122 9160
rect 39080 9120 39086 9132
rect 40110 9129 40122 9132
rect 40156 9129 40168 9163
rect 40110 9123 40168 9129
rect 40678 9120 40684 9172
rect 40736 9160 40742 9172
rect 43254 9160 43260 9172
rect 40736 9132 43260 9160
rect 40736 9120 40742 9132
rect 26620 9092 26648 9120
rect 26160 9064 26648 9092
rect 24946 8984 24952 9036
rect 25004 9024 25010 9036
rect 25590 9024 25596 9036
rect 25004 8996 25596 9024
rect 25004 8984 25010 8996
rect 25590 8984 25596 8996
rect 25648 8984 25654 9036
rect 23569 8959 23627 8965
rect 23569 8925 23581 8959
rect 23615 8925 23627 8959
rect 23569 8919 23627 8925
rect 23584 8888 23612 8919
rect 23658 8888 23664 8900
rect 23584 8860 23664 8888
rect 23658 8848 23664 8860
rect 23716 8888 23722 8900
rect 24394 8888 24400 8900
rect 23716 8860 24400 8888
rect 23716 8848 23722 8860
rect 24394 8848 24400 8860
rect 24452 8848 24458 8900
rect 24670 8848 24676 8900
rect 24728 8888 24734 8900
rect 25777 8891 25835 8897
rect 25777 8888 25789 8891
rect 24728 8860 25789 8888
rect 24728 8848 24734 8860
rect 25777 8857 25789 8860
rect 25823 8857 25835 8891
rect 25777 8851 25835 8857
rect 25993 8891 26051 8897
rect 25993 8857 26005 8891
rect 26039 8888 26051 8891
rect 26160 8888 26188 9064
rect 26421 8959 26479 8965
rect 26421 8925 26433 8959
rect 26467 8958 26479 8959
rect 26510 8958 26516 8968
rect 26467 8930 26516 8958
rect 26467 8925 26479 8930
rect 26421 8919 26479 8925
rect 26510 8916 26516 8930
rect 26568 8916 26574 8968
rect 26620 8956 26648 9064
rect 26697 8959 26755 8965
rect 26697 8956 26709 8959
rect 26620 8928 26709 8956
rect 26697 8925 26709 8928
rect 26743 8925 26755 8959
rect 26697 8919 26755 8925
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8956 27215 8959
rect 27264 8956 27292 9120
rect 27433 9027 27491 9033
rect 27433 8993 27445 9027
rect 27479 9024 27491 9027
rect 27724 9024 27752 9120
rect 31665 9095 31723 9101
rect 31665 9061 31677 9095
rect 31711 9061 31723 9095
rect 31665 9055 31723 9061
rect 27893 9027 27951 9033
rect 27893 9024 27905 9027
rect 27479 8996 27568 9024
rect 27724 8996 27905 9024
rect 27479 8993 27491 8996
rect 27433 8987 27491 8993
rect 27203 8928 27292 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 26039 8860 26188 8888
rect 26237 8891 26295 8897
rect 26039 8857 26051 8860
rect 25993 8851 26051 8857
rect 26237 8857 26249 8891
rect 26283 8888 26295 8891
rect 27249 8891 27307 8897
rect 27249 8888 27261 8891
rect 26283 8860 27261 8888
rect 26283 8857 26295 8860
rect 26237 8851 26295 8857
rect 25792 8820 25820 8851
rect 26712 8832 26740 8860
rect 27249 8857 27261 8860
rect 27295 8857 27307 8891
rect 27249 8851 27307 8857
rect 26602 8820 26608 8832
rect 25792 8792 26608 8820
rect 26602 8780 26608 8792
rect 26660 8780 26666 8832
rect 26694 8780 26700 8832
rect 26752 8780 26758 8832
rect 27540 8820 27568 8996
rect 27893 8993 27905 8996
rect 27939 8993 27951 9027
rect 31680 9024 31708 9055
rect 32125 9027 32183 9033
rect 32125 9024 32137 9027
rect 31680 8996 32137 9024
rect 27893 8987 27951 8993
rect 32125 8993 32137 8996
rect 32171 8993 32183 9027
rect 34808 9024 34836 9120
rect 35802 9052 35808 9104
rect 35860 9092 35866 9104
rect 35860 9064 36308 9092
rect 35860 9052 35866 9064
rect 32125 8987 32183 8993
rect 34348 8996 34836 9024
rect 27614 8916 27620 8968
rect 27672 8916 27678 8968
rect 29549 8959 29607 8965
rect 29549 8925 29561 8959
rect 29595 8956 29607 8959
rect 30006 8956 30012 8968
rect 29595 8928 30012 8956
rect 29595 8925 29607 8928
rect 29549 8919 29607 8925
rect 30006 8916 30012 8928
rect 30064 8916 30070 8968
rect 30285 8959 30343 8965
rect 30285 8925 30297 8959
rect 30331 8956 30343 8959
rect 30374 8956 30380 8968
rect 30331 8928 30380 8956
rect 30331 8925 30343 8928
rect 30285 8919 30343 8925
rect 30374 8916 30380 8928
rect 30432 8916 30438 8968
rect 30552 8959 30610 8965
rect 30552 8925 30564 8959
rect 30598 8956 30610 8959
rect 31294 8956 31300 8968
rect 30598 8928 31300 8956
rect 30598 8925 30610 8928
rect 30552 8919 30610 8925
rect 31294 8916 31300 8928
rect 31352 8916 31358 8968
rect 33137 8959 33195 8965
rect 33137 8925 33149 8959
rect 33183 8956 33195 8959
rect 33594 8956 33600 8968
rect 33183 8928 33600 8956
rect 33183 8925 33195 8928
rect 33137 8919 33195 8925
rect 33594 8916 33600 8928
rect 33652 8916 33658 8968
rect 34348 8965 34376 8996
rect 34333 8959 34391 8965
rect 34333 8925 34345 8959
rect 34379 8925 34391 8959
rect 34333 8919 34391 8925
rect 35437 8959 35495 8965
rect 35437 8925 35449 8959
rect 35483 8956 35495 8959
rect 35802 8956 35808 8968
rect 35483 8928 35808 8956
rect 35483 8925 35495 8928
rect 35437 8919 35495 8925
rect 35802 8916 35808 8928
rect 35860 8916 35866 8968
rect 36280 8965 36308 9064
rect 36446 9052 36452 9104
rect 36504 9052 36510 9104
rect 39114 9052 39120 9104
rect 39172 9092 39178 9104
rect 39255 9095 39313 9101
rect 39255 9092 39267 9095
rect 39172 9064 39267 9092
rect 39172 9052 39178 9064
rect 39255 9061 39267 9064
rect 39301 9061 39313 9095
rect 39255 9055 39313 9061
rect 39853 9027 39911 9033
rect 39853 9024 39865 9027
rect 37476 8996 39865 9024
rect 37476 8968 37504 8996
rect 39853 8993 39865 8996
rect 39899 9024 39911 9027
rect 40126 9024 40132 9036
rect 39899 8996 40132 9024
rect 39899 8993 39911 8996
rect 39853 8987 39911 8993
rect 40126 8984 40132 8996
rect 40184 9024 40190 9036
rect 41322 9024 41328 9036
rect 40184 8996 41328 9024
rect 40184 8984 40190 8996
rect 41322 8984 41328 8996
rect 41380 9024 41386 9036
rect 41785 9027 41843 9033
rect 41785 9024 41797 9027
rect 41380 8996 41797 9024
rect 41380 8984 41386 8996
rect 41785 8993 41797 8996
rect 41831 8993 41843 9027
rect 43088 9024 43116 9132
rect 43254 9120 43260 9132
rect 43312 9120 43318 9172
rect 46648 9163 46706 9169
rect 46648 9129 46660 9163
rect 46694 9160 46706 9163
rect 47670 9160 47676 9172
rect 46694 9132 47676 9160
rect 46694 9129 46706 9132
rect 46648 9123 46706 9129
rect 47670 9120 47676 9132
rect 47728 9120 47734 9172
rect 47854 9120 47860 9172
rect 47912 9120 47918 9172
rect 48038 9120 48044 9172
rect 48096 9160 48102 9172
rect 48133 9163 48191 9169
rect 48133 9160 48145 9163
rect 48096 9132 48145 9160
rect 48096 9120 48102 9132
rect 48133 9129 48145 9132
rect 48179 9129 48191 9163
rect 48133 9123 48191 9129
rect 48222 9120 48228 9172
rect 48280 9160 48286 9172
rect 49050 9160 49056 9172
rect 48280 9132 49056 9160
rect 48280 9120 48286 9132
rect 49050 9120 49056 9132
rect 49108 9120 49114 9172
rect 49142 9120 49148 9172
rect 49200 9120 49206 9172
rect 43165 9095 43223 9101
rect 43165 9061 43177 9095
rect 43211 9092 43223 9095
rect 47872 9092 47900 9120
rect 49697 9095 49755 9101
rect 49697 9092 49709 9095
rect 43211 9064 44128 9092
rect 47872 9064 49709 9092
rect 43211 9061 43223 9064
rect 43165 9055 43223 9061
rect 44100 9033 44128 9064
rect 49697 9061 49709 9064
rect 49743 9092 49755 9095
rect 49743 9064 50016 9092
rect 49743 9061 49755 9064
rect 49697 9055 49755 9061
rect 43717 9027 43775 9033
rect 43717 9024 43729 9027
rect 43088 8996 43729 9024
rect 41785 8987 41843 8993
rect 43717 8993 43729 8996
rect 43763 8993 43775 9027
rect 43717 8987 43775 8993
rect 43901 9027 43959 9033
rect 43901 8993 43913 9027
rect 43947 8993 43959 9027
rect 43901 8987 43959 8993
rect 44085 9027 44143 9033
rect 44085 8993 44097 9027
rect 44131 8993 44143 9027
rect 44266 9024 44272 9036
rect 44085 8987 44143 8993
rect 44192 8996 44272 9024
rect 36265 8959 36323 8965
rect 36265 8925 36277 8959
rect 36311 8925 36323 8959
rect 36265 8919 36323 8925
rect 36357 8959 36415 8965
rect 36357 8925 36369 8959
rect 36403 8925 36415 8959
rect 36357 8919 36415 8925
rect 36541 8959 36599 8965
rect 36541 8925 36553 8959
rect 36587 8925 36599 8959
rect 36541 8919 36599 8925
rect 36725 8959 36783 8965
rect 36725 8925 36737 8959
rect 36771 8956 36783 8959
rect 37090 8956 37096 8968
rect 36771 8928 37096 8956
rect 36771 8925 36783 8928
rect 36725 8919 36783 8925
rect 29641 8891 29699 8897
rect 29641 8888 29653 8891
rect 29118 8860 29653 8888
rect 29641 8857 29653 8860
rect 29687 8857 29699 8891
rect 29641 8851 29699 8857
rect 33965 8891 34023 8897
rect 33965 8857 33977 8891
rect 34011 8888 34023 8891
rect 34422 8888 34428 8900
rect 34011 8860 34428 8888
rect 34011 8857 34023 8860
rect 33965 8851 34023 8857
rect 34422 8848 34428 8860
rect 34480 8848 34486 8900
rect 35342 8848 35348 8900
rect 35400 8888 35406 8900
rect 35894 8888 35900 8900
rect 35400 8860 35900 8888
rect 35400 8848 35406 8860
rect 35894 8848 35900 8860
rect 35952 8848 35958 8900
rect 29362 8820 29368 8832
rect 27540 8792 29368 8820
rect 29362 8780 29368 8792
rect 29420 8780 29426 8832
rect 32766 8780 32772 8832
rect 32824 8780 32830 8832
rect 35710 8780 35716 8832
rect 35768 8820 35774 8832
rect 35989 8823 36047 8829
rect 35989 8820 36001 8823
rect 35768 8792 36001 8820
rect 35768 8780 35774 8792
rect 35989 8789 36001 8792
rect 36035 8789 36047 8823
rect 36372 8820 36400 8919
rect 36556 8888 36584 8919
rect 37090 8916 37096 8928
rect 37148 8916 37154 8968
rect 37366 8916 37372 8968
rect 37424 8916 37430 8968
rect 37458 8916 37464 8968
rect 37516 8916 37522 8968
rect 37826 8916 37832 8968
rect 37884 8916 37890 8968
rect 43916 8956 43944 8987
rect 44192 8956 44220 8996
rect 44266 8984 44272 8996
rect 44324 9024 44330 9036
rect 44324 8996 45600 9024
rect 44324 8984 44330 8996
rect 45572 8968 45600 8996
rect 45646 8984 45652 9036
rect 45704 8984 45710 9036
rect 46385 9027 46443 9033
rect 46385 8993 46397 9027
rect 46431 9024 46443 9027
rect 47026 9024 47032 9036
rect 46431 8996 47032 9024
rect 46431 8993 46443 8996
rect 46385 8987 46443 8993
rect 47026 8984 47032 8996
rect 47084 8984 47090 9036
rect 48608 8996 49740 9024
rect 43916 8928 44220 8956
rect 45094 8916 45100 8968
rect 45152 8916 45158 8968
rect 45186 8916 45192 8968
rect 45244 8956 45250 8968
rect 45281 8959 45339 8965
rect 45281 8956 45293 8959
rect 45244 8928 45293 8956
rect 45244 8916 45250 8928
rect 45281 8925 45293 8928
rect 45327 8925 45339 8959
rect 45281 8919 45339 8925
rect 45554 8916 45560 8968
rect 45612 8916 45618 8968
rect 45664 8956 45692 8984
rect 48608 8968 48636 8996
rect 45741 8959 45799 8965
rect 45741 8956 45753 8959
rect 45664 8928 45753 8956
rect 45741 8925 45753 8928
rect 45787 8925 45799 8959
rect 45741 8919 45799 8925
rect 37384 8888 37412 8916
rect 36556 8860 37412 8888
rect 38378 8848 38384 8900
rect 38436 8848 38442 8900
rect 40678 8848 40684 8900
rect 40736 8848 40742 8900
rect 42052 8891 42110 8897
rect 42052 8857 42064 8891
rect 42098 8857 42110 8891
rect 42052 8851 42110 8857
rect 37182 8820 37188 8832
rect 36372 8792 37188 8820
rect 35989 8783 36047 8789
rect 37182 8780 37188 8792
rect 37240 8820 37246 8832
rect 37366 8820 37372 8832
rect 37240 8792 37372 8820
rect 37240 8780 37246 8792
rect 37366 8780 37372 8792
rect 37424 8780 37430 8832
rect 39574 8780 39580 8832
rect 39632 8820 39638 8832
rect 41601 8823 41659 8829
rect 41601 8820 41613 8823
rect 39632 8792 41613 8820
rect 39632 8780 39638 8792
rect 41601 8789 41613 8792
rect 41647 8789 41659 8823
rect 41601 8783 41659 8789
rect 41966 8780 41972 8832
rect 42024 8820 42030 8832
rect 42076 8820 42104 8851
rect 42978 8848 42984 8900
rect 43036 8888 43042 8900
rect 43625 8891 43683 8897
rect 43036 8860 43300 8888
rect 43036 8848 43042 8860
rect 43272 8829 43300 8860
rect 43625 8857 43637 8891
rect 43671 8888 43683 8891
rect 44729 8891 44787 8897
rect 44729 8888 44741 8891
rect 43671 8860 44741 8888
rect 43671 8857 43683 8860
rect 43625 8851 43683 8857
rect 44729 8857 44741 8860
rect 44775 8857 44787 8891
rect 45756 8888 45784 8919
rect 48590 8916 48596 8968
rect 48648 8916 48654 8968
rect 48774 8916 48780 8968
rect 48832 8916 48838 8968
rect 48866 8916 48872 8968
rect 48924 8916 48930 8968
rect 48958 8916 48964 8968
rect 49016 8956 49022 8968
rect 49712 8965 49740 8996
rect 49605 8959 49663 8965
rect 49605 8956 49617 8959
rect 49016 8928 49617 8956
rect 49016 8916 49022 8928
rect 49605 8925 49617 8928
rect 49651 8925 49663 8959
rect 49605 8919 49663 8925
rect 49697 8959 49755 8965
rect 49697 8925 49709 8959
rect 49743 8925 49755 8959
rect 49697 8919 49755 8925
rect 49786 8916 49792 8968
rect 49844 8956 49850 8968
rect 49881 8959 49939 8965
rect 49881 8956 49893 8959
rect 49844 8928 49893 8956
rect 49844 8916 49850 8928
rect 49881 8925 49893 8928
rect 49927 8925 49939 8959
rect 49881 8919 49939 8925
rect 46750 8888 46756 8900
rect 45756 8860 46756 8888
rect 44729 8851 44787 8857
rect 46750 8848 46756 8860
rect 46808 8848 46814 8900
rect 47302 8848 47308 8900
rect 47360 8848 47366 8900
rect 49050 8848 49056 8900
rect 49108 8888 49114 8900
rect 49237 8891 49295 8897
rect 49237 8888 49249 8891
rect 49108 8860 49249 8888
rect 49108 8848 49114 8860
rect 49237 8857 49249 8860
rect 49283 8857 49295 8891
rect 49237 8851 49295 8857
rect 49421 8891 49479 8897
rect 49421 8857 49433 8891
rect 49467 8888 49479 8891
rect 49988 8888 50016 9064
rect 50062 8916 50068 8968
rect 50120 8916 50126 8968
rect 68462 8916 68468 8968
rect 68520 8916 68526 8968
rect 49467 8860 50016 8888
rect 49467 8857 49479 8860
rect 49421 8851 49479 8857
rect 42024 8792 42104 8820
rect 43257 8823 43315 8829
rect 42024 8780 42030 8792
rect 43257 8789 43269 8823
rect 43303 8789 43315 8823
rect 43257 8783 43315 8789
rect 45370 8780 45376 8832
rect 45428 8820 45434 8832
rect 45465 8823 45523 8829
rect 45465 8820 45477 8823
rect 45428 8792 45477 8820
rect 45428 8780 45434 8792
rect 45465 8789 45477 8792
rect 45511 8789 45523 8823
rect 45465 8783 45523 8789
rect 45925 8823 45983 8829
rect 45925 8789 45937 8823
rect 45971 8820 45983 8823
rect 48222 8820 48228 8832
rect 45971 8792 48228 8820
rect 45971 8789 45983 8792
rect 45925 8783 45983 8789
rect 48222 8780 48228 8792
rect 48280 8780 48286 8832
rect 48958 8780 48964 8832
rect 49016 8820 49022 8832
rect 50080 8820 50108 8916
rect 49016 8792 50108 8820
rect 49016 8780 49022 8792
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 23198 8576 23204 8628
rect 23256 8616 23262 8628
rect 25590 8616 25596 8628
rect 23256 8588 25596 8616
rect 23256 8576 23262 8588
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 26142 8576 26148 8628
rect 26200 8576 26206 8628
rect 29362 8616 29368 8628
rect 27908 8588 29368 8616
rect 23216 8489 23244 8576
rect 23474 8508 23480 8560
rect 23532 8508 23538 8560
rect 24486 8508 24492 8560
rect 24544 8508 24550 8560
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 26160 8480 26188 8576
rect 27908 8557 27936 8588
rect 29362 8576 29368 8588
rect 29420 8576 29426 8628
rect 32398 8576 32404 8628
rect 32456 8576 32462 8628
rect 32493 8619 32551 8625
rect 32493 8585 32505 8619
rect 32539 8616 32551 8619
rect 32766 8616 32772 8628
rect 32539 8588 32772 8616
rect 32539 8585 32551 8588
rect 32493 8579 32551 8585
rect 32766 8576 32772 8588
rect 32824 8576 32830 8628
rect 33962 8576 33968 8628
rect 34020 8576 34026 8628
rect 35526 8576 35532 8628
rect 35584 8576 35590 8628
rect 37826 8576 37832 8628
rect 37884 8616 37890 8628
rect 37921 8619 37979 8625
rect 37921 8616 37933 8619
rect 37884 8588 37933 8616
rect 37884 8576 37890 8588
rect 37921 8585 37933 8588
rect 37967 8585 37979 8619
rect 37921 8579 37979 8585
rect 38378 8576 38384 8628
rect 38436 8616 38442 8628
rect 38473 8619 38531 8625
rect 38473 8616 38485 8619
rect 38436 8588 38485 8616
rect 38436 8576 38442 8588
rect 38473 8585 38485 8588
rect 38519 8585 38531 8619
rect 38473 8579 38531 8585
rect 40678 8576 40684 8628
rect 40736 8576 40742 8628
rect 46934 8616 46940 8628
rect 41386 8588 46940 8616
rect 26605 8551 26663 8557
rect 26605 8517 26617 8551
rect 26651 8548 26663 8551
rect 27617 8551 27675 8557
rect 27617 8548 27629 8551
rect 26651 8520 27629 8548
rect 26651 8517 26663 8520
rect 26605 8511 26663 8517
rect 27617 8517 27629 8520
rect 27663 8517 27675 8551
rect 27617 8511 27675 8517
rect 27893 8551 27951 8557
rect 27893 8517 27905 8551
rect 27939 8517 27951 8551
rect 27893 8511 27951 8517
rect 28074 8508 28080 8560
rect 28132 8508 28138 8560
rect 32416 8548 32444 8576
rect 32585 8551 32643 8557
rect 32585 8548 32597 8551
rect 32416 8520 32597 8548
rect 32585 8517 32597 8520
rect 32631 8517 32643 8551
rect 32585 8511 32643 8517
rect 26421 8483 26479 8489
rect 26421 8480 26433 8483
rect 26160 8452 26433 8480
rect 23201 8443 23259 8449
rect 26421 8449 26433 8452
rect 26467 8449 26479 8483
rect 26421 8443 26479 8449
rect 26694 8440 26700 8492
rect 26752 8440 26758 8492
rect 26970 8440 26976 8492
rect 27028 8480 27034 8492
rect 27709 8483 27767 8489
rect 27709 8480 27721 8483
rect 27028 8452 27721 8480
rect 27028 8440 27034 8452
rect 27709 8449 27721 8452
rect 27755 8449 27767 8483
rect 27709 8443 27767 8449
rect 31021 8483 31079 8489
rect 31021 8449 31033 8483
rect 31067 8480 31079 8483
rect 33229 8483 33287 8489
rect 31067 8452 31754 8480
rect 31067 8449 31079 8452
rect 31021 8443 31079 8449
rect 24946 8304 24952 8356
rect 25004 8304 25010 8356
rect 31726 8344 31754 8452
rect 33229 8449 33241 8483
rect 33275 8449 33287 8483
rect 33229 8443 33287 8449
rect 33873 8483 33931 8489
rect 33873 8449 33885 8483
rect 33919 8480 33931 8483
rect 33980 8480 34008 8576
rect 33919 8452 34008 8480
rect 34348 8520 35480 8548
rect 33919 8449 33931 8452
rect 33873 8443 33931 8449
rect 32766 8372 32772 8424
rect 32824 8372 32830 8424
rect 33244 8356 33272 8443
rect 33965 8415 34023 8421
rect 33965 8381 33977 8415
rect 34011 8412 34023 8415
rect 34238 8412 34244 8424
rect 34011 8384 34244 8412
rect 34011 8381 34023 8384
rect 33965 8375 34023 8381
rect 34238 8372 34244 8384
rect 34296 8372 34302 8424
rect 32125 8347 32183 8353
rect 32125 8344 32137 8347
rect 31726 8316 32137 8344
rect 32125 8313 32137 8316
rect 32171 8313 32183 8347
rect 32125 8307 32183 8313
rect 33226 8304 33232 8356
rect 33284 8344 33290 8356
rect 34348 8344 34376 8520
rect 34698 8489 34704 8492
rect 34692 8443 34704 8489
rect 34698 8440 34704 8443
rect 34756 8440 34762 8492
rect 34422 8372 34428 8424
rect 34480 8372 34486 8424
rect 35452 8412 35480 8520
rect 35544 8480 35572 8576
rect 36280 8520 36860 8548
rect 36280 8492 36308 8520
rect 35897 8483 35955 8489
rect 35897 8480 35909 8483
rect 35544 8452 35909 8480
rect 35897 8449 35909 8452
rect 35943 8449 35955 8483
rect 35897 8443 35955 8449
rect 36262 8440 36268 8492
rect 36320 8440 36326 8492
rect 36630 8440 36636 8492
rect 36688 8440 36694 8492
rect 36832 8489 36860 8520
rect 37550 8508 37556 8560
rect 37608 8508 37614 8560
rect 39669 8551 39727 8557
rect 39669 8548 39681 8551
rect 38028 8520 39681 8548
rect 36817 8483 36875 8489
rect 36817 8449 36829 8483
rect 36863 8449 36875 8483
rect 36817 8443 36875 8449
rect 37568 8412 37596 8508
rect 37829 8483 37887 8489
rect 37829 8449 37841 8483
rect 37875 8480 37887 8483
rect 37918 8480 37924 8492
rect 37875 8452 37924 8480
rect 37875 8449 37887 8452
rect 37829 8443 37887 8449
rect 37918 8440 37924 8452
rect 37976 8440 37982 8492
rect 38028 8489 38056 8520
rect 39669 8517 39681 8520
rect 39715 8517 39727 8551
rect 39669 8511 39727 8517
rect 40770 8508 40776 8560
rect 40828 8548 40834 8560
rect 40865 8551 40923 8557
rect 40865 8548 40877 8551
rect 40828 8520 40877 8548
rect 40828 8508 40834 8520
rect 40865 8517 40877 8520
rect 40911 8548 40923 8551
rect 41386 8548 41414 8588
rect 40911 8520 41414 8548
rect 40911 8517 40923 8520
rect 40865 8511 40923 8517
rect 41966 8508 41972 8560
rect 42024 8508 42030 8560
rect 46400 8557 46428 8588
rect 46934 8576 46940 8588
rect 46992 8576 46998 8628
rect 47946 8576 47952 8628
rect 48004 8616 48010 8628
rect 48425 8619 48483 8625
rect 48425 8616 48437 8619
rect 48004 8588 48437 8616
rect 48004 8576 48010 8588
rect 48425 8585 48437 8588
rect 48471 8585 48483 8619
rect 48425 8579 48483 8585
rect 48590 8576 48596 8628
rect 48648 8576 48654 8628
rect 48774 8576 48780 8628
rect 48832 8576 48838 8628
rect 49326 8576 49332 8628
rect 49384 8616 49390 8628
rect 51261 8619 51319 8625
rect 51261 8616 51273 8619
rect 49384 8588 51273 8616
rect 49384 8576 49390 8588
rect 51261 8585 51273 8588
rect 51307 8585 51319 8619
rect 51261 8579 51319 8585
rect 43349 8551 43407 8557
rect 43349 8548 43361 8551
rect 42720 8520 43361 8548
rect 38013 8483 38071 8489
rect 38013 8449 38025 8483
rect 38059 8449 38071 8483
rect 38013 8443 38071 8449
rect 38194 8440 38200 8492
rect 38252 8480 38258 8492
rect 38381 8483 38439 8489
rect 38381 8480 38393 8483
rect 38252 8452 38393 8480
rect 38252 8440 38258 8452
rect 38381 8449 38393 8452
rect 38427 8449 38439 8483
rect 38381 8443 38439 8449
rect 40589 8483 40647 8489
rect 40589 8449 40601 8483
rect 40635 8449 40647 8483
rect 40589 8443 40647 8449
rect 35452 8384 37596 8412
rect 38654 8372 38660 8424
rect 38712 8412 38718 8424
rect 39117 8415 39175 8421
rect 39117 8412 39129 8415
rect 38712 8384 39129 8412
rect 38712 8372 38718 8384
rect 39117 8381 39129 8384
rect 39163 8412 39175 8415
rect 39942 8412 39948 8424
rect 39163 8384 39948 8412
rect 39163 8381 39175 8384
rect 39117 8375 39175 8381
rect 39942 8372 39948 8384
rect 40000 8372 40006 8424
rect 33284 8316 34376 8344
rect 33284 8304 33290 8316
rect 35802 8304 35808 8356
rect 35860 8304 35866 8356
rect 26234 8236 26240 8288
rect 26292 8236 26298 8288
rect 30742 8236 30748 8288
rect 30800 8276 30806 8288
rect 30837 8279 30895 8285
rect 30837 8276 30849 8279
rect 30800 8248 30849 8276
rect 30800 8236 30806 8248
rect 30837 8245 30849 8248
rect 30883 8245 30895 8279
rect 30837 8239 30895 8245
rect 33318 8236 33324 8288
rect 33376 8236 33382 8288
rect 34790 8236 34796 8288
rect 34848 8276 34854 8288
rect 36541 8279 36599 8285
rect 36541 8276 36553 8279
rect 34848 8248 36553 8276
rect 34848 8236 34854 8248
rect 36541 8245 36553 8248
rect 36587 8245 36599 8279
rect 36541 8239 36599 8245
rect 36630 8236 36636 8288
rect 36688 8236 36694 8288
rect 40604 8276 40632 8443
rect 41874 8440 41880 8492
rect 41932 8440 41938 8492
rect 42058 8440 42064 8492
rect 42116 8440 42122 8492
rect 41322 8372 41328 8424
rect 41380 8412 41386 8424
rect 41601 8415 41659 8421
rect 41601 8412 41613 8415
rect 41380 8384 41613 8412
rect 41380 8372 41386 8384
rect 41601 8381 41613 8384
rect 41647 8381 41659 8415
rect 41601 8375 41659 8381
rect 42720 8353 42748 8520
rect 43349 8517 43361 8520
rect 43395 8517 43407 8551
rect 45005 8551 45063 8557
rect 45005 8548 45017 8551
rect 44574 8520 45017 8548
rect 43349 8511 43407 8517
rect 45005 8517 45017 8520
rect 45051 8517 45063 8551
rect 45005 8511 45063 8517
rect 46385 8551 46443 8557
rect 46385 8517 46397 8551
rect 46431 8517 46443 8551
rect 46385 8511 46443 8517
rect 46566 8508 46572 8560
rect 46624 8508 46630 8560
rect 48038 8508 48044 8560
rect 48096 8548 48102 8560
rect 48225 8551 48283 8557
rect 48225 8548 48237 8551
rect 48096 8520 48237 8548
rect 48096 8508 48102 8520
rect 48225 8517 48237 8520
rect 48271 8517 48283 8551
rect 49694 8548 49700 8560
rect 48225 8511 48283 8517
rect 48700 8520 49700 8548
rect 42889 8483 42947 8489
rect 42889 8449 42901 8483
rect 42935 8480 42947 8483
rect 42978 8480 42984 8492
rect 42935 8452 42984 8480
rect 42935 8449 42947 8452
rect 42889 8443 42947 8449
rect 42978 8440 42984 8452
rect 43036 8440 43042 8492
rect 44726 8440 44732 8492
rect 44784 8480 44790 8492
rect 44913 8483 44971 8489
rect 44913 8480 44925 8483
rect 44784 8452 44925 8480
rect 44784 8440 44790 8452
rect 44913 8449 44925 8452
rect 44959 8480 44971 8483
rect 45462 8480 45468 8492
rect 44959 8452 45468 8480
rect 44959 8449 44971 8452
rect 44913 8443 44971 8449
rect 45462 8440 45468 8452
rect 45520 8440 45526 8492
rect 45738 8440 45744 8492
rect 45796 8480 45802 8492
rect 45889 8483 45947 8489
rect 45889 8480 45901 8483
rect 45796 8452 45901 8480
rect 45796 8440 45802 8452
rect 45889 8449 45901 8452
rect 45935 8449 45947 8483
rect 45889 8443 45947 8449
rect 46014 8440 46020 8492
rect 46072 8440 46078 8492
rect 46109 8483 46167 8489
rect 46109 8449 46121 8483
rect 46155 8480 46167 8483
rect 46198 8480 46204 8492
rect 46155 8452 46204 8480
rect 46155 8449 46167 8452
rect 46109 8443 46167 8449
rect 46198 8440 46204 8452
rect 46256 8440 46262 8492
rect 46293 8483 46351 8489
rect 46293 8449 46305 8483
rect 46339 8480 46351 8483
rect 46584 8480 46612 8508
rect 46339 8452 46612 8480
rect 46339 8449 46351 8452
rect 46293 8443 46351 8449
rect 46750 8440 46756 8492
rect 46808 8480 46814 8492
rect 48700 8489 48728 8520
rect 49694 8508 49700 8520
rect 49752 8508 49758 8560
rect 51537 8551 51595 8557
rect 51537 8548 51549 8551
rect 51014 8520 51549 8548
rect 51537 8517 51549 8520
rect 51583 8517 51595 8551
rect 51537 8511 51595 8517
rect 48685 8483 48743 8489
rect 48685 8480 48697 8483
rect 46808 8452 48697 8480
rect 46808 8440 46814 8452
rect 48685 8449 48697 8452
rect 48731 8449 48743 8483
rect 48685 8443 48743 8449
rect 48866 8440 48872 8492
rect 48924 8440 48930 8492
rect 51442 8440 51448 8492
rect 51500 8440 51506 8492
rect 43073 8415 43131 8421
rect 43073 8381 43085 8415
rect 43119 8412 43131 8415
rect 47026 8412 47032 8424
rect 43119 8384 47032 8412
rect 43119 8381 43131 8384
rect 43073 8375 43131 8381
rect 47026 8372 47032 8384
rect 47084 8412 47090 8424
rect 47121 8415 47179 8421
rect 47121 8412 47133 8415
rect 47084 8384 47133 8412
rect 47084 8372 47090 8384
rect 47121 8381 47133 8384
rect 47167 8412 47179 8415
rect 49513 8415 49571 8421
rect 49513 8412 49525 8415
rect 47167 8384 49525 8412
rect 47167 8381 47179 8384
rect 47121 8375 47179 8381
rect 49513 8381 49525 8384
rect 49559 8381 49571 8415
rect 49513 8375 49571 8381
rect 49786 8372 49792 8424
rect 49844 8372 49850 8424
rect 42705 8347 42763 8353
rect 42705 8313 42717 8347
rect 42751 8313 42763 8347
rect 42705 8307 42763 8313
rect 44821 8347 44879 8353
rect 44821 8313 44833 8347
rect 44867 8344 44879 8347
rect 45554 8344 45560 8356
rect 44867 8316 45560 8344
rect 44867 8313 44879 8316
rect 44821 8307 44879 8313
rect 45554 8304 45560 8316
rect 45612 8304 45618 8356
rect 46014 8304 46020 8356
rect 46072 8344 46078 8356
rect 46072 8316 48452 8344
rect 46072 8304 46078 8316
rect 44726 8276 44732 8288
rect 40604 8248 44732 8276
rect 44726 8236 44732 8248
rect 44784 8236 44790 8288
rect 48424 8285 48452 8316
rect 48409 8279 48467 8285
rect 48409 8245 48421 8279
rect 48455 8276 48467 8279
rect 49326 8276 49332 8288
rect 48455 8248 49332 8276
rect 48455 8245 48467 8248
rect 48409 8239 48467 8245
rect 49326 8236 49332 8248
rect 49384 8236 49390 8288
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 24486 8032 24492 8084
rect 24544 8032 24550 8084
rect 26970 8032 26976 8084
rect 27028 8072 27034 8084
rect 27065 8075 27123 8081
rect 27065 8072 27077 8075
rect 27028 8044 27077 8072
rect 27028 8032 27034 8044
rect 27065 8041 27077 8044
rect 27111 8041 27123 8075
rect 27065 8035 27123 8041
rect 32125 8075 32183 8081
rect 32125 8041 32137 8075
rect 32171 8072 32183 8075
rect 32214 8072 32220 8084
rect 32171 8044 32220 8072
rect 32171 8041 32183 8044
rect 32125 8035 32183 8041
rect 32214 8032 32220 8044
rect 32272 8072 32278 8084
rect 32766 8072 32772 8084
rect 32272 8044 32772 8072
rect 32272 8032 32278 8044
rect 32766 8032 32772 8044
rect 32824 8032 32830 8084
rect 34514 8032 34520 8084
rect 34572 8032 34578 8084
rect 34698 8032 34704 8084
rect 34756 8032 34762 8084
rect 36280 8044 39712 8072
rect 34532 8004 34560 8032
rect 36280 8016 36308 8044
rect 36262 8004 36268 8016
rect 34532 7976 36268 8004
rect 36262 7964 36268 7976
rect 36320 7964 36326 8016
rect 37737 8007 37795 8013
rect 37737 7973 37749 8007
rect 37783 8004 37795 8007
rect 37783 7976 38700 8004
rect 37783 7973 37795 7976
rect 37737 7967 37795 7973
rect 25317 7939 25375 7945
rect 25317 7905 25329 7939
rect 25363 7936 25375 7939
rect 25590 7936 25596 7948
rect 25363 7908 25596 7936
rect 25363 7905 25375 7908
rect 25317 7899 25375 7905
rect 25590 7896 25596 7908
rect 25648 7936 25654 7948
rect 27614 7936 27620 7948
rect 25648 7908 27620 7936
rect 25648 7896 25654 7908
rect 27614 7896 27620 7908
rect 27672 7896 27678 7948
rect 29365 7939 29423 7945
rect 29365 7905 29377 7939
rect 29411 7936 29423 7939
rect 29914 7936 29920 7948
rect 29411 7908 29920 7936
rect 29411 7905 29423 7908
rect 29365 7899 29423 7905
rect 29914 7896 29920 7908
rect 29972 7896 29978 7948
rect 30374 7896 30380 7948
rect 30432 7936 30438 7948
rect 32217 7939 32275 7945
rect 32217 7936 32229 7939
rect 30432 7908 32229 7936
rect 30432 7896 30438 7908
rect 32217 7905 32229 7908
rect 32263 7936 32275 7939
rect 32766 7936 32772 7948
rect 32263 7908 32772 7936
rect 32263 7905 32275 7908
rect 32217 7899 32275 7905
rect 32766 7896 32772 7908
rect 32824 7896 32830 7948
rect 36357 7939 36415 7945
rect 36357 7936 36369 7939
rect 34440 7908 36369 7936
rect 34440 7880 34468 7908
rect 36357 7905 36369 7908
rect 36403 7905 36415 7939
rect 36357 7899 36415 7905
rect 37918 7896 37924 7948
rect 37976 7936 37982 7948
rect 38289 7939 38347 7945
rect 38289 7936 38301 7939
rect 37976 7908 38301 7936
rect 37976 7896 37982 7908
rect 38289 7905 38301 7908
rect 38335 7905 38347 7939
rect 38289 7899 38347 7905
rect 38473 7939 38531 7945
rect 38473 7905 38485 7939
rect 38519 7936 38531 7939
rect 38562 7936 38568 7948
rect 38519 7908 38568 7936
rect 38519 7905 38531 7908
rect 38473 7899 38531 7905
rect 38562 7896 38568 7908
rect 38620 7896 38626 7948
rect 38672 7945 38700 7976
rect 38657 7939 38715 7945
rect 38657 7905 38669 7939
rect 38703 7905 38715 7939
rect 38657 7899 38715 7905
rect 934 7828 940 7880
rect 992 7868 998 7880
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 992 7840 1593 7868
rect 992 7828 998 7840
rect 1581 7837 1593 7840
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 24394 7828 24400 7880
rect 24452 7868 24458 7880
rect 24452 7840 24808 7868
rect 24452 7828 24458 7840
rect 24780 7812 24808 7840
rect 29822 7828 29828 7880
rect 29880 7828 29886 7880
rect 30009 7871 30067 7877
rect 30009 7837 30021 7871
rect 30055 7837 30067 7871
rect 30009 7831 30067 7837
rect 24762 7760 24768 7812
rect 24820 7760 24826 7812
rect 25593 7803 25651 7809
rect 25593 7769 25605 7803
rect 25639 7769 25651 7803
rect 25593 7763 25651 7769
rect 25608 7732 25636 7763
rect 26326 7760 26332 7812
rect 26384 7760 26390 7812
rect 27890 7760 27896 7812
rect 27948 7760 27954 7812
rect 29270 7800 29276 7812
rect 29118 7772 29276 7800
rect 29270 7760 29276 7772
rect 29328 7760 29334 7812
rect 30024 7800 30052 7831
rect 31938 7828 31944 7880
rect 31996 7868 32002 7880
rect 32585 7871 32643 7877
rect 32585 7868 32597 7871
rect 31996 7840 32597 7868
rect 31996 7828 32002 7840
rect 32585 7837 32597 7840
rect 32631 7837 32643 7871
rect 32585 7831 32643 7837
rect 34422 7828 34428 7880
rect 34480 7828 34486 7880
rect 34514 7828 34520 7880
rect 34572 7828 34578 7880
rect 34701 7871 34759 7877
rect 34701 7837 34713 7871
rect 34747 7868 34759 7871
rect 34790 7868 34796 7880
rect 34747 7840 34796 7868
rect 34747 7837 34759 7840
rect 34701 7831 34759 7837
rect 34790 7828 34796 7840
rect 34848 7828 34854 7880
rect 34885 7871 34943 7877
rect 34885 7837 34897 7871
rect 34931 7868 34943 7871
rect 34977 7871 35035 7877
rect 34977 7868 34989 7871
rect 34931 7840 34989 7868
rect 34931 7837 34943 7840
rect 34885 7831 34943 7837
rect 34977 7837 34989 7840
rect 35023 7837 35035 7871
rect 34977 7831 35035 7837
rect 30374 7800 30380 7812
rect 30024 7772 30380 7800
rect 30374 7760 30380 7772
rect 30432 7760 30438 7812
rect 30653 7803 30711 7809
rect 30653 7769 30665 7803
rect 30699 7800 30711 7803
rect 30742 7800 30748 7812
rect 30699 7772 30748 7800
rect 30699 7769 30711 7772
rect 30653 7763 30711 7769
rect 30742 7760 30748 7772
rect 30800 7760 30806 7812
rect 31662 7760 31668 7812
rect 31720 7760 31726 7812
rect 33318 7760 33324 7812
rect 33376 7760 33382 7812
rect 34532 7800 34560 7828
rect 34900 7800 34928 7831
rect 35250 7828 35256 7880
rect 35308 7828 35314 7880
rect 36630 7877 36636 7880
rect 35345 7871 35403 7877
rect 35345 7837 35357 7871
rect 35391 7837 35403 7871
rect 36624 7868 36636 7877
rect 36591 7840 36636 7868
rect 35345 7831 35403 7837
rect 36624 7831 36636 7840
rect 35360 7800 35388 7831
rect 36630 7828 36636 7831
rect 36688 7828 36694 7880
rect 39577 7871 39635 7877
rect 39577 7868 39589 7871
rect 37844 7840 39589 7868
rect 34532 7772 34928 7800
rect 35084 7772 35388 7800
rect 26234 7732 26240 7744
rect 25608 7704 26240 7732
rect 26234 7692 26240 7704
rect 26292 7692 26298 7744
rect 29546 7692 29552 7744
rect 29604 7732 29610 7744
rect 29641 7735 29699 7741
rect 29641 7732 29653 7735
rect 29604 7704 29653 7732
rect 29604 7692 29610 7704
rect 29641 7701 29653 7704
rect 29687 7701 29699 7735
rect 29641 7695 29699 7701
rect 30006 7692 30012 7744
rect 30064 7732 30070 7744
rect 30101 7735 30159 7741
rect 30101 7732 30113 7735
rect 30064 7704 30113 7732
rect 30064 7692 30070 7704
rect 30101 7701 30113 7704
rect 30147 7701 30159 7735
rect 30101 7695 30159 7701
rect 33410 7692 33416 7744
rect 33468 7732 33474 7744
rect 35084 7741 35112 7772
rect 34011 7735 34069 7741
rect 34011 7732 34023 7735
rect 33468 7704 34023 7732
rect 33468 7692 33474 7704
rect 34011 7701 34023 7704
rect 34057 7701 34069 7735
rect 34011 7695 34069 7701
rect 35075 7735 35133 7741
rect 35075 7701 35087 7735
rect 35121 7701 35133 7735
rect 35075 7695 35133 7701
rect 35161 7735 35219 7741
rect 35161 7701 35173 7735
rect 35207 7732 35219 7735
rect 35894 7732 35900 7744
rect 35207 7704 35900 7732
rect 35207 7701 35219 7704
rect 35161 7695 35219 7701
rect 35894 7692 35900 7704
rect 35952 7692 35958 7744
rect 35986 7692 35992 7744
rect 36044 7692 36050 7744
rect 37844 7741 37872 7840
rect 39577 7837 39589 7840
rect 39623 7837 39635 7871
rect 39577 7831 39635 7837
rect 38197 7803 38255 7809
rect 38197 7769 38209 7803
rect 38243 7800 38255 7803
rect 39301 7803 39359 7809
rect 39301 7800 39313 7803
rect 38243 7772 39313 7800
rect 38243 7769 38255 7772
rect 38197 7763 38255 7769
rect 39301 7769 39313 7772
rect 39347 7769 39359 7803
rect 39684 7800 39712 8044
rect 45738 8032 45744 8084
rect 45796 8032 45802 8084
rect 45830 8032 45836 8084
rect 45888 8032 45894 8084
rect 46753 8075 46811 8081
rect 46753 8041 46765 8075
rect 46799 8041 46811 8075
rect 47946 8072 47952 8084
rect 46753 8035 46811 8041
rect 47504 8044 47952 8072
rect 42337 8007 42395 8013
rect 42337 8004 42349 8007
rect 41064 7976 42349 8004
rect 41064 7877 41092 7976
rect 42337 7973 42349 7976
rect 42383 7973 42395 8007
rect 45756 8004 45784 8032
rect 46106 8004 46112 8016
rect 45756 7976 46112 8004
rect 42337 7967 42395 7973
rect 46106 7964 46112 7976
rect 46164 8004 46170 8016
rect 46768 8004 46796 8035
rect 46164 7976 46796 8004
rect 46937 8007 46995 8013
rect 46164 7964 46170 7976
rect 46937 7973 46949 8007
rect 46983 7973 46995 8007
rect 46937 7967 46995 7973
rect 41397 7939 41455 7945
rect 41397 7905 41409 7939
rect 41443 7936 41455 7939
rect 41693 7939 41751 7945
rect 41693 7936 41705 7939
rect 41443 7908 41705 7936
rect 41443 7905 41455 7908
rect 41397 7899 41455 7905
rect 41693 7905 41705 7908
rect 41739 7905 41751 7939
rect 44085 7939 44143 7945
rect 44085 7936 44097 7939
rect 41693 7899 41751 7905
rect 43180 7908 44097 7936
rect 41049 7871 41107 7877
rect 41049 7837 41061 7871
rect 41095 7837 41107 7871
rect 41049 7831 41107 7837
rect 41233 7871 41291 7877
rect 41233 7837 41245 7871
rect 41279 7837 41291 7871
rect 41233 7831 41291 7837
rect 41601 7871 41659 7877
rect 41601 7837 41613 7871
rect 41647 7868 41659 7871
rect 41782 7868 41788 7880
rect 41647 7840 41788 7868
rect 41647 7837 41659 7840
rect 41601 7831 41659 7837
rect 41248 7800 41276 7831
rect 41782 7828 41788 7840
rect 41840 7868 41846 7880
rect 42150 7868 42156 7880
rect 41840 7840 42156 7868
rect 41840 7828 41846 7840
rect 42150 7828 42156 7840
rect 42208 7828 42214 7880
rect 42426 7828 42432 7880
rect 42484 7828 42490 7880
rect 43180 7877 43208 7908
rect 44085 7905 44097 7908
rect 44131 7905 44143 7939
rect 46952 7936 46980 7967
rect 44085 7899 44143 7905
rect 46308 7908 46980 7936
rect 43165 7871 43223 7877
rect 43165 7837 43177 7871
rect 43211 7837 43223 7871
rect 43165 7831 43223 7837
rect 43530 7828 43536 7880
rect 43588 7828 43594 7880
rect 46014 7871 46072 7877
rect 46014 7837 46026 7871
rect 46060 7868 46072 7871
rect 46308 7868 46336 7908
rect 46060 7840 46336 7868
rect 46060 7837 46072 7840
rect 46014 7831 46072 7837
rect 46382 7828 46388 7880
rect 46440 7828 46446 7880
rect 46477 7871 46535 7877
rect 46477 7837 46489 7871
rect 46523 7837 46535 7871
rect 46477 7831 46535 7837
rect 39684 7772 41276 7800
rect 39301 7763 39359 7769
rect 37829 7735 37887 7741
rect 37829 7701 37841 7735
rect 37875 7701 37887 7735
rect 37829 7695 37887 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 41138 7692 41144 7744
rect 41196 7692 41202 7744
rect 41248 7732 41276 7772
rect 41325 7803 41383 7809
rect 41325 7769 41337 7803
rect 41371 7800 41383 7803
rect 41414 7800 41420 7812
rect 41371 7772 41420 7800
rect 41371 7769 41383 7772
rect 41325 7763 41383 7769
rect 41414 7760 41420 7772
rect 41472 7760 41478 7812
rect 41509 7803 41567 7809
rect 41509 7769 41521 7803
rect 41555 7800 41567 7803
rect 43073 7803 43131 7809
rect 43073 7800 43085 7803
rect 41555 7772 43085 7800
rect 41555 7769 41567 7772
rect 41509 7763 41567 7769
rect 43073 7769 43085 7772
rect 43119 7769 43131 7803
rect 43073 7763 43131 7769
rect 46198 7760 46204 7812
rect 46256 7800 46262 7812
rect 46492 7800 46520 7831
rect 46658 7828 46664 7880
rect 46716 7828 46722 7880
rect 47504 7877 47532 8044
rect 47946 8032 47952 8044
rect 48004 8072 48010 8084
rect 48133 8075 48191 8081
rect 48133 8072 48145 8075
rect 48004 8044 48145 8072
rect 48004 8032 48010 8044
rect 48133 8041 48145 8044
rect 48179 8041 48191 8075
rect 48133 8035 48191 8041
rect 48409 8075 48467 8081
rect 48409 8041 48421 8075
rect 48455 8041 48467 8075
rect 48409 8035 48467 8041
rect 49605 8075 49663 8081
rect 49605 8041 49617 8075
rect 49651 8072 49663 8075
rect 49786 8072 49792 8084
rect 49651 8044 49792 8072
rect 49651 8041 49663 8044
rect 49605 8035 49663 8041
rect 48424 8004 48452 8035
rect 49786 8032 49792 8044
rect 49844 8032 49850 8084
rect 47872 7976 48452 8004
rect 48777 8007 48835 8013
rect 47762 7896 47768 7948
rect 47820 7896 47826 7948
rect 47489 7871 47547 7877
rect 47489 7837 47501 7871
rect 47535 7837 47547 7871
rect 47489 7831 47547 7837
rect 47670 7828 47676 7880
rect 47728 7868 47734 7880
rect 47872 7878 47900 7976
rect 48777 7973 48789 8007
rect 48823 8004 48835 8007
rect 48823 7976 49832 8004
rect 48823 7973 48835 7976
rect 48777 7967 48835 7973
rect 48286 7908 48452 7936
rect 47935 7881 47993 7887
rect 47935 7878 47947 7881
rect 47872 7868 47947 7878
rect 47728 7850 47947 7868
rect 47728 7840 47900 7850
rect 47935 7847 47947 7850
rect 47981 7847 47993 7881
rect 48286 7868 48314 7908
rect 48148 7864 48314 7868
rect 47935 7841 47993 7847
rect 48056 7840 48314 7864
rect 47728 7828 47734 7840
rect 48056 7836 48176 7840
rect 46569 7803 46627 7809
rect 46569 7800 46581 7803
rect 46256 7772 46581 7800
rect 46256 7760 46262 7772
rect 46569 7769 46581 7772
rect 46615 7769 46627 7803
rect 46676 7800 46704 7828
rect 46769 7803 46827 7809
rect 46769 7800 46781 7803
rect 46676 7772 46781 7800
rect 46569 7763 46627 7769
rect 46769 7769 46781 7772
rect 46815 7769 46827 7803
rect 46769 7763 46827 7769
rect 47581 7803 47639 7809
rect 47581 7769 47593 7803
rect 47627 7800 47639 7803
rect 48056 7800 48084 7836
rect 48424 7812 48452 7908
rect 49326 7896 49332 7948
rect 49384 7896 49390 7948
rect 49804 7877 49832 7976
rect 49789 7871 49847 7877
rect 49789 7837 49801 7871
rect 49835 7837 49847 7871
rect 49789 7831 49847 7837
rect 48225 7803 48283 7809
rect 48225 7800 48237 7803
rect 47627 7772 48084 7800
rect 48148 7772 48237 7800
rect 47627 7769 47639 7772
rect 47581 7763 47639 7769
rect 42058 7732 42064 7744
rect 41248 7704 42064 7732
rect 42058 7692 42064 7704
rect 42116 7692 42122 7744
rect 42794 7692 42800 7744
rect 42852 7732 42858 7744
rect 43257 7735 43315 7741
rect 43257 7732 43269 7735
rect 42852 7704 43269 7732
rect 42852 7692 42858 7704
rect 43257 7701 43269 7704
rect 43303 7701 43315 7735
rect 43257 7695 43315 7701
rect 46014 7692 46020 7744
rect 46072 7692 46078 7744
rect 46584 7732 46612 7763
rect 48148 7744 48176 7772
rect 48225 7769 48237 7772
rect 48271 7769 48283 7803
rect 48225 7763 48283 7769
rect 48406 7760 48412 7812
rect 48464 7809 48470 7812
rect 48464 7803 48483 7809
rect 48471 7769 48483 7803
rect 49237 7803 49295 7809
rect 49237 7800 49249 7803
rect 48464 7763 48483 7769
rect 48516 7772 49249 7800
rect 48464 7760 48470 7763
rect 47762 7732 47768 7744
rect 46584 7704 47768 7732
rect 47762 7692 47768 7704
rect 47820 7692 47826 7744
rect 48130 7692 48136 7744
rect 48188 7692 48194 7744
rect 48314 7692 48320 7744
rect 48372 7732 48378 7744
rect 48516 7732 48544 7772
rect 49237 7769 49249 7772
rect 49283 7800 49295 7803
rect 49510 7800 49516 7812
rect 49283 7772 49516 7800
rect 49283 7769 49295 7772
rect 49237 7763 49295 7769
rect 49510 7760 49516 7772
rect 49568 7760 49574 7812
rect 48372 7704 48544 7732
rect 48372 7692 48378 7704
rect 48590 7692 48596 7744
rect 48648 7692 48654 7744
rect 49142 7692 49148 7744
rect 49200 7692 49206 7744
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 26326 7488 26332 7540
rect 26384 7488 26390 7540
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 28905 7531 28963 7537
rect 28905 7528 28917 7531
rect 27948 7500 28917 7528
rect 27948 7488 27954 7500
rect 28905 7497 28917 7500
rect 28951 7497 28963 7531
rect 28905 7491 28963 7497
rect 29270 7488 29276 7540
rect 29328 7488 29334 7540
rect 31573 7531 31631 7537
rect 29380 7500 31524 7528
rect 24762 7420 24768 7472
rect 24820 7460 24826 7472
rect 29380 7460 29408 7500
rect 29546 7460 29552 7472
rect 24820 7432 29408 7460
rect 24820 7420 24826 7432
rect 26252 7401 26280 7432
rect 26237 7395 26295 7401
rect 26237 7361 26249 7395
rect 26283 7361 26295 7395
rect 26237 7355 26295 7361
rect 28445 7395 28503 7401
rect 28445 7361 28457 7395
rect 28491 7392 28503 7395
rect 28994 7392 29000 7404
rect 28491 7364 29000 7392
rect 28491 7361 28503 7364
rect 28445 7355 28503 7361
rect 28994 7352 29000 7364
rect 29052 7352 29058 7404
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 29181 7395 29239 7401
rect 29181 7361 29193 7395
rect 29227 7392 29239 7395
rect 29380 7392 29408 7432
rect 29472 7432 29552 7460
rect 29472 7401 29500 7432
rect 29546 7420 29552 7432
rect 29604 7420 29610 7472
rect 30745 7463 30803 7469
rect 30745 7429 30757 7463
rect 30791 7460 30803 7463
rect 31110 7460 31116 7472
rect 30791 7432 31116 7460
rect 30791 7429 30803 7432
rect 30745 7423 30803 7429
rect 31110 7420 31116 7432
rect 31168 7420 31174 7472
rect 29227 7364 29408 7392
rect 29457 7395 29515 7401
rect 29227 7361 29239 7364
rect 29181 7355 29239 7361
rect 29457 7361 29469 7395
rect 29503 7361 29515 7395
rect 29641 7395 29699 7401
rect 29641 7392 29653 7395
rect 29457 7355 29515 7361
rect 29564 7364 29653 7392
rect 28534 7284 28540 7336
rect 28592 7284 28598 7336
rect 28626 7284 28632 7336
rect 28684 7333 28690 7336
rect 28684 7327 28733 7333
rect 28684 7293 28687 7327
rect 28721 7293 28733 7327
rect 28684 7287 28733 7293
rect 28684 7284 28690 7287
rect 28810 7284 28816 7336
rect 28868 7324 28874 7336
rect 29104 7324 29132 7355
rect 28868 7296 29132 7324
rect 28868 7284 28874 7296
rect 28077 7259 28135 7265
rect 28077 7225 28089 7259
rect 28123 7256 28135 7259
rect 28442 7256 28448 7268
rect 28123 7228 28448 7256
rect 28123 7225 28135 7228
rect 28077 7219 28135 7225
rect 28442 7216 28448 7228
rect 28500 7216 28506 7268
rect 29564 7256 29592 7364
rect 29641 7361 29653 7364
rect 29687 7361 29699 7395
rect 29641 7355 29699 7361
rect 30098 7352 30104 7404
rect 30156 7392 30162 7404
rect 31496 7401 31524 7500
rect 31573 7497 31585 7531
rect 31619 7528 31631 7531
rect 31662 7528 31668 7540
rect 31619 7500 31668 7528
rect 31619 7497 31631 7500
rect 31573 7491 31631 7497
rect 31662 7488 31668 7500
rect 31720 7488 31726 7540
rect 31938 7488 31944 7540
rect 31996 7488 32002 7540
rect 32861 7531 32919 7537
rect 32861 7528 32873 7531
rect 32600 7500 32873 7528
rect 32398 7460 32404 7472
rect 31772 7432 32404 7460
rect 30193 7395 30251 7401
rect 30193 7392 30205 7395
rect 30156 7364 30205 7392
rect 30156 7352 30162 7364
rect 30193 7361 30205 7364
rect 30239 7361 30251 7395
rect 30193 7355 30251 7361
rect 30377 7395 30435 7401
rect 30377 7361 30389 7395
rect 30423 7392 30435 7395
rect 31481 7395 31539 7401
rect 30423 7364 31064 7392
rect 30423 7361 30435 7364
rect 30377 7355 30435 7361
rect 30374 7256 30380 7268
rect 29564 7228 30380 7256
rect 30374 7216 30380 7228
rect 30432 7216 30438 7268
rect 28626 7148 28632 7200
rect 28684 7188 28690 7200
rect 29914 7188 29920 7200
rect 28684 7160 29920 7188
rect 28684 7148 28690 7160
rect 29914 7148 29920 7160
rect 29972 7148 29978 7200
rect 31036 7188 31064 7364
rect 31481 7361 31493 7395
rect 31527 7392 31539 7395
rect 31570 7392 31576 7404
rect 31527 7364 31576 7392
rect 31527 7361 31539 7364
rect 31481 7355 31539 7361
rect 31570 7352 31576 7364
rect 31628 7352 31634 7404
rect 31662 7352 31668 7404
rect 31720 7392 31726 7404
rect 31772 7401 31800 7432
rect 32398 7420 32404 7432
rect 32456 7420 32462 7472
rect 31757 7395 31815 7401
rect 31757 7392 31769 7395
rect 31720 7364 31769 7392
rect 31720 7352 31726 7364
rect 31757 7361 31769 7364
rect 31803 7361 31815 7395
rect 31757 7355 31815 7361
rect 31941 7395 31999 7401
rect 31941 7361 31953 7395
rect 31987 7392 31999 7395
rect 32600 7392 32628 7500
rect 32861 7497 32873 7500
rect 32907 7497 32919 7531
rect 32861 7491 32919 7497
rect 33410 7488 33416 7540
rect 33468 7488 33474 7540
rect 33505 7531 33563 7537
rect 33505 7497 33517 7531
rect 33551 7528 33563 7531
rect 33686 7528 33692 7540
rect 33551 7500 33692 7528
rect 33551 7497 33563 7500
rect 33505 7491 33563 7497
rect 33686 7488 33692 7500
rect 33744 7488 33750 7540
rect 35986 7488 35992 7540
rect 36044 7488 36050 7540
rect 39390 7528 39396 7540
rect 38488 7500 39396 7528
rect 35152 7463 35210 7469
rect 35152 7429 35164 7463
rect 35198 7460 35210 7463
rect 36004 7460 36032 7488
rect 38488 7469 38516 7500
rect 39390 7488 39396 7500
rect 39448 7488 39454 7540
rect 40129 7531 40187 7537
rect 40129 7497 40141 7531
rect 40175 7497 40187 7531
rect 40129 7491 40187 7497
rect 42245 7531 42303 7537
rect 42245 7497 42257 7531
rect 42291 7528 42303 7531
rect 42426 7528 42432 7540
rect 42291 7500 42432 7528
rect 42291 7497 42303 7500
rect 42245 7491 42303 7497
rect 35198 7432 36032 7460
rect 38473 7463 38531 7469
rect 35198 7429 35210 7432
rect 35152 7423 35210 7429
rect 38473 7429 38485 7463
rect 38519 7429 38531 7463
rect 40144 7460 40172 7491
rect 41322 7460 41328 7472
rect 39698 7432 40172 7460
rect 40880 7432 41328 7460
rect 38473 7423 38531 7429
rect 34422 7392 34428 7404
rect 31987 7364 32628 7392
rect 32784 7364 34428 7392
rect 31987 7361 31999 7364
rect 31941 7355 31999 7361
rect 32784 7336 32812 7364
rect 34422 7352 34428 7364
rect 34480 7392 34486 7404
rect 34480 7364 34928 7392
rect 34480 7352 34486 7364
rect 32214 7284 32220 7336
rect 32272 7284 32278 7336
rect 32766 7284 32772 7336
rect 32824 7284 32830 7336
rect 33226 7284 33232 7336
rect 33284 7324 33290 7336
rect 33689 7327 33747 7333
rect 33689 7324 33701 7327
rect 33284 7296 33701 7324
rect 33284 7284 33290 7296
rect 33689 7293 33701 7296
rect 33735 7324 33747 7327
rect 34238 7324 34244 7336
rect 33735 7296 34244 7324
rect 33735 7293 33747 7296
rect 33689 7287 33747 7293
rect 34238 7284 34244 7296
rect 34296 7284 34302 7336
rect 34900 7333 34928 7364
rect 37458 7352 37464 7404
rect 37516 7392 37522 7404
rect 38197 7395 38255 7401
rect 38197 7392 38209 7395
rect 37516 7364 38209 7392
rect 37516 7352 37522 7364
rect 38197 7361 38209 7364
rect 38243 7361 38255 7395
rect 38197 7355 38255 7361
rect 40034 7352 40040 7404
rect 40092 7352 40098 7404
rect 40126 7352 40132 7404
rect 40184 7392 40190 7404
rect 40880 7401 40908 7432
rect 41322 7420 41328 7432
rect 41380 7460 41386 7472
rect 42260 7460 42288 7491
rect 42426 7488 42432 7500
rect 42484 7488 42490 7540
rect 43530 7488 43536 7540
rect 43588 7528 43594 7540
rect 43809 7531 43867 7537
rect 43809 7528 43821 7531
rect 43588 7500 43821 7528
rect 43588 7488 43594 7500
rect 43809 7497 43821 7500
rect 43855 7528 43867 7531
rect 44729 7531 44787 7537
rect 44729 7528 44741 7531
rect 43855 7500 44741 7528
rect 43855 7497 43867 7500
rect 43809 7491 43867 7497
rect 44729 7497 44741 7500
rect 44775 7497 44787 7531
rect 44729 7491 44787 7497
rect 46014 7488 46020 7540
rect 46072 7488 46078 7540
rect 46293 7531 46351 7537
rect 46293 7497 46305 7531
rect 46339 7528 46351 7531
rect 47670 7528 47676 7540
rect 46339 7500 47676 7528
rect 46339 7497 46351 7500
rect 46293 7491 46351 7497
rect 44821 7463 44879 7469
rect 44821 7460 44833 7463
rect 41380 7420 41414 7460
rect 42260 7432 44833 7460
rect 44821 7429 44833 7432
rect 44867 7429 44879 7463
rect 44821 7423 44879 7429
rect 45922 7420 45928 7472
rect 45980 7420 45986 7472
rect 41138 7401 41144 7404
rect 40865 7395 40923 7401
rect 40865 7392 40877 7395
rect 40184 7364 40877 7392
rect 40184 7352 40190 7364
rect 40865 7361 40877 7364
rect 40911 7361 40923 7395
rect 41132 7392 41144 7401
rect 41099 7364 41144 7392
rect 40865 7355 40923 7361
rect 41132 7355 41144 7364
rect 41138 7352 41144 7355
rect 41196 7352 41202 7404
rect 41386 7392 41414 7420
rect 42426 7392 42432 7404
rect 41386 7364 42432 7392
rect 42426 7352 42432 7364
rect 42484 7352 42490 7404
rect 42518 7352 42524 7404
rect 42576 7392 42582 7404
rect 42685 7395 42743 7401
rect 42685 7392 42697 7395
rect 42576 7364 42697 7392
rect 42576 7352 42582 7364
rect 42685 7361 42697 7364
rect 42731 7361 42743 7395
rect 46032 7392 46060 7488
rect 42685 7355 42743 7361
rect 44928 7364 46060 7392
rect 46155 7429 46213 7435
rect 46155 7395 46167 7429
rect 46201 7395 46213 7429
rect 46400 7401 46428 7500
rect 47670 7488 47676 7500
rect 47728 7488 47734 7540
rect 47765 7531 47823 7537
rect 47765 7497 47777 7531
rect 47811 7528 47823 7531
rect 48314 7528 48320 7540
rect 47811 7500 48320 7528
rect 47811 7497 47823 7500
rect 47765 7491 47823 7497
rect 48314 7488 48320 7500
rect 48372 7488 48378 7540
rect 48406 7488 48412 7540
rect 48464 7488 48470 7540
rect 48590 7488 48596 7540
rect 48648 7488 48654 7540
rect 49142 7488 49148 7540
rect 49200 7528 49206 7540
rect 49697 7531 49755 7537
rect 49697 7528 49709 7531
rect 49200 7500 49709 7528
rect 49200 7488 49206 7500
rect 49697 7497 49709 7500
rect 49743 7497 49755 7531
rect 49697 7491 49755 7497
rect 48130 7420 48136 7472
rect 48188 7420 48194 7472
rect 46155 7392 46213 7395
rect 46385 7395 46443 7401
rect 46155 7389 46244 7392
rect 46156 7364 46244 7389
rect 34885 7327 34943 7333
rect 34885 7293 34897 7327
rect 34931 7293 34943 7327
rect 36357 7327 36415 7333
rect 36357 7324 36369 7327
rect 34885 7287 34943 7293
rect 36280 7296 36369 7324
rect 32784 7228 34008 7256
rect 32784 7188 32812 7228
rect 33980 7200 34008 7228
rect 36280 7200 36308 7296
rect 36357 7293 36369 7296
rect 36403 7293 36415 7327
rect 36357 7287 36415 7293
rect 44361 7259 44419 7265
rect 44361 7225 44373 7259
rect 44407 7256 44419 7259
rect 44928 7256 44956 7364
rect 45005 7327 45063 7333
rect 45005 7293 45017 7327
rect 45051 7324 45063 7327
rect 46216 7324 46244 7364
rect 46385 7361 46397 7395
rect 46431 7361 46443 7395
rect 46385 7355 46443 7361
rect 46661 7395 46719 7401
rect 46661 7361 46673 7395
rect 46707 7361 46719 7395
rect 46661 7355 46719 7361
rect 45051 7296 46244 7324
rect 45051 7293 45063 7296
rect 45005 7287 45063 7293
rect 44407 7228 44956 7256
rect 46216 7256 46244 7296
rect 46676 7324 46704 7355
rect 46750 7352 46756 7404
rect 46808 7392 46814 7404
rect 46845 7395 46903 7401
rect 46845 7392 46857 7395
rect 46808 7364 46857 7392
rect 46808 7352 46814 7364
rect 46845 7361 46857 7364
rect 46891 7361 46903 7395
rect 46845 7355 46903 7361
rect 47949 7395 48007 7401
rect 47949 7361 47961 7395
rect 47995 7392 48007 7395
rect 48038 7392 48044 7404
rect 47995 7364 48044 7392
rect 47995 7361 48007 7364
rect 47949 7355 48007 7361
rect 48038 7352 48044 7364
rect 48096 7352 48102 7404
rect 48225 7395 48283 7401
rect 48225 7361 48237 7395
rect 48271 7392 48283 7395
rect 48424 7392 48452 7488
rect 48271 7364 48452 7392
rect 48608 7392 48636 7488
rect 48961 7463 49019 7469
rect 48961 7429 48973 7463
rect 49007 7460 49019 7463
rect 49421 7463 49479 7469
rect 49421 7460 49433 7463
rect 49007 7432 49433 7460
rect 49007 7429 49019 7432
rect 48961 7423 49019 7429
rect 49421 7429 49433 7432
rect 49467 7429 49479 7463
rect 49421 7423 49479 7429
rect 49510 7420 49516 7472
rect 49568 7420 49574 7472
rect 49510 7417 49568 7420
rect 49237 7395 49295 7401
rect 49237 7392 49249 7395
rect 48608 7364 49249 7392
rect 48271 7361 48283 7364
rect 48225 7355 48283 7361
rect 46676 7296 46888 7324
rect 46676 7256 46704 7296
rect 46216 7228 46704 7256
rect 44407 7225 44419 7228
rect 44361 7219 44419 7225
rect 46860 7200 46888 7296
rect 47762 7284 47768 7336
rect 47820 7324 47826 7336
rect 48317 7327 48375 7333
rect 48317 7324 48329 7327
rect 47820 7296 48329 7324
rect 47820 7284 47826 7296
rect 48317 7293 48329 7296
rect 48363 7293 48375 7327
rect 48424 7324 48452 7364
rect 49237 7361 49249 7364
rect 49283 7361 49295 7395
rect 49510 7383 49522 7417
rect 49556 7383 49568 7417
rect 49510 7377 49568 7383
rect 49605 7395 49663 7401
rect 49237 7355 49295 7361
rect 49605 7361 49617 7395
rect 49651 7361 49663 7395
rect 49605 7355 49663 7361
rect 49620 7324 49648 7355
rect 49694 7352 49700 7404
rect 49752 7392 49758 7404
rect 49789 7395 49847 7401
rect 49789 7392 49801 7395
rect 49752 7364 49801 7392
rect 49752 7352 49758 7364
rect 49789 7361 49801 7364
rect 49835 7361 49847 7395
rect 49789 7355 49847 7361
rect 48424 7296 49648 7324
rect 48317 7287 48375 7293
rect 48332 7256 48360 7287
rect 49786 7256 49792 7268
rect 48332 7228 49792 7256
rect 49786 7216 49792 7228
rect 49844 7216 49850 7268
rect 31036 7160 32812 7188
rect 32858 7148 32864 7200
rect 32916 7188 32922 7200
rect 33045 7191 33103 7197
rect 33045 7188 33057 7191
rect 32916 7160 33057 7188
rect 32916 7148 32922 7160
rect 33045 7157 33057 7160
rect 33091 7157 33103 7191
rect 33045 7151 33103 7157
rect 33962 7148 33968 7200
rect 34020 7148 34026 7200
rect 36262 7148 36268 7200
rect 36320 7148 36326 7200
rect 36998 7148 37004 7200
rect 37056 7148 37062 7200
rect 39942 7148 39948 7200
rect 40000 7148 40006 7200
rect 46106 7148 46112 7200
rect 46164 7148 46170 7200
rect 46474 7148 46480 7200
rect 46532 7148 46538 7200
rect 46658 7148 46664 7200
rect 46716 7148 46722 7200
rect 46842 7148 46848 7200
rect 46900 7148 46906 7200
rect 49050 7148 49056 7200
rect 49108 7148 49114 7200
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 25856 6987 25914 6993
rect 25856 6953 25868 6987
rect 25902 6984 25914 6987
rect 29181 6987 29239 6993
rect 29181 6984 29193 6987
rect 25902 6956 29193 6984
rect 25902 6953 25914 6956
rect 25856 6947 25914 6953
rect 29181 6953 29193 6956
rect 29227 6953 29239 6987
rect 29181 6947 29239 6953
rect 29546 6944 29552 6996
rect 29604 6984 29610 6996
rect 29733 6987 29791 6993
rect 29733 6984 29745 6987
rect 29604 6956 29745 6984
rect 29604 6944 29610 6956
rect 29733 6953 29745 6956
rect 29779 6953 29791 6987
rect 29733 6947 29791 6953
rect 35894 6944 35900 6996
rect 35952 6984 35958 6996
rect 36449 6987 36507 6993
rect 36449 6984 36461 6987
rect 35952 6956 36461 6984
rect 35952 6944 35958 6956
rect 36449 6953 36461 6956
rect 36495 6953 36507 6987
rect 36449 6947 36507 6953
rect 37918 6944 37924 6996
rect 37976 6984 37982 6996
rect 39114 6984 39120 6996
rect 37976 6956 39120 6984
rect 37976 6944 37982 6956
rect 39114 6944 39120 6956
rect 39172 6944 39178 6996
rect 41877 6987 41935 6993
rect 41877 6953 41889 6987
rect 41923 6984 41935 6987
rect 42518 6984 42524 6996
rect 41923 6956 42524 6984
rect 41923 6953 41935 6956
rect 41877 6947 41935 6953
rect 42518 6944 42524 6956
rect 42576 6944 42582 6996
rect 43244 6987 43302 6993
rect 43244 6953 43256 6987
rect 43290 6984 43302 6987
rect 45005 6987 45063 6993
rect 45005 6984 45017 6987
rect 43290 6956 45017 6984
rect 43290 6953 43302 6956
rect 43244 6947 43302 6953
rect 45005 6953 45017 6956
rect 45051 6953 45063 6987
rect 45922 6984 45928 6996
rect 45005 6947 45063 6953
rect 45480 6956 45928 6984
rect 28534 6876 28540 6928
rect 28592 6876 28598 6928
rect 33410 6876 33416 6928
rect 33468 6876 33474 6928
rect 33502 6876 33508 6928
rect 33560 6876 33566 6928
rect 27341 6851 27399 6857
rect 27341 6817 27353 6851
rect 27387 6848 27399 6851
rect 27890 6848 27896 6860
rect 27387 6820 27896 6848
rect 27387 6817 27399 6820
rect 27341 6811 27399 6817
rect 25590 6740 25596 6792
rect 25648 6740 25654 6792
rect 27632 6789 27660 6820
rect 27890 6808 27896 6820
rect 27948 6808 27954 6860
rect 28552 6848 28580 6876
rect 28552 6820 28856 6848
rect 28828 6792 28856 6820
rect 28902 6808 28908 6860
rect 28960 6848 28966 6860
rect 29825 6851 29883 6857
rect 29825 6848 29837 6851
rect 28960 6820 29837 6848
rect 28960 6808 28966 6820
rect 27617 6783 27675 6789
rect 27617 6749 27629 6783
rect 27663 6749 27675 6783
rect 27617 6743 27675 6749
rect 27709 6783 27767 6789
rect 27709 6749 27721 6783
rect 27755 6780 27767 6783
rect 28442 6780 28448 6792
rect 27755 6752 28448 6780
rect 27755 6749 27767 6752
rect 27709 6743 27767 6749
rect 28442 6740 28448 6752
rect 28500 6740 28506 6792
rect 28537 6783 28595 6789
rect 28537 6749 28549 6783
rect 28583 6780 28595 6783
rect 28629 6783 28687 6789
rect 28629 6780 28641 6783
rect 28583 6752 28641 6780
rect 28583 6749 28595 6752
rect 28537 6743 28595 6749
rect 28629 6749 28641 6752
rect 28675 6749 28687 6783
rect 28629 6743 28687 6749
rect 28810 6740 28816 6792
rect 28868 6740 28874 6792
rect 28997 6783 29055 6789
rect 28997 6749 29009 6783
rect 29043 6749 29055 6783
rect 28997 6743 29055 6749
rect 26602 6672 26608 6724
rect 26660 6672 26666 6724
rect 27430 6672 27436 6724
rect 27488 6672 27494 6724
rect 27540 6684 28856 6712
rect 27540 6656 27568 6684
rect 27522 6604 27528 6656
rect 27580 6653 27586 6656
rect 27580 6607 27589 6653
rect 28828 6644 28856 6684
rect 28902 6672 28908 6724
rect 28960 6672 28966 6724
rect 29012 6644 29040 6743
rect 28828 6616 29040 6644
rect 29656 6644 29684 6820
rect 29825 6817 29837 6820
rect 29871 6817 29883 6851
rect 29825 6811 29883 6817
rect 31573 6851 31631 6857
rect 31573 6817 31585 6851
rect 31619 6848 31631 6851
rect 32214 6848 32220 6860
rect 31619 6820 32220 6848
rect 31619 6817 31631 6820
rect 31573 6811 31631 6817
rect 32214 6808 32220 6820
rect 32272 6808 32278 6860
rect 29733 6783 29791 6789
rect 29733 6749 29745 6783
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 29748 6712 29776 6743
rect 31754 6740 31760 6792
rect 31812 6740 31818 6792
rect 32490 6740 32496 6792
rect 32548 6780 32554 6792
rect 33321 6783 33379 6789
rect 33321 6780 33333 6783
rect 32548 6752 33333 6780
rect 32548 6740 32554 6752
rect 33321 6749 33333 6752
rect 33367 6749 33379 6783
rect 33428 6780 33456 6876
rect 33520 6848 33548 6876
rect 33520 6820 33824 6848
rect 33796 6789 33824 6820
rect 34238 6808 34244 6860
rect 34296 6808 34302 6860
rect 35253 6851 35311 6857
rect 35253 6817 35265 6851
rect 35299 6817 35311 6851
rect 37645 6851 37703 6857
rect 35253 6811 35311 6817
rect 37200 6820 37596 6848
rect 33505 6783 33563 6789
rect 33505 6780 33517 6783
rect 33428 6752 33517 6780
rect 33321 6743 33379 6749
rect 33505 6749 33517 6752
rect 33551 6749 33563 6783
rect 33505 6743 33563 6749
rect 33781 6783 33839 6789
rect 33781 6749 33793 6783
rect 33827 6780 33839 6783
rect 34054 6780 34060 6792
rect 33827 6752 34060 6780
rect 33827 6749 33839 6752
rect 33781 6743 33839 6749
rect 34054 6740 34060 6752
rect 34112 6740 34118 6792
rect 34256 6780 34284 6808
rect 35268 6780 35296 6811
rect 37200 6792 37228 6820
rect 34256 6752 35296 6780
rect 36078 6740 36084 6792
rect 36136 6740 36142 6792
rect 36357 6783 36415 6789
rect 36357 6749 36369 6783
rect 36403 6780 36415 6783
rect 36998 6780 37004 6792
rect 36403 6752 37004 6780
rect 36403 6749 36415 6752
rect 36357 6743 36415 6749
rect 36998 6740 37004 6752
rect 37056 6740 37062 6792
rect 37182 6740 37188 6792
rect 37240 6740 37246 6792
rect 37458 6780 37464 6792
rect 37384 6752 37464 6780
rect 33226 6712 33232 6724
rect 29748 6684 33232 6712
rect 33226 6672 33232 6684
rect 33284 6672 33290 6724
rect 35069 6715 35127 6721
rect 35069 6712 35081 6715
rect 34532 6684 35081 6712
rect 34532 6656 34560 6684
rect 35069 6681 35081 6684
rect 35115 6681 35127 6715
rect 36096 6712 36124 6740
rect 37384 6712 37412 6752
rect 37458 6740 37464 6752
rect 37516 6740 37522 6792
rect 37568 6780 37596 6820
rect 37645 6817 37657 6851
rect 37691 6848 37703 6851
rect 39132 6848 39160 6944
rect 39574 6876 39580 6928
rect 39632 6916 39638 6928
rect 39632 6888 40540 6916
rect 39632 6876 39638 6888
rect 37691 6820 38240 6848
rect 39132 6820 40448 6848
rect 37691 6817 37703 6820
rect 37645 6811 37703 6817
rect 38212 6792 38240 6820
rect 37737 6783 37795 6789
rect 37737 6780 37749 6783
rect 37568 6752 37749 6780
rect 37737 6749 37749 6752
rect 37783 6749 37795 6783
rect 37737 6743 37795 6749
rect 38194 6740 38200 6792
rect 38252 6740 38258 6792
rect 38381 6783 38439 6789
rect 38381 6749 38393 6783
rect 38427 6780 38439 6783
rect 39574 6780 39580 6792
rect 38427 6752 39580 6780
rect 38427 6749 38439 6752
rect 38381 6743 38439 6749
rect 39574 6740 39580 6752
rect 39632 6740 39638 6792
rect 39942 6740 39948 6792
rect 40000 6740 40006 6792
rect 40420 6789 40448 6820
rect 40037 6783 40095 6789
rect 40037 6749 40049 6783
rect 40083 6749 40095 6783
rect 40037 6743 40095 6749
rect 40405 6783 40463 6789
rect 40405 6749 40417 6783
rect 40451 6749 40463 6783
rect 40512 6780 40540 6888
rect 42058 6876 42064 6928
rect 42116 6876 42122 6928
rect 40589 6783 40647 6789
rect 40589 6780 40601 6783
rect 40512 6752 40601 6780
rect 40405 6743 40463 6749
rect 40589 6749 40601 6752
rect 40635 6749 40647 6783
rect 40589 6743 40647 6749
rect 41877 6783 41935 6789
rect 41877 6749 41889 6783
rect 41923 6780 41935 6783
rect 42076 6780 42104 6876
rect 42426 6808 42432 6860
rect 42484 6848 42490 6860
rect 42981 6851 43039 6857
rect 42981 6848 42993 6851
rect 42484 6820 42993 6848
rect 42484 6808 42490 6820
rect 42981 6817 42993 6820
rect 43027 6817 43039 6851
rect 42981 6811 43039 6817
rect 44729 6851 44787 6857
rect 44729 6817 44741 6851
rect 44775 6848 44787 6851
rect 45480 6848 45508 6956
rect 45922 6944 45928 6956
rect 45980 6984 45986 6996
rect 48304 6987 48362 6993
rect 45980 6956 46612 6984
rect 45980 6944 45986 6956
rect 46474 6916 46480 6928
rect 44775 6820 45508 6848
rect 45572 6888 46480 6916
rect 44775 6817 44787 6820
rect 44729 6811 44787 6817
rect 41923 6752 42104 6780
rect 41923 6749 41935 6752
rect 41877 6743 41935 6749
rect 36096 6684 37412 6712
rect 40052 6712 40080 6743
rect 42150 6740 42156 6792
rect 42208 6740 42214 6792
rect 42794 6740 42800 6792
rect 42852 6740 42858 6792
rect 45189 6783 45247 6789
rect 45189 6749 45201 6783
rect 45235 6749 45247 6783
rect 45189 6743 45247 6749
rect 45281 6783 45339 6789
rect 45281 6749 45293 6783
rect 45327 6780 45339 6783
rect 45572 6780 45600 6888
rect 46474 6876 46480 6888
rect 46532 6876 46538 6928
rect 45649 6851 45707 6857
rect 45649 6817 45661 6851
rect 45695 6848 45707 6851
rect 46385 6851 46443 6857
rect 46385 6848 46397 6851
rect 45695 6820 46397 6848
rect 45695 6817 45707 6820
rect 45649 6811 45707 6817
rect 46385 6817 46397 6820
rect 46431 6817 46443 6851
rect 46584 6848 46612 6956
rect 48304 6953 48316 6987
rect 48350 6984 48362 6987
rect 49050 6984 49056 6996
rect 48350 6956 49056 6984
rect 48350 6953 48362 6956
rect 48304 6947 48362 6953
rect 49050 6944 49056 6956
rect 49108 6944 49114 6996
rect 49786 6944 49792 6996
rect 49844 6944 49850 6996
rect 46937 6851 46995 6857
rect 46937 6848 46949 6851
rect 46584 6820 46949 6848
rect 46385 6811 46443 6817
rect 46937 6817 46949 6820
rect 46983 6817 46995 6851
rect 46937 6811 46995 6817
rect 45327 6752 45600 6780
rect 45833 6783 45891 6789
rect 45327 6749 45339 6752
rect 45281 6743 45339 6749
rect 45833 6749 45845 6783
rect 45879 6780 45891 6783
rect 45922 6780 45928 6792
rect 45879 6752 45928 6780
rect 45879 6749 45891 6752
rect 45833 6743 45891 6749
rect 40497 6715 40555 6721
rect 40497 6712 40509 6715
rect 40052 6684 40509 6712
rect 35069 6675 35127 6681
rect 40497 6681 40509 6684
rect 40543 6681 40555 6715
rect 40497 6675 40555 6681
rect 42061 6715 42119 6721
rect 42061 6681 42073 6715
rect 42107 6712 42119 6715
rect 42812 6712 42840 6740
rect 42107 6684 42840 6712
rect 42107 6681 42119 6684
rect 42061 6675 42119 6681
rect 29730 6644 29736 6656
rect 29656 6616 29736 6644
rect 27580 6604 27586 6607
rect 29730 6604 29736 6616
rect 29788 6604 29794 6656
rect 30098 6604 30104 6656
rect 30156 6604 30162 6656
rect 30834 6604 30840 6656
rect 30892 6644 30898 6656
rect 31941 6647 31999 6653
rect 31941 6644 31953 6647
rect 30892 6616 31953 6644
rect 30892 6604 30898 6616
rect 31941 6613 31953 6616
rect 31987 6644 31999 6647
rect 32582 6644 32588 6656
rect 31987 6616 32588 6644
rect 31987 6613 31999 6616
rect 31941 6607 31999 6613
rect 32582 6604 32588 6616
rect 32640 6604 32646 6656
rect 33686 6604 33692 6656
rect 33744 6604 33750 6656
rect 33778 6604 33784 6656
rect 33836 6644 33842 6656
rect 33873 6647 33931 6653
rect 33873 6644 33885 6647
rect 33836 6616 33885 6644
rect 33836 6604 33842 6616
rect 33873 6613 33885 6616
rect 33919 6613 33931 6647
rect 33873 6607 33931 6613
rect 34514 6604 34520 6656
rect 34572 6604 34578 6656
rect 34698 6604 34704 6656
rect 34756 6604 34762 6656
rect 35161 6647 35219 6653
rect 35161 6613 35173 6647
rect 35207 6644 35219 6647
rect 35618 6644 35624 6656
rect 35207 6616 35624 6644
rect 35207 6613 35219 6616
rect 35161 6607 35219 6613
rect 35618 6604 35624 6616
rect 35676 6604 35682 6656
rect 37274 6604 37280 6656
rect 37332 6604 37338 6656
rect 38654 6604 38660 6656
rect 38712 6644 38718 6656
rect 38933 6647 38991 6653
rect 38933 6644 38945 6647
rect 38712 6616 38945 6644
rect 38712 6604 38718 6616
rect 38933 6613 38945 6616
rect 38979 6613 38991 6647
rect 38933 6607 38991 6613
rect 40218 6604 40224 6656
rect 40276 6604 40282 6656
rect 40512 6644 40540 6675
rect 44266 6672 44272 6724
rect 44324 6672 44330 6724
rect 40586 6644 40592 6656
rect 40512 6616 40592 6644
rect 40586 6604 40592 6616
rect 40644 6604 40650 6656
rect 45204 6644 45232 6743
rect 45922 6740 45928 6752
rect 45980 6740 45986 6792
rect 46106 6740 46112 6792
rect 46164 6780 46170 6792
rect 46661 6783 46719 6789
rect 46661 6780 46673 6783
rect 46164 6752 46673 6780
rect 46164 6740 46170 6752
rect 46661 6749 46673 6752
rect 46707 6749 46719 6783
rect 46661 6743 46719 6749
rect 46750 6740 46756 6792
rect 46808 6740 46814 6792
rect 46845 6783 46903 6789
rect 46845 6749 46857 6783
rect 46891 6749 46903 6783
rect 46845 6743 46903 6749
rect 45370 6672 45376 6724
rect 45428 6672 45434 6724
rect 45511 6715 45569 6721
rect 45511 6681 45523 6715
rect 45557 6712 45569 6715
rect 46014 6712 46020 6724
rect 45557 6684 46020 6712
rect 45557 6681 45569 6684
rect 45511 6675 45569 6681
rect 46014 6672 46020 6684
rect 46072 6672 46078 6724
rect 46198 6672 46204 6724
rect 46256 6712 46262 6724
rect 46860 6712 46888 6743
rect 47026 6740 47032 6792
rect 47084 6780 47090 6792
rect 48041 6783 48099 6789
rect 48041 6780 48053 6783
rect 47084 6752 48053 6780
rect 47084 6740 47090 6752
rect 48041 6749 48053 6752
rect 48087 6749 48099 6783
rect 48041 6743 48099 6749
rect 46256 6684 46888 6712
rect 46256 6672 46262 6684
rect 48774 6672 48780 6724
rect 48832 6672 48838 6724
rect 46477 6647 46535 6653
rect 46477 6644 46489 6647
rect 45204 6616 46489 6644
rect 46477 6613 46489 6616
rect 46523 6613 46535 6647
rect 46477 6607 46535 6613
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 26602 6400 26608 6452
rect 26660 6440 26666 6452
rect 26697 6443 26755 6449
rect 26697 6440 26709 6443
rect 26660 6412 26709 6440
rect 26660 6400 26666 6412
rect 26697 6409 26709 6412
rect 26743 6409 26755 6443
rect 26697 6403 26755 6409
rect 27522 6400 27528 6452
rect 27580 6400 27586 6452
rect 28626 6400 28632 6452
rect 28684 6400 28690 6452
rect 28810 6400 28816 6452
rect 28868 6400 28874 6452
rect 28994 6400 29000 6452
rect 29052 6440 29058 6452
rect 29273 6443 29331 6449
rect 29273 6440 29285 6443
rect 29052 6412 29285 6440
rect 29052 6400 29058 6412
rect 29273 6409 29285 6412
rect 29319 6409 29331 6443
rect 29273 6403 29331 6409
rect 29822 6400 29828 6452
rect 29880 6400 29886 6452
rect 30098 6400 30104 6452
rect 30156 6400 30162 6452
rect 31754 6440 31760 6452
rect 31496 6412 31760 6440
rect 27540 6372 27568 6400
rect 28445 6375 28503 6381
rect 28445 6372 28457 6375
rect 27540 6344 28457 6372
rect 28445 6341 28457 6344
rect 28491 6341 28503 6375
rect 28644 6372 28672 6400
rect 28905 6375 28963 6381
rect 28905 6372 28917 6375
rect 28644 6344 28917 6372
rect 28445 6335 28503 6341
rect 28905 6341 28917 6344
rect 28951 6341 28963 6375
rect 29105 6375 29163 6381
rect 29105 6372 29117 6375
rect 28905 6335 28963 6341
rect 29012 6344 29117 6372
rect 26605 6307 26663 6313
rect 26605 6273 26617 6307
rect 26651 6304 26663 6307
rect 26970 6304 26976 6316
rect 26651 6276 26976 6304
rect 26651 6273 26663 6276
rect 26605 6267 26663 6273
rect 26970 6264 26976 6276
rect 27028 6264 27034 6316
rect 27890 6264 27896 6316
rect 27948 6264 27954 6316
rect 28350 6264 28356 6316
rect 28408 6304 28414 6316
rect 28629 6307 28687 6313
rect 28629 6304 28641 6307
rect 28408 6276 28641 6304
rect 28408 6264 28414 6276
rect 28629 6273 28641 6276
rect 28675 6304 28687 6307
rect 28810 6304 28816 6316
rect 28675 6276 28816 6304
rect 28675 6273 28687 6276
rect 28629 6267 28687 6273
rect 28810 6264 28816 6276
rect 28868 6264 28874 6316
rect 29012 6304 29040 6344
rect 29105 6341 29117 6344
rect 29151 6341 29163 6375
rect 29840 6372 29868 6400
rect 30009 6375 30067 6381
rect 30009 6372 30021 6375
rect 29105 6335 29163 6341
rect 29472 6344 29776 6372
rect 29840 6344 30021 6372
rect 29472 6304 29500 6344
rect 28920 6276 29040 6304
rect 29104 6276 29500 6304
rect 27908 6100 27936 6264
rect 28920 6248 28948 6276
rect 28442 6196 28448 6248
rect 28500 6236 28506 6248
rect 28902 6236 28908 6248
rect 28500 6208 28908 6236
rect 28500 6196 28506 6208
rect 28902 6196 28908 6208
rect 28960 6196 28966 6248
rect 27982 6128 27988 6180
rect 28040 6168 28046 6180
rect 28718 6168 28724 6180
rect 28040 6140 28724 6168
rect 28040 6128 28046 6140
rect 28718 6128 28724 6140
rect 28776 6128 28782 6180
rect 29104 6168 29132 6276
rect 29546 6264 29552 6316
rect 29604 6264 29610 6316
rect 29641 6307 29699 6313
rect 29641 6273 29653 6307
rect 29687 6273 29699 6307
rect 29748 6304 29776 6344
rect 30009 6341 30021 6344
rect 30055 6341 30067 6375
rect 30116 6372 30144 6400
rect 30116 6344 30420 6372
rect 30009 6335 30067 6341
rect 29825 6307 29883 6313
rect 29825 6304 29837 6307
rect 29748 6276 29837 6304
rect 29641 6267 29699 6273
rect 29825 6273 29837 6276
rect 29871 6273 29883 6307
rect 29825 6267 29883 6273
rect 29656 6236 29684 6267
rect 29914 6264 29920 6316
rect 29972 6304 29978 6316
rect 30392 6313 30420 6344
rect 30576 6344 30972 6372
rect 30576 6316 30604 6344
rect 30377 6307 30435 6313
rect 29972 6276 30328 6304
rect 29972 6264 29978 6276
rect 30006 6236 30012 6248
rect 29656 6208 30012 6236
rect 30006 6196 30012 6208
rect 30064 6196 30070 6248
rect 30300 6245 30328 6276
rect 30377 6273 30389 6307
rect 30423 6273 30435 6307
rect 30377 6267 30435 6273
rect 30466 6264 30472 6316
rect 30524 6264 30530 6316
rect 30558 6264 30564 6316
rect 30616 6264 30622 6316
rect 30650 6264 30656 6316
rect 30708 6264 30714 6316
rect 30944 6313 30972 6344
rect 30929 6307 30987 6313
rect 30929 6273 30941 6307
rect 30975 6273 30987 6307
rect 30929 6267 30987 6273
rect 30285 6239 30343 6245
rect 30285 6205 30297 6239
rect 30331 6205 30343 6239
rect 31496 6236 31524 6412
rect 31754 6400 31760 6412
rect 31812 6400 31818 6452
rect 36081 6443 36139 6449
rect 36081 6409 36093 6443
rect 36127 6440 36139 6443
rect 36127 6412 36860 6440
rect 36127 6409 36139 6412
rect 36081 6403 36139 6409
rect 31662 6332 31668 6384
rect 31720 6332 31726 6384
rect 33778 6332 33784 6384
rect 33836 6332 33842 6384
rect 36262 6372 36268 6384
rect 35728 6344 36268 6372
rect 31573 6307 31631 6313
rect 31573 6273 31585 6307
rect 31619 6304 31631 6307
rect 31680 6304 31708 6332
rect 35728 6313 35756 6344
rect 36262 6332 36268 6344
rect 36320 6332 36326 6384
rect 31619 6276 31708 6304
rect 31757 6307 31815 6313
rect 31619 6273 31631 6276
rect 31573 6267 31631 6273
rect 31757 6273 31769 6307
rect 31803 6273 31815 6307
rect 31757 6267 31815 6273
rect 35529 6307 35587 6313
rect 35529 6273 35541 6307
rect 35575 6273 35587 6307
rect 35529 6267 35587 6273
rect 35713 6307 35771 6313
rect 35713 6273 35725 6307
rect 35759 6273 35771 6307
rect 35713 6267 35771 6273
rect 31665 6239 31723 6245
rect 31665 6236 31677 6239
rect 30285 6199 30343 6205
rect 30392 6208 31677 6236
rect 30193 6171 30251 6177
rect 30193 6168 30205 6171
rect 29104 6140 30205 6168
rect 29104 6109 29132 6140
rect 30193 6137 30205 6140
rect 30239 6137 30251 6171
rect 30392 6168 30420 6208
rect 31665 6205 31677 6208
rect 31711 6205 31723 6239
rect 31665 6199 31723 6205
rect 31772 6168 31800 6267
rect 32766 6196 32772 6248
rect 32824 6196 32830 6248
rect 33042 6196 33048 6248
rect 33100 6196 33106 6248
rect 32490 6168 32496 6180
rect 30193 6131 30251 6137
rect 30300 6140 30420 6168
rect 31588 6140 32496 6168
rect 30300 6112 30328 6140
rect 31588 6112 31616 6140
rect 32490 6128 32496 6140
rect 32548 6128 32554 6180
rect 29089 6103 29147 6109
rect 29089 6100 29101 6103
rect 27908 6072 29101 6100
rect 29089 6069 29101 6072
rect 29135 6069 29147 6103
rect 29089 6063 29147 6069
rect 29365 6103 29423 6109
rect 29365 6069 29377 6103
rect 29411 6100 29423 6103
rect 30098 6100 30104 6112
rect 29411 6072 30104 6100
rect 29411 6069 29423 6072
rect 29365 6063 29423 6069
rect 30098 6060 30104 6072
rect 30156 6060 30162 6112
rect 30282 6060 30288 6112
rect 30340 6060 30346 6112
rect 31018 6060 31024 6112
rect 31076 6060 31082 6112
rect 31570 6060 31576 6112
rect 31628 6060 31634 6112
rect 34514 6060 34520 6112
rect 34572 6060 34578 6112
rect 35544 6100 35572 6267
rect 35802 6264 35808 6316
rect 35860 6264 35866 6316
rect 35897 6307 35955 6313
rect 35897 6273 35909 6307
rect 35943 6304 35955 6307
rect 35943 6276 36216 6304
rect 35943 6273 35955 6276
rect 35897 6267 35955 6273
rect 36188 6248 36216 6276
rect 36354 6264 36360 6316
rect 36412 6264 36418 6316
rect 36832 6313 36860 6412
rect 38838 6400 38844 6452
rect 38896 6400 38902 6452
rect 39114 6400 39120 6452
rect 39172 6400 39178 6452
rect 40773 6443 40831 6449
rect 40773 6409 40785 6443
rect 40819 6440 40831 6443
rect 41506 6440 41512 6452
rect 40819 6412 41512 6440
rect 40819 6409 40831 6412
rect 40773 6403 40831 6409
rect 41506 6400 41512 6412
rect 41564 6400 41570 6452
rect 44266 6400 44272 6452
rect 44324 6400 44330 6452
rect 45925 6443 45983 6449
rect 45925 6409 45937 6443
rect 45971 6440 45983 6443
rect 45971 6412 46612 6440
rect 45971 6409 45983 6412
rect 45925 6403 45983 6409
rect 38197 6375 38255 6381
rect 38197 6341 38209 6375
rect 38243 6372 38255 6375
rect 38286 6372 38292 6384
rect 38243 6344 38292 6372
rect 38243 6341 38255 6344
rect 38197 6335 38255 6341
rect 38286 6332 38292 6344
rect 38344 6332 38350 6384
rect 40497 6375 40555 6381
rect 40497 6341 40509 6375
rect 40543 6372 40555 6375
rect 41141 6375 41199 6381
rect 41141 6372 41153 6375
rect 40543 6344 41153 6372
rect 40543 6341 40555 6344
rect 40497 6335 40555 6341
rect 41141 6341 41153 6344
rect 41187 6341 41199 6375
rect 41141 6335 41199 6341
rect 43898 6332 43904 6384
rect 43956 6372 43962 6384
rect 45557 6375 45615 6381
rect 43956 6344 44220 6372
rect 43956 6332 43962 6344
rect 36450 6307 36508 6313
rect 36450 6273 36462 6307
rect 36496 6273 36508 6307
rect 36450 6267 36508 6273
rect 36633 6307 36691 6313
rect 36633 6273 36645 6307
rect 36679 6273 36691 6307
rect 36633 6267 36691 6273
rect 36725 6307 36783 6313
rect 36725 6273 36737 6307
rect 36771 6273 36783 6307
rect 36725 6267 36783 6273
rect 36822 6307 36880 6313
rect 36822 6273 36834 6307
rect 36868 6273 36880 6307
rect 36822 6267 36880 6273
rect 36078 6196 36084 6248
rect 36136 6196 36142 6248
rect 36170 6196 36176 6248
rect 36228 6236 36234 6248
rect 36464 6236 36492 6267
rect 36648 6236 36676 6267
rect 36228 6208 36492 6236
rect 36556 6208 36676 6236
rect 36740 6236 36768 6267
rect 37090 6264 37096 6316
rect 37148 6264 37154 6316
rect 37366 6264 37372 6316
rect 37424 6304 37430 6316
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 37424 6276 37473 6304
rect 37424 6264 37430 6276
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 38657 6307 38715 6313
rect 38657 6273 38669 6307
rect 38703 6273 38715 6307
rect 38657 6267 38715 6273
rect 37108 6236 37136 6264
rect 36740 6208 37136 6236
rect 37553 6239 37611 6245
rect 36228 6196 36234 6208
rect 35621 6171 35679 6177
rect 35621 6137 35633 6171
rect 35667 6168 35679 6171
rect 36556 6168 36584 6208
rect 35667 6140 36584 6168
rect 35667 6137 35679 6140
rect 35621 6131 35679 6137
rect 36740 6100 36768 6208
rect 37553 6205 37565 6239
rect 37599 6236 37611 6239
rect 38286 6236 38292 6248
rect 37599 6208 38292 6236
rect 37599 6205 37611 6208
rect 37553 6199 37611 6205
rect 38286 6196 38292 6208
rect 38344 6236 38350 6248
rect 38473 6239 38531 6245
rect 38473 6236 38485 6239
rect 38344 6208 38485 6236
rect 38344 6196 38350 6208
rect 38473 6205 38485 6208
rect 38519 6205 38531 6239
rect 38672 6236 38700 6267
rect 38930 6264 38936 6316
rect 38988 6264 38994 6316
rect 39298 6264 39304 6316
rect 39356 6264 39362 6316
rect 40402 6264 40408 6316
rect 40460 6264 40466 6316
rect 40586 6264 40592 6316
rect 40644 6264 40650 6316
rect 44192 6313 44220 6344
rect 45557 6341 45569 6375
rect 45603 6372 45615 6375
rect 46106 6372 46112 6384
rect 45603 6344 46112 6372
rect 45603 6341 45615 6344
rect 45557 6335 45615 6341
rect 46106 6332 46112 6344
rect 46164 6332 46170 6384
rect 46198 6332 46204 6384
rect 46256 6372 46262 6384
rect 46385 6375 46443 6381
rect 46385 6372 46397 6375
rect 46256 6344 46397 6372
rect 46256 6332 46262 6344
rect 46385 6341 46397 6344
rect 46431 6341 46443 6375
rect 46385 6335 46443 6341
rect 44177 6307 44235 6313
rect 44177 6273 44189 6307
rect 44223 6273 44235 6307
rect 44177 6267 44235 6273
rect 45741 6307 45799 6313
rect 45741 6273 45753 6307
rect 45787 6273 45799 6307
rect 45741 6267 45799 6273
rect 46017 6307 46075 6313
rect 46017 6273 46029 6307
rect 46063 6304 46075 6307
rect 46124 6304 46152 6332
rect 46584 6316 46612 6412
rect 48774 6400 48780 6452
rect 48832 6400 48838 6452
rect 46658 6332 46664 6384
rect 46716 6372 46722 6384
rect 46753 6375 46811 6381
rect 46753 6372 46765 6375
rect 46716 6344 46765 6372
rect 46716 6332 46722 6344
rect 46753 6341 46765 6344
rect 46799 6341 46811 6375
rect 46753 6335 46811 6341
rect 46845 6375 46903 6381
rect 46845 6341 46857 6375
rect 46891 6372 46903 6375
rect 48593 6375 48651 6381
rect 48593 6372 48605 6375
rect 46891 6344 48605 6372
rect 46891 6341 46903 6344
rect 46845 6335 46903 6341
rect 48593 6341 48605 6344
rect 48639 6341 48651 6375
rect 48593 6335 48651 6341
rect 46063 6276 46152 6304
rect 46477 6307 46535 6313
rect 46063 6273 46075 6276
rect 46017 6267 46075 6273
rect 46477 6273 46489 6307
rect 46523 6273 46535 6307
rect 46477 6267 46535 6273
rect 39316 6236 39344 6264
rect 38672 6208 39344 6236
rect 38473 6199 38531 6205
rect 41230 6196 41236 6248
rect 41288 6196 41294 6248
rect 41414 6196 41420 6248
rect 41472 6196 41478 6248
rect 45756 6236 45784 6267
rect 45830 6236 45836 6248
rect 45756 6208 45836 6236
rect 45830 6196 45836 6208
rect 45888 6236 45894 6248
rect 46492 6236 46520 6267
rect 46566 6264 46572 6316
rect 46624 6264 46630 6316
rect 46937 6307 46995 6313
rect 46937 6273 46949 6307
rect 46983 6304 46995 6307
rect 47946 6304 47952 6316
rect 46983 6276 47952 6304
rect 46983 6273 46995 6276
rect 46937 6267 46995 6273
rect 46750 6236 46756 6248
rect 45888 6208 46756 6236
rect 45888 6196 45894 6208
rect 46750 6196 46756 6208
rect 46808 6196 46814 6248
rect 46014 6128 46020 6180
rect 46072 6168 46078 6180
rect 46566 6168 46572 6180
rect 46072 6140 46572 6168
rect 46072 6128 46078 6140
rect 46566 6128 46572 6140
rect 46624 6168 46630 6180
rect 46952 6168 46980 6267
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 48314 6264 48320 6316
rect 48372 6304 48378 6316
rect 48685 6307 48743 6313
rect 48685 6304 48697 6307
rect 48372 6276 48697 6304
rect 48372 6264 48378 6276
rect 48685 6273 48697 6276
rect 48731 6273 48743 6307
rect 48685 6267 48743 6273
rect 48041 6239 48099 6245
rect 48041 6205 48053 6239
rect 48087 6236 48099 6239
rect 48087 6208 48912 6236
rect 48087 6205 48099 6208
rect 48041 6199 48099 6205
rect 46624 6140 46980 6168
rect 46624 6128 46630 6140
rect 48884 6112 48912 6208
rect 68462 6128 68468 6180
rect 68520 6128 68526 6180
rect 35544 6072 36768 6100
rect 36998 6060 37004 6112
rect 37056 6060 37062 6112
rect 37826 6060 37832 6112
rect 37884 6060 37890 6112
rect 38562 6060 38568 6112
rect 38620 6100 38626 6112
rect 40862 6100 40868 6112
rect 38620 6072 40868 6100
rect 38620 6060 38626 6072
rect 40862 6060 40868 6072
rect 40920 6060 40926 6112
rect 46198 6060 46204 6112
rect 46256 6060 46262 6112
rect 47121 6103 47179 6109
rect 47121 6069 47133 6103
rect 47167 6100 47179 6103
rect 47394 6100 47400 6112
rect 47167 6072 47400 6100
rect 47167 6069 47179 6072
rect 47121 6063 47179 6069
rect 47394 6060 47400 6072
rect 47452 6060 47458 6112
rect 48866 6060 48872 6112
rect 48924 6060 48930 6112
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 27430 5856 27436 5908
rect 27488 5856 27494 5908
rect 29546 5856 29552 5908
rect 29604 5896 29610 5908
rect 29641 5899 29699 5905
rect 29641 5896 29653 5899
rect 29604 5868 29653 5896
rect 29604 5856 29610 5868
rect 29641 5865 29653 5868
rect 29687 5865 29699 5899
rect 30282 5896 30288 5908
rect 29641 5859 29699 5865
rect 29932 5868 30288 5896
rect 27448 5828 27476 5856
rect 29932 5828 29960 5868
rect 30282 5856 30288 5868
rect 30340 5856 30346 5908
rect 30374 5856 30380 5908
rect 30432 5856 30438 5908
rect 31297 5899 31355 5905
rect 30668 5868 31156 5896
rect 27448 5800 29960 5828
rect 30009 5831 30067 5837
rect 27157 5763 27215 5769
rect 27157 5729 27169 5763
rect 27203 5760 27215 5763
rect 27893 5763 27951 5769
rect 27893 5760 27905 5763
rect 27203 5732 27905 5760
rect 27203 5729 27215 5732
rect 27157 5723 27215 5729
rect 27893 5729 27905 5732
rect 27939 5760 27951 5763
rect 27982 5760 27988 5772
rect 27939 5732 27988 5760
rect 27939 5729 27951 5732
rect 27893 5723 27951 5729
rect 27982 5720 27988 5732
rect 28040 5720 28046 5772
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5661 25467 5695
rect 25409 5655 25467 5661
rect 25424 5624 25452 5655
rect 28074 5652 28080 5704
rect 28132 5652 28138 5704
rect 28276 5701 28304 5800
rect 30009 5797 30021 5831
rect 30055 5828 30067 5831
rect 30668 5828 30696 5868
rect 30055 5800 30696 5828
rect 30055 5797 30067 5800
rect 30009 5791 30067 5797
rect 28552 5732 29868 5760
rect 28552 5704 28580 5732
rect 29840 5704 29868 5732
rect 29914 5720 29920 5772
rect 29972 5720 29978 5772
rect 30558 5720 30564 5772
rect 30616 5720 30622 5772
rect 30742 5720 30748 5772
rect 30800 5720 30806 5772
rect 31128 5769 31156 5868
rect 31297 5865 31309 5899
rect 31343 5896 31355 5899
rect 31938 5896 31944 5908
rect 31343 5868 31944 5896
rect 31343 5865 31355 5868
rect 31297 5859 31355 5865
rect 31938 5856 31944 5868
rect 31996 5856 32002 5908
rect 32416 5868 32996 5896
rect 31113 5763 31171 5769
rect 31113 5729 31125 5763
rect 31159 5729 31171 5763
rect 31113 5723 31171 5729
rect 31662 5720 31668 5772
rect 31720 5760 31726 5772
rect 32416 5760 32444 5868
rect 31720 5732 32444 5760
rect 32968 5760 32996 5868
rect 33042 5856 33048 5908
rect 33100 5856 33106 5908
rect 33413 5899 33471 5905
rect 33413 5865 33425 5899
rect 33459 5896 33471 5899
rect 33686 5896 33692 5908
rect 33459 5868 33692 5896
rect 33459 5865 33471 5868
rect 33413 5859 33471 5865
rect 33686 5856 33692 5868
rect 33744 5856 33750 5908
rect 36170 5856 36176 5908
rect 36228 5856 36234 5908
rect 36998 5856 37004 5908
rect 37056 5856 37062 5908
rect 37274 5856 37280 5908
rect 37332 5856 37338 5908
rect 37458 5856 37464 5908
rect 37516 5896 37522 5908
rect 37829 5899 37887 5905
rect 37829 5896 37841 5899
rect 37516 5868 37841 5896
rect 37516 5856 37522 5868
rect 37829 5865 37841 5868
rect 37875 5865 37887 5899
rect 38562 5896 38568 5908
rect 37829 5859 37887 5865
rect 38212 5868 38568 5896
rect 33505 5763 33563 5769
rect 32968 5732 33272 5760
rect 31720 5720 31726 5732
rect 28261 5695 28319 5701
rect 28261 5661 28273 5695
rect 28307 5661 28319 5695
rect 28261 5655 28319 5661
rect 28353 5695 28411 5701
rect 28353 5661 28365 5695
rect 28399 5661 28411 5695
rect 28353 5655 28411 5661
rect 25590 5624 25596 5636
rect 25424 5596 25596 5624
rect 25590 5584 25596 5596
rect 25648 5584 25654 5636
rect 25682 5584 25688 5636
rect 25740 5584 25746 5636
rect 26418 5584 26424 5636
rect 26476 5584 26482 5636
rect 27617 5627 27675 5633
rect 27617 5593 27629 5627
rect 27663 5624 27675 5627
rect 28169 5627 28227 5633
rect 28169 5624 28181 5627
rect 27663 5596 28181 5624
rect 27663 5593 27675 5596
rect 27617 5587 27675 5593
rect 28169 5593 28181 5596
rect 28215 5593 28227 5627
rect 28169 5587 28227 5593
rect 27246 5516 27252 5568
rect 27304 5516 27310 5568
rect 27706 5516 27712 5568
rect 27764 5516 27770 5568
rect 28368 5556 28396 5655
rect 28534 5652 28540 5704
rect 28592 5652 28598 5704
rect 28626 5652 28632 5704
rect 28684 5652 28690 5704
rect 29549 5695 29607 5701
rect 29549 5661 29561 5695
rect 29595 5661 29607 5695
rect 29549 5655 29607 5661
rect 28644 5624 28672 5652
rect 29564 5624 29592 5655
rect 29822 5652 29828 5704
rect 29880 5652 29886 5704
rect 30006 5652 30012 5704
rect 30064 5652 30070 5704
rect 30098 5652 30104 5704
rect 30156 5652 30162 5704
rect 30374 5652 30380 5704
rect 30432 5692 30438 5704
rect 30653 5695 30711 5701
rect 30653 5692 30665 5695
rect 30432 5664 30665 5692
rect 30432 5652 30438 5664
rect 30653 5661 30665 5664
rect 30699 5661 30711 5695
rect 30653 5655 30711 5661
rect 30834 5652 30840 5704
rect 30892 5652 30898 5704
rect 31297 5695 31355 5701
rect 31297 5661 31309 5695
rect 31343 5661 31355 5695
rect 31570 5692 31576 5704
rect 31297 5655 31355 5661
rect 31404 5664 31576 5692
rect 30024 5624 30052 5652
rect 28644 5596 28994 5624
rect 29564 5596 30052 5624
rect 30116 5624 30144 5652
rect 31021 5627 31079 5633
rect 31021 5624 31033 5627
rect 30116 5596 31033 5624
rect 28442 5556 28448 5568
rect 28368 5528 28448 5556
rect 28442 5516 28448 5528
rect 28500 5516 28506 5568
rect 28537 5559 28595 5565
rect 28537 5525 28549 5559
rect 28583 5556 28595 5559
rect 28810 5556 28816 5568
rect 28583 5528 28816 5556
rect 28583 5525 28595 5528
rect 28537 5519 28595 5525
rect 28810 5516 28816 5528
rect 28868 5516 28874 5568
rect 28966 5556 28994 5596
rect 31021 5593 31033 5596
rect 31067 5593 31079 5627
rect 31021 5587 31079 5593
rect 31202 5584 31208 5636
rect 31260 5624 31266 5636
rect 31312 5624 31340 5655
rect 31260 5596 31340 5624
rect 31260 5584 31266 5596
rect 31404 5556 31432 5664
rect 31570 5652 31576 5664
rect 31628 5652 31634 5704
rect 31680 5692 31708 5720
rect 31757 5695 31815 5701
rect 31757 5692 31769 5695
rect 31680 5664 31769 5692
rect 31757 5661 31769 5664
rect 31803 5661 31815 5695
rect 31757 5655 31815 5661
rect 31938 5652 31944 5704
rect 31996 5652 32002 5704
rect 32306 5652 32312 5704
rect 32364 5652 32370 5704
rect 32490 5652 32496 5704
rect 32548 5652 32554 5704
rect 32582 5652 32588 5704
rect 32640 5701 32646 5704
rect 32640 5695 32669 5701
rect 32657 5661 32669 5695
rect 32640 5655 32669 5661
rect 32769 5695 32827 5701
rect 32769 5661 32781 5695
rect 32815 5692 32827 5695
rect 33134 5692 33140 5704
rect 32815 5664 33140 5692
rect 32815 5661 32827 5664
rect 32769 5655 32827 5661
rect 32640 5652 32646 5655
rect 33134 5652 33140 5664
rect 33192 5652 33198 5704
rect 33244 5701 33272 5732
rect 33505 5729 33517 5763
rect 33551 5760 33563 5763
rect 33689 5763 33747 5769
rect 33689 5760 33701 5763
rect 33551 5732 33701 5760
rect 33551 5729 33563 5732
rect 33505 5723 33563 5729
rect 33689 5729 33701 5732
rect 33735 5729 33747 5763
rect 33689 5723 33747 5729
rect 33229 5695 33287 5701
rect 33229 5661 33241 5695
rect 33275 5661 33287 5695
rect 33229 5655 33287 5661
rect 33410 5652 33416 5704
rect 33468 5692 33474 5704
rect 33597 5695 33655 5701
rect 33597 5692 33609 5695
rect 33468 5664 33609 5692
rect 33468 5652 33474 5664
rect 33597 5661 33609 5664
rect 33643 5661 33655 5695
rect 33597 5655 33655 5661
rect 33781 5695 33839 5701
rect 33781 5661 33793 5695
rect 33827 5692 33839 5695
rect 34514 5692 34520 5704
rect 33827 5664 34520 5692
rect 33827 5661 33839 5664
rect 33781 5655 33839 5661
rect 31956 5624 31984 5652
rect 32401 5627 32459 5633
rect 32401 5624 32413 5627
rect 31956 5596 32413 5624
rect 32401 5593 32413 5596
rect 32447 5593 32459 5627
rect 32508 5624 32536 5652
rect 33796 5624 33824 5655
rect 34514 5652 34520 5664
rect 34572 5652 34578 5704
rect 36081 5695 36139 5701
rect 36081 5661 36093 5695
rect 36127 5692 36139 5695
rect 36357 5695 36415 5701
rect 36127 5664 36216 5692
rect 36127 5661 36139 5664
rect 36081 5655 36139 5661
rect 32508 5596 33824 5624
rect 32401 5587 32459 5593
rect 36188 5568 36216 5664
rect 36357 5661 36369 5695
rect 36403 5692 36415 5695
rect 37016 5692 37044 5856
rect 37090 5788 37096 5840
rect 37148 5828 37154 5840
rect 37148 5800 37964 5828
rect 37148 5788 37154 5800
rect 37384 5769 37412 5800
rect 37369 5763 37427 5769
rect 37369 5729 37381 5763
rect 37415 5760 37427 5763
rect 37415 5732 37449 5760
rect 37415 5729 37427 5732
rect 37369 5723 37427 5729
rect 37734 5720 37740 5772
rect 37792 5720 37798 5772
rect 37826 5720 37832 5772
rect 37884 5720 37890 5772
rect 37093 5695 37151 5701
rect 37093 5692 37105 5695
rect 36403 5664 36860 5692
rect 37016 5664 37105 5692
rect 36403 5661 36415 5664
rect 36357 5655 36415 5661
rect 36832 5568 36860 5664
rect 37093 5661 37105 5664
rect 37139 5661 37151 5695
rect 37093 5655 37151 5661
rect 36909 5627 36967 5633
rect 36909 5593 36921 5627
rect 36955 5624 36967 5627
rect 37752 5624 37780 5720
rect 37844 5633 37872 5720
rect 36955 5596 37780 5624
rect 37829 5627 37887 5633
rect 36955 5593 36967 5596
rect 36909 5587 36967 5593
rect 37829 5593 37841 5627
rect 37875 5593 37887 5627
rect 37936 5624 37964 5800
rect 38013 5763 38071 5769
rect 38013 5729 38025 5763
rect 38059 5760 38071 5763
rect 38212 5760 38240 5868
rect 38562 5856 38568 5868
rect 38620 5856 38626 5908
rect 38841 5899 38899 5905
rect 38841 5865 38853 5899
rect 38887 5865 38899 5899
rect 38841 5859 38899 5865
rect 38289 5831 38347 5837
rect 38289 5797 38301 5831
rect 38335 5797 38347 5831
rect 38856 5828 38884 5859
rect 38930 5856 38936 5908
rect 38988 5896 38994 5908
rect 39025 5899 39083 5905
rect 39025 5896 39037 5899
rect 38988 5868 39037 5896
rect 38988 5856 38994 5868
rect 39025 5865 39037 5868
rect 39071 5865 39083 5899
rect 39025 5859 39083 5865
rect 39393 5899 39451 5905
rect 39393 5865 39405 5899
rect 39439 5896 39451 5899
rect 40494 5896 40500 5908
rect 39439 5868 40500 5896
rect 39439 5865 39451 5868
rect 39393 5859 39451 5865
rect 40494 5856 40500 5868
rect 40552 5896 40558 5908
rect 40773 5899 40831 5905
rect 40773 5896 40785 5899
rect 40552 5868 40785 5896
rect 40552 5856 40558 5868
rect 40773 5865 40785 5868
rect 40819 5865 40831 5899
rect 40773 5859 40831 5865
rect 40862 5856 40868 5908
rect 40920 5896 40926 5908
rect 41509 5899 41567 5905
rect 41509 5896 41521 5899
rect 40920 5868 41521 5896
rect 40920 5856 40926 5868
rect 41509 5865 41521 5868
rect 41555 5865 41567 5899
rect 41509 5859 41567 5865
rect 46198 5856 46204 5908
rect 46256 5856 46262 5908
rect 46382 5856 46388 5908
rect 46440 5856 46446 5908
rect 46750 5856 46756 5908
rect 46808 5896 46814 5908
rect 48866 5896 48872 5908
rect 46808 5868 48872 5896
rect 46808 5856 46814 5868
rect 48866 5856 48872 5868
rect 48924 5856 48930 5908
rect 39209 5831 39267 5837
rect 39209 5828 39221 5831
rect 38856 5800 39221 5828
rect 38289 5791 38347 5797
rect 39209 5797 39221 5800
rect 39255 5797 39267 5831
rect 39209 5791 39267 5797
rect 40037 5831 40095 5837
rect 40037 5797 40049 5831
rect 40083 5828 40095 5831
rect 41230 5828 41236 5840
rect 40083 5800 41236 5828
rect 40083 5797 40095 5800
rect 40037 5791 40095 5797
rect 38059 5732 38240 5760
rect 38059 5729 38071 5732
rect 38013 5723 38071 5729
rect 38105 5695 38163 5701
rect 38105 5661 38117 5695
rect 38151 5692 38163 5695
rect 38194 5692 38200 5704
rect 38151 5664 38200 5692
rect 38151 5661 38163 5664
rect 38105 5655 38163 5661
rect 38194 5652 38200 5664
rect 38252 5652 38258 5704
rect 38304 5692 38332 5791
rect 39224 5760 39252 5791
rect 41230 5788 41236 5800
rect 41288 5788 41294 5840
rect 46106 5788 46112 5840
rect 46164 5788 46170 5840
rect 38764 5732 39160 5760
rect 39224 5732 39620 5760
rect 38657 5695 38715 5701
rect 38657 5692 38669 5695
rect 38304 5664 38669 5692
rect 38657 5661 38669 5664
rect 38703 5661 38715 5695
rect 38657 5655 38715 5661
rect 38764 5624 38792 5732
rect 39132 5701 39160 5732
rect 38841 5695 38899 5701
rect 38841 5661 38853 5695
rect 38887 5692 38899 5695
rect 39117 5695 39175 5701
rect 38887 5664 38976 5692
rect 38887 5661 38899 5664
rect 38841 5655 38899 5661
rect 37936 5596 38792 5624
rect 37829 5587 37887 5593
rect 28966 5528 31432 5556
rect 31478 5516 31484 5568
rect 31536 5516 31542 5568
rect 31570 5516 31576 5568
rect 31628 5556 31634 5568
rect 31941 5559 31999 5565
rect 31941 5556 31953 5559
rect 31628 5528 31953 5556
rect 31628 5516 31634 5528
rect 31941 5525 31953 5528
rect 31987 5525 31999 5559
rect 31941 5519 31999 5525
rect 32122 5516 32128 5568
rect 32180 5516 32186 5568
rect 36170 5516 36176 5568
rect 36228 5516 36234 5568
rect 36446 5516 36452 5568
rect 36504 5516 36510 5568
rect 36814 5516 36820 5568
rect 36872 5556 36878 5568
rect 37182 5556 37188 5568
rect 36872 5528 37188 5556
rect 36872 5516 36878 5528
rect 37182 5516 37188 5528
rect 37240 5556 37246 5568
rect 38948 5556 38976 5664
rect 39117 5661 39129 5695
rect 39163 5692 39175 5695
rect 39301 5695 39359 5701
rect 39163 5664 39252 5692
rect 39163 5661 39175 5664
rect 39117 5655 39175 5661
rect 39224 5568 39252 5664
rect 39301 5661 39313 5695
rect 39347 5661 39359 5695
rect 39301 5655 39359 5661
rect 39316 5568 39344 5655
rect 39390 5652 39396 5704
rect 39448 5652 39454 5704
rect 39592 5701 39620 5732
rect 40402 5720 40408 5772
rect 40460 5720 40466 5772
rect 41322 5720 41328 5772
rect 41380 5760 41386 5772
rect 41693 5763 41751 5769
rect 41693 5760 41705 5763
rect 41380 5732 41705 5760
rect 41380 5720 41386 5732
rect 41693 5729 41705 5732
rect 41739 5729 41751 5763
rect 41693 5723 41751 5729
rect 45741 5763 45799 5769
rect 45741 5729 45753 5763
rect 45787 5760 45799 5763
rect 45830 5760 45836 5772
rect 45787 5732 45836 5760
rect 45787 5729 45799 5732
rect 45741 5723 45799 5729
rect 45830 5720 45836 5732
rect 45888 5720 45894 5772
rect 39577 5695 39635 5701
rect 39577 5661 39589 5695
rect 39623 5661 39635 5695
rect 39577 5655 39635 5661
rect 40218 5652 40224 5704
rect 40276 5652 40282 5704
rect 40420 5692 40448 5720
rect 40497 5695 40555 5701
rect 40497 5692 40509 5695
rect 40420 5664 40509 5692
rect 40497 5661 40509 5664
rect 40543 5692 40555 5695
rect 43533 5695 43591 5701
rect 40543 5664 40724 5692
rect 40543 5661 40555 5664
rect 40497 5655 40555 5661
rect 40696 5636 40724 5664
rect 43533 5661 43545 5695
rect 43579 5692 43591 5695
rect 43898 5692 43904 5704
rect 43579 5664 43904 5692
rect 43579 5661 43591 5664
rect 43533 5655 43591 5661
rect 43898 5652 43904 5664
rect 43956 5652 43962 5704
rect 45925 5695 45983 5701
rect 45925 5661 45937 5695
rect 45971 5692 45983 5695
rect 46124 5692 46152 5788
rect 45971 5664 46152 5692
rect 46216 5692 46244 5856
rect 46290 5720 46296 5772
rect 46348 5760 46354 5772
rect 46845 5763 46903 5769
rect 46845 5760 46857 5763
rect 46348 5732 46857 5760
rect 46348 5720 46354 5732
rect 46845 5729 46857 5732
rect 46891 5760 46903 5763
rect 46934 5760 46940 5772
rect 46891 5732 46940 5760
rect 46891 5729 46903 5732
rect 46845 5723 46903 5729
rect 46934 5720 46940 5732
rect 46992 5720 46998 5772
rect 47394 5720 47400 5772
rect 47452 5720 47458 5772
rect 48424 5732 49004 5760
rect 48424 5704 48452 5732
rect 46569 5695 46627 5701
rect 46569 5692 46581 5695
rect 46216 5664 46581 5692
rect 45971 5661 45983 5664
rect 45925 5655 45983 5661
rect 46569 5661 46581 5664
rect 46615 5661 46627 5695
rect 46569 5655 46627 5661
rect 47026 5652 47032 5704
rect 47084 5692 47090 5704
rect 47121 5695 47179 5701
rect 47121 5692 47133 5695
rect 47084 5664 47133 5692
rect 47084 5652 47090 5664
rect 47121 5661 47133 5664
rect 47167 5661 47179 5695
rect 47121 5655 47179 5661
rect 48406 5652 48412 5704
rect 48464 5652 48470 5704
rect 48976 5701 49004 5732
rect 48961 5695 49019 5701
rect 48961 5661 48973 5695
rect 49007 5661 49019 5695
rect 48961 5655 49019 5661
rect 40589 5627 40647 5633
rect 40589 5593 40601 5627
rect 40635 5593 40647 5627
rect 40589 5587 40647 5593
rect 37240 5528 38976 5556
rect 37240 5516 37246 5528
rect 39206 5516 39212 5568
rect 39264 5516 39270 5568
rect 39298 5516 39304 5568
rect 39356 5516 39362 5568
rect 39666 5516 39672 5568
rect 39724 5556 39730 5568
rect 40405 5559 40463 5565
rect 40405 5556 40417 5559
rect 39724 5528 40417 5556
rect 39724 5516 39730 5528
rect 40405 5525 40417 5528
rect 40451 5556 40463 5559
rect 40604 5556 40632 5587
rect 40678 5584 40684 5636
rect 40736 5624 40742 5636
rect 40789 5627 40847 5633
rect 40789 5624 40801 5627
rect 40736 5596 40801 5624
rect 40736 5584 40742 5596
rect 40789 5593 40801 5596
rect 40835 5593 40847 5627
rect 40789 5587 40847 5593
rect 41138 5584 41144 5636
rect 41196 5584 41202 5636
rect 41325 5627 41383 5633
rect 41325 5593 41337 5627
rect 41371 5593 41383 5627
rect 41325 5587 41383 5593
rect 40451 5528 40632 5556
rect 40451 5525 40463 5528
rect 40405 5519 40463 5525
rect 40954 5516 40960 5568
rect 41012 5516 41018 5568
rect 41340 5556 41368 5587
rect 41966 5584 41972 5636
rect 42024 5584 42030 5636
rect 43625 5627 43683 5633
rect 43625 5624 43637 5627
rect 43194 5596 43637 5624
rect 43625 5593 43637 5596
rect 43671 5593 43683 5627
rect 49053 5627 49111 5633
rect 49053 5624 49065 5627
rect 48622 5596 49065 5624
rect 43625 5587 43683 5593
rect 49053 5593 49065 5596
rect 49099 5593 49111 5627
rect 49053 5587 49111 5593
rect 41414 5556 41420 5568
rect 41340 5528 41420 5556
rect 41414 5516 41420 5528
rect 41472 5556 41478 5568
rect 43441 5559 43499 5565
rect 43441 5556 43453 5559
rect 41472 5528 43453 5556
rect 41472 5516 41478 5528
rect 43441 5525 43453 5528
rect 43487 5525 43499 5559
rect 43441 5519 43499 5525
rect 46109 5559 46167 5565
rect 46109 5525 46121 5559
rect 46155 5556 46167 5559
rect 46842 5556 46848 5568
rect 46155 5528 46848 5556
rect 46155 5525 46167 5528
rect 46109 5519 46167 5525
rect 46842 5516 46848 5528
rect 46900 5516 46906 5568
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 25682 5312 25688 5364
rect 25740 5352 25746 5364
rect 25961 5355 26019 5361
rect 25961 5352 25973 5355
rect 25740 5324 25973 5352
rect 25740 5312 25746 5324
rect 25961 5321 25973 5324
rect 26007 5321 26019 5355
rect 25961 5315 26019 5321
rect 26418 5312 26424 5364
rect 26476 5352 26482 5364
rect 26513 5355 26571 5361
rect 26513 5352 26525 5355
rect 26476 5324 26525 5352
rect 26476 5312 26482 5324
rect 26513 5321 26525 5324
rect 26559 5321 26571 5355
rect 26513 5315 26571 5321
rect 27246 5312 27252 5364
rect 27304 5312 27310 5364
rect 28350 5312 28356 5364
rect 28408 5312 28414 5364
rect 28442 5312 28448 5364
rect 28500 5352 28506 5364
rect 28994 5352 29000 5364
rect 28500 5324 29000 5352
rect 28500 5312 28506 5324
rect 28994 5312 29000 5324
rect 29052 5352 29058 5364
rect 29105 5355 29163 5361
rect 29105 5352 29117 5355
rect 29052 5324 29117 5352
rect 29052 5312 29058 5324
rect 29105 5321 29117 5324
rect 29151 5321 29163 5355
rect 29105 5315 29163 5321
rect 29454 5312 29460 5364
rect 29512 5312 29518 5364
rect 29822 5312 29828 5364
rect 29880 5312 29886 5364
rect 30650 5312 30656 5364
rect 30708 5352 30714 5364
rect 30837 5355 30895 5361
rect 30837 5352 30849 5355
rect 30708 5324 30849 5352
rect 30708 5312 30714 5324
rect 30837 5321 30849 5324
rect 30883 5321 30895 5355
rect 30837 5315 30895 5321
rect 31297 5355 31355 5361
rect 31297 5321 31309 5355
rect 31343 5352 31355 5355
rect 31662 5352 31668 5364
rect 31343 5324 31668 5352
rect 31343 5321 31355 5324
rect 31297 5315 31355 5321
rect 31662 5312 31668 5324
rect 31720 5312 31726 5364
rect 31938 5312 31944 5364
rect 31996 5312 32002 5364
rect 32306 5312 32312 5364
rect 32364 5352 32370 5364
rect 32953 5355 33011 5361
rect 32953 5352 32965 5355
rect 32364 5324 32965 5352
rect 32364 5312 32370 5324
rect 32953 5321 32965 5324
rect 32999 5321 33011 5355
rect 32953 5315 33011 5321
rect 33134 5312 33140 5364
rect 33192 5352 33198 5364
rect 33873 5355 33931 5361
rect 33873 5352 33885 5355
rect 33192 5324 33885 5352
rect 33192 5312 33198 5324
rect 33873 5321 33885 5324
rect 33919 5321 33931 5355
rect 33873 5315 33931 5321
rect 39114 5312 39120 5364
rect 39172 5312 39178 5364
rect 40494 5312 40500 5364
rect 40552 5312 40558 5364
rect 40678 5312 40684 5364
rect 40736 5312 40742 5364
rect 41325 5355 41383 5361
rect 41325 5321 41337 5355
rect 41371 5352 41383 5355
rect 41966 5352 41972 5364
rect 41371 5324 41972 5352
rect 41371 5321 41383 5324
rect 41325 5315 41383 5321
rect 41966 5312 41972 5324
rect 42024 5312 42030 5364
rect 45370 5312 45376 5364
rect 45428 5352 45434 5364
rect 45649 5355 45707 5361
rect 45649 5352 45661 5355
rect 45428 5324 45661 5352
rect 45428 5312 45434 5324
rect 45649 5321 45661 5324
rect 45695 5352 45707 5355
rect 46474 5352 46480 5364
rect 45695 5324 46480 5352
rect 45695 5321 45707 5324
rect 45649 5315 45707 5321
rect 46474 5312 46480 5324
rect 46532 5312 46538 5364
rect 46842 5312 46848 5364
rect 46900 5352 46906 5364
rect 46900 5324 48360 5352
rect 46900 5312 46906 5324
rect 27264 5284 27292 5312
rect 26160 5256 27292 5284
rect 27433 5287 27491 5293
rect 26160 5225 26188 5256
rect 27433 5253 27445 5287
rect 27479 5284 27491 5287
rect 28261 5287 28319 5293
rect 28261 5284 28273 5287
rect 27479 5256 28273 5284
rect 27479 5253 27491 5256
rect 27433 5247 27491 5253
rect 28261 5253 28273 5256
rect 28307 5253 28319 5287
rect 28368 5284 28396 5312
rect 28368 5256 28580 5284
rect 28261 5247 28319 5253
rect 26145 5219 26203 5225
rect 26145 5185 26157 5219
rect 26191 5185 26203 5219
rect 26145 5179 26203 5185
rect 26421 5219 26479 5225
rect 26421 5185 26433 5219
rect 26467 5216 26479 5219
rect 26970 5216 26976 5228
rect 26467 5188 26976 5216
rect 26467 5185 26479 5188
rect 26421 5179 26479 5185
rect 26970 5176 26976 5188
rect 27028 5176 27034 5228
rect 27249 5219 27307 5225
rect 27249 5185 27261 5219
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 27525 5219 27583 5225
rect 27525 5185 27537 5219
rect 27571 5216 27583 5219
rect 27706 5216 27712 5228
rect 27571 5188 27712 5216
rect 27571 5185 27583 5188
rect 27525 5179 27583 5185
rect 27264 5080 27292 5179
rect 27706 5176 27712 5188
rect 27764 5216 27770 5228
rect 28552 5225 28580 5256
rect 28626 5244 28632 5296
rect 28684 5284 28690 5296
rect 28905 5287 28963 5293
rect 28905 5284 28917 5287
rect 28684 5256 28917 5284
rect 28684 5244 28690 5256
rect 28905 5253 28917 5256
rect 28951 5253 28963 5287
rect 28905 5247 28963 5253
rect 28353 5219 28411 5225
rect 28353 5216 28365 5219
rect 27764 5188 28365 5216
rect 27764 5176 27770 5188
rect 28353 5185 28365 5188
rect 28399 5185 28411 5219
rect 28353 5179 28411 5185
rect 28537 5219 28595 5225
rect 28537 5185 28549 5219
rect 28583 5185 28595 5219
rect 28537 5179 28595 5185
rect 28718 5176 28724 5228
rect 28776 5176 28782 5228
rect 28810 5176 28816 5228
rect 28868 5176 28874 5228
rect 29365 5219 29423 5225
rect 29365 5185 29377 5219
rect 29411 5216 29423 5219
rect 29840 5216 29868 5312
rect 30926 5284 30932 5296
rect 30576 5256 30932 5284
rect 30576 5225 30604 5256
rect 30926 5244 30932 5256
rect 30984 5284 30990 5296
rect 31757 5287 31815 5293
rect 31757 5284 31769 5287
rect 30984 5256 31769 5284
rect 30984 5244 30990 5256
rect 31757 5253 31769 5256
rect 31803 5284 31815 5287
rect 31803 5256 33088 5284
rect 31803 5253 31815 5256
rect 31757 5247 31815 5253
rect 29411 5188 29868 5216
rect 30561 5219 30619 5225
rect 29411 5185 29423 5188
rect 29365 5179 29423 5185
rect 30561 5185 30573 5219
rect 30607 5185 30619 5219
rect 30561 5179 30619 5185
rect 30653 5219 30711 5225
rect 30653 5185 30665 5219
rect 30699 5216 30711 5219
rect 31018 5216 31024 5228
rect 30699 5188 31024 5216
rect 30699 5185 30711 5188
rect 30653 5179 30711 5185
rect 31018 5176 31024 5188
rect 31076 5176 31082 5228
rect 31113 5219 31171 5225
rect 31113 5185 31125 5219
rect 31159 5216 31171 5219
rect 31478 5216 31484 5228
rect 31159 5188 31484 5216
rect 31159 5185 31171 5188
rect 31113 5179 31171 5185
rect 31478 5176 31484 5188
rect 31536 5176 31542 5228
rect 31573 5219 31631 5225
rect 31573 5185 31585 5219
rect 31619 5185 31631 5219
rect 31573 5179 31631 5185
rect 27614 5108 27620 5160
rect 27672 5108 27678 5160
rect 28074 5108 28080 5160
rect 28132 5148 28138 5160
rect 28828 5148 28856 5176
rect 28132 5120 28856 5148
rect 28132 5108 28138 5120
rect 30374 5108 30380 5160
rect 30432 5148 30438 5160
rect 30837 5151 30895 5157
rect 30837 5148 30849 5151
rect 30432 5120 30849 5148
rect 30432 5108 30438 5120
rect 29273 5083 29331 5089
rect 29273 5080 29285 5083
rect 27264 5052 29285 5080
rect 29273 5049 29285 5052
rect 29319 5049 29331 5083
rect 29273 5043 29331 5049
rect 30668 5024 30696 5120
rect 30837 5117 30849 5120
rect 30883 5148 30895 5151
rect 31202 5148 31208 5160
rect 30883 5120 31208 5148
rect 30883 5117 30895 5120
rect 30837 5111 30895 5117
rect 31202 5108 31208 5120
rect 31260 5108 31266 5160
rect 31588 5148 31616 5179
rect 32122 5176 32128 5228
rect 32180 5176 32186 5228
rect 33060 5225 33088 5256
rect 35434 5244 35440 5296
rect 35492 5244 35498 5296
rect 36446 5284 36452 5296
rect 36004 5256 36452 5284
rect 36004 5228 36032 5256
rect 36446 5244 36452 5256
rect 36504 5244 36510 5296
rect 32861 5219 32919 5225
rect 32861 5185 32873 5219
rect 32907 5185 32919 5219
rect 32861 5179 32919 5185
rect 33045 5219 33103 5225
rect 33045 5185 33057 5219
rect 33091 5216 33103 5219
rect 33091 5188 33364 5216
rect 33091 5185 33103 5188
rect 33045 5179 33103 5185
rect 32876 5148 32904 5179
rect 33336 5157 33364 5188
rect 35986 5176 35992 5228
rect 36044 5176 36050 5228
rect 36262 5176 36268 5228
rect 36320 5176 36326 5228
rect 39132 5216 39160 5312
rect 39482 5216 39488 5228
rect 39132 5188 39488 5216
rect 39482 5176 39488 5188
rect 39540 5176 39546 5228
rect 39574 5176 39580 5228
rect 39632 5176 39638 5228
rect 40512 5225 40540 5312
rect 41141 5287 41199 5293
rect 41141 5253 41153 5287
rect 41187 5284 41199 5287
rect 43073 5287 43131 5293
rect 43073 5284 43085 5287
rect 41187 5256 43085 5284
rect 41187 5253 41199 5256
rect 41141 5247 41199 5253
rect 43073 5253 43085 5256
rect 43119 5253 43131 5287
rect 43073 5247 43131 5253
rect 44450 5244 44456 5296
rect 44508 5244 44514 5296
rect 45741 5287 45799 5293
rect 45741 5253 45753 5287
rect 45787 5284 45799 5287
rect 46014 5284 46020 5296
rect 45787 5256 46020 5284
rect 45787 5253 45799 5256
rect 45741 5247 45799 5253
rect 46014 5244 46020 5256
rect 46072 5244 46078 5296
rect 47213 5287 47271 5293
rect 47213 5284 47225 5287
rect 46308 5256 47225 5284
rect 40497 5219 40555 5225
rect 40497 5185 40509 5219
rect 40543 5185 40555 5219
rect 40497 5179 40555 5185
rect 40681 5219 40739 5225
rect 40681 5185 40693 5219
rect 40727 5185 40739 5219
rect 40681 5179 40739 5185
rect 33321 5151 33379 5157
rect 31588 5120 33088 5148
rect 33060 5024 33088 5120
rect 33321 5117 33333 5151
rect 33367 5148 33379 5151
rect 33367 5120 33640 5148
rect 33367 5117 33379 5120
rect 33321 5111 33379 5117
rect 33612 5024 33640 5120
rect 33870 5108 33876 5160
rect 33928 5148 33934 5160
rect 34149 5151 34207 5157
rect 34149 5148 34161 5151
rect 33928 5120 34161 5148
rect 33928 5108 33934 5120
rect 34149 5117 34161 5120
rect 34195 5117 34207 5151
rect 34149 5111 34207 5117
rect 34425 5151 34483 5157
rect 34425 5117 34437 5151
rect 34471 5148 34483 5151
rect 36078 5148 36084 5160
rect 34471 5120 36084 5148
rect 34471 5117 34483 5120
rect 34425 5111 34483 5117
rect 36078 5108 36084 5120
rect 36136 5108 36142 5160
rect 36170 5108 36176 5160
rect 36228 5148 36234 5160
rect 36722 5148 36728 5160
rect 36228 5120 36728 5148
rect 36228 5108 36234 5120
rect 36722 5108 36728 5120
rect 36780 5108 36786 5160
rect 39301 5151 39359 5157
rect 39301 5117 39313 5151
rect 39347 5148 39359 5151
rect 39592 5148 39620 5176
rect 39347 5120 39620 5148
rect 40696 5148 40724 5179
rect 40954 5176 40960 5228
rect 41012 5176 41018 5228
rect 41230 5176 41236 5228
rect 41288 5176 41294 5228
rect 41506 5176 41512 5228
rect 41564 5176 41570 5228
rect 46308 5225 46336 5256
rect 47213 5253 47225 5256
rect 47259 5253 47271 5287
rect 47213 5247 47271 5253
rect 46293 5219 46351 5225
rect 46293 5185 46305 5219
rect 46339 5185 46351 5219
rect 46293 5179 46351 5185
rect 46385 5219 46443 5225
rect 46385 5185 46397 5219
rect 46431 5185 46443 5219
rect 46385 5179 46443 5185
rect 41138 5148 41144 5160
rect 40696 5120 41144 5148
rect 39347 5117 39359 5120
rect 39301 5111 39359 5117
rect 41138 5108 41144 5120
rect 41196 5148 41202 5160
rect 42426 5148 42432 5160
rect 41196 5120 42432 5148
rect 41196 5108 41202 5120
rect 42426 5108 42432 5120
rect 42484 5108 42490 5160
rect 43441 5151 43499 5157
rect 43441 5117 43453 5151
rect 43487 5117 43499 5151
rect 43441 5111 43499 5117
rect 36538 5040 36544 5092
rect 36596 5080 36602 5092
rect 36596 5052 40356 5080
rect 36596 5040 36602 5052
rect 40328 5024 40356 5052
rect 27062 4972 27068 5024
rect 27120 4972 27126 5024
rect 29089 5015 29147 5021
rect 29089 4981 29101 5015
rect 29135 5012 29147 5015
rect 29454 5012 29460 5024
rect 29135 4984 29460 5012
rect 29135 4981 29147 4984
rect 29089 4975 29147 4981
rect 29454 4972 29460 4984
rect 29512 4972 29518 5024
rect 30650 4972 30656 5024
rect 30708 4972 30714 5024
rect 32490 4972 32496 5024
rect 32548 5012 32554 5024
rect 32769 5015 32827 5021
rect 32769 5012 32781 5015
rect 32548 4984 32781 5012
rect 32548 4972 32554 4984
rect 32769 4981 32781 4984
rect 32815 4981 32827 5015
rect 32769 4975 32827 4981
rect 33042 4972 33048 5024
rect 33100 4972 33106 5024
rect 33594 4972 33600 5024
rect 33652 4972 33658 5024
rect 36630 4972 36636 5024
rect 36688 4972 36694 5024
rect 37182 4972 37188 5024
rect 37240 5012 37246 5024
rect 39666 5012 39672 5024
rect 37240 4984 39672 5012
rect 37240 4972 37246 4984
rect 39666 4972 39672 4984
rect 39724 4972 39730 5024
rect 40310 4972 40316 5024
rect 40368 4972 40374 5024
rect 40770 4972 40776 5024
rect 40828 4972 40834 5024
rect 43456 5012 43484 5111
rect 43714 5108 43720 5160
rect 43772 5108 43778 5160
rect 45925 5151 45983 5157
rect 45925 5117 45937 5151
rect 45971 5148 45983 5151
rect 46106 5148 46112 5160
rect 45971 5120 46112 5148
rect 45971 5117 45983 5120
rect 45925 5111 45983 5117
rect 45189 5083 45247 5089
rect 45189 5049 45201 5083
rect 45235 5080 45247 5083
rect 45940 5080 45968 5111
rect 46106 5108 46112 5120
rect 46164 5108 46170 5160
rect 45235 5052 45968 5080
rect 45235 5049 45247 5052
rect 45189 5043 45247 5049
rect 45094 5012 45100 5024
rect 43456 4984 45100 5012
rect 45094 4972 45100 4984
rect 45152 4972 45158 5024
rect 45278 4972 45284 5024
rect 45336 4972 45342 5024
rect 45922 4972 45928 5024
rect 45980 5012 45986 5024
rect 46109 5015 46167 5021
rect 46109 5012 46121 5015
rect 45980 4984 46121 5012
rect 45980 4972 45986 4984
rect 46109 4981 46121 4984
rect 46155 4981 46167 5015
rect 46400 5012 46428 5179
rect 46474 5176 46480 5228
rect 46532 5176 46538 5228
rect 46566 5176 46572 5228
rect 46624 5225 46630 5228
rect 46624 5219 46653 5225
rect 46641 5185 46653 5219
rect 46624 5179 46653 5185
rect 46624 5176 46630 5179
rect 46842 5176 46848 5228
rect 46900 5176 46906 5228
rect 46934 5176 46940 5228
rect 46992 5216 46998 5228
rect 47029 5219 47087 5225
rect 47029 5216 47041 5219
rect 46992 5188 47041 5216
rect 46992 5176 46998 5188
rect 47029 5185 47041 5188
rect 47075 5216 47087 5219
rect 47578 5216 47584 5228
rect 47075 5188 47584 5216
rect 47075 5185 47087 5188
rect 47029 5179 47087 5185
rect 47578 5176 47584 5188
rect 47636 5176 47642 5228
rect 48332 5225 48360 5324
rect 48317 5219 48375 5225
rect 48317 5185 48329 5219
rect 48363 5185 48375 5219
rect 48317 5179 48375 5185
rect 48501 5219 48559 5225
rect 48501 5185 48513 5219
rect 48547 5185 48559 5219
rect 48501 5179 48559 5185
rect 46753 5151 46811 5157
rect 46753 5117 46765 5151
rect 46799 5117 46811 5151
rect 47596 5148 47624 5176
rect 48516 5148 48544 5179
rect 47596 5120 48544 5148
rect 46753 5111 46811 5117
rect 46768 5080 46796 5111
rect 48225 5083 48283 5089
rect 48225 5080 48237 5083
rect 46768 5052 48237 5080
rect 48225 5049 48237 5052
rect 48271 5049 48283 5083
rect 48225 5043 48283 5049
rect 48409 5015 48467 5021
rect 48409 5012 48421 5015
rect 46400 4984 48421 5012
rect 46109 4975 46167 4981
rect 48409 4981 48421 4984
rect 48455 4981 48467 5015
rect 48409 4975 48467 4981
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 26040 4811 26098 4817
rect 26040 4777 26052 4811
rect 26086 4808 26098 4811
rect 27062 4808 27068 4820
rect 26086 4780 27068 4808
rect 26086 4777 26098 4780
rect 26040 4771 26098 4777
rect 27062 4768 27068 4780
rect 27120 4768 27126 4820
rect 27525 4811 27583 4817
rect 27525 4777 27537 4811
rect 27571 4808 27583 4811
rect 27614 4808 27620 4820
rect 27571 4780 27620 4808
rect 27571 4777 27583 4780
rect 27525 4771 27583 4777
rect 27614 4768 27620 4780
rect 27672 4808 27678 4820
rect 28169 4811 28227 4817
rect 28169 4808 28181 4811
rect 27672 4780 28181 4808
rect 27672 4768 27678 4780
rect 28169 4777 28181 4780
rect 28215 4808 28227 4811
rect 28534 4808 28540 4820
rect 28215 4780 28540 4808
rect 28215 4777 28227 4780
rect 28169 4771 28227 4777
rect 28534 4768 28540 4780
rect 28592 4768 28598 4820
rect 30466 4768 30472 4820
rect 30524 4808 30530 4820
rect 30561 4811 30619 4817
rect 30561 4808 30573 4811
rect 30524 4780 30573 4808
rect 30524 4768 30530 4780
rect 30561 4777 30573 4780
rect 30607 4777 30619 4811
rect 30561 4771 30619 4777
rect 32112 4811 32170 4817
rect 32112 4777 32124 4811
rect 32158 4808 32170 4811
rect 32490 4808 32496 4820
rect 32158 4780 32496 4808
rect 32158 4777 32170 4780
rect 32112 4771 32170 4777
rect 32490 4768 32496 4780
rect 32548 4768 32554 4820
rect 33594 4768 33600 4820
rect 33652 4768 33658 4820
rect 35069 4811 35127 4817
rect 35069 4777 35081 4811
rect 35115 4808 35127 4811
rect 35434 4808 35440 4820
rect 35115 4780 35440 4808
rect 35115 4777 35127 4780
rect 35069 4771 35127 4777
rect 35434 4768 35440 4780
rect 35492 4768 35498 4820
rect 36078 4768 36084 4820
rect 36136 4768 36142 4820
rect 37458 4768 37464 4820
rect 37516 4808 37522 4820
rect 37516 4780 38240 4808
rect 37516 4768 37522 4780
rect 28353 4743 28411 4749
rect 28353 4709 28365 4743
rect 28399 4740 28411 4743
rect 28902 4740 28908 4752
rect 28399 4712 28908 4740
rect 28399 4709 28411 4712
rect 28353 4703 28411 4709
rect 28902 4700 28908 4712
rect 28960 4700 28966 4752
rect 34054 4700 34060 4752
rect 34112 4700 34118 4752
rect 36262 4700 36268 4752
rect 36320 4740 36326 4752
rect 38105 4743 38163 4749
rect 38105 4740 38117 4743
rect 36320 4712 38117 4740
rect 36320 4700 36326 4712
rect 38105 4709 38117 4712
rect 38151 4709 38163 4743
rect 38105 4703 38163 4709
rect 25590 4632 25596 4684
rect 25648 4672 25654 4684
rect 25777 4675 25835 4681
rect 25777 4672 25789 4675
rect 25648 4644 25789 4672
rect 25648 4632 25654 4644
rect 25777 4641 25789 4644
rect 25823 4672 25835 4675
rect 25823 4644 27476 4672
rect 25823 4641 25835 4644
rect 25777 4635 25835 4641
rect 27448 4616 27476 4644
rect 31846 4632 31852 4684
rect 31904 4672 31910 4684
rect 32766 4672 32772 4684
rect 31904 4644 32772 4672
rect 31904 4632 31910 4644
rect 32766 4632 32772 4644
rect 32824 4672 32830 4684
rect 33870 4672 33876 4684
rect 32824 4644 33876 4672
rect 32824 4632 32830 4644
rect 33870 4632 33876 4644
rect 33928 4632 33934 4684
rect 27430 4564 27436 4616
rect 27488 4564 27494 4616
rect 30650 4564 30656 4616
rect 30708 4604 30714 4616
rect 30745 4607 30803 4613
rect 30745 4604 30757 4607
rect 30708 4576 30757 4604
rect 30708 4564 30714 4576
rect 30745 4573 30757 4576
rect 30791 4573 30803 4607
rect 30745 4567 30803 4573
rect 30926 4564 30932 4616
rect 30984 4564 30990 4616
rect 31021 4607 31079 4613
rect 31021 4573 31033 4607
rect 31067 4573 31079 4607
rect 34072 4604 34100 4700
rect 36280 4672 36308 4700
rect 37921 4675 37979 4681
rect 37921 4672 37933 4675
rect 35820 4644 36308 4672
rect 34606 4604 34612 4616
rect 34072 4576 34612 4604
rect 31021 4567 31079 4573
rect 27062 4496 27068 4548
rect 27120 4496 27126 4548
rect 27982 4496 27988 4548
rect 28040 4496 28046 4548
rect 28201 4539 28259 4545
rect 28201 4505 28213 4539
rect 28247 4536 28259 4539
rect 28247 4508 29040 4536
rect 28247 4505 28259 4508
rect 28201 4499 28259 4505
rect 29012 4480 29040 4508
rect 30558 4496 30564 4548
rect 30616 4536 30622 4548
rect 31036 4536 31064 4567
rect 34606 4564 34612 4576
rect 34664 4604 34670 4616
rect 35820 4613 35848 4644
rect 34977 4607 35035 4613
rect 34977 4604 34989 4607
rect 34664 4576 34989 4604
rect 34664 4564 34670 4576
rect 34977 4573 34989 4576
rect 35023 4573 35035 4607
rect 34977 4567 35035 4573
rect 35805 4607 35863 4613
rect 35805 4573 35817 4607
rect 35851 4573 35863 4607
rect 35805 4567 35863 4573
rect 35986 4564 35992 4616
rect 36044 4564 36050 4616
rect 36280 4613 36308 4644
rect 36372 4644 37933 4672
rect 36372 4613 36400 4644
rect 37921 4641 37933 4644
rect 37967 4641 37979 4675
rect 38212 4672 38240 4780
rect 39482 4768 39488 4820
rect 39540 4768 39546 4820
rect 40770 4768 40776 4820
rect 40828 4768 40834 4820
rect 42426 4768 42432 4820
rect 42484 4808 42490 4820
rect 42889 4811 42947 4817
rect 42889 4808 42901 4811
rect 42484 4780 42901 4808
rect 42484 4768 42490 4780
rect 42889 4777 42901 4780
rect 42935 4777 42947 4811
rect 42889 4771 42947 4777
rect 43714 4768 43720 4820
rect 43772 4808 43778 4820
rect 43993 4811 44051 4817
rect 43993 4808 44005 4811
rect 43772 4780 44005 4808
rect 43772 4768 43778 4780
rect 43993 4777 44005 4780
rect 44039 4777 44051 4811
rect 43993 4771 44051 4777
rect 44450 4768 44456 4820
rect 44508 4768 44514 4820
rect 45278 4768 45284 4820
rect 45336 4768 45342 4820
rect 45820 4811 45878 4817
rect 45820 4777 45832 4811
rect 45866 4808 45878 4811
rect 45922 4808 45928 4820
rect 45866 4780 45928 4808
rect 45866 4777 45878 4780
rect 45820 4771 45878 4777
rect 45922 4768 45928 4780
rect 45980 4768 45986 4820
rect 38378 4700 38384 4752
rect 38436 4740 38442 4752
rect 39390 4740 39396 4752
rect 38436 4712 39396 4740
rect 38436 4700 38442 4712
rect 39390 4700 39396 4712
rect 39448 4700 39454 4752
rect 39574 4672 39580 4684
rect 37921 4635 37979 4641
rect 38028 4644 38240 4672
rect 39316 4644 39580 4672
rect 36265 4607 36323 4613
rect 36265 4573 36277 4607
rect 36311 4573 36323 4607
rect 36265 4567 36323 4573
rect 36357 4607 36415 4613
rect 36357 4573 36369 4607
rect 36403 4573 36415 4607
rect 36357 4567 36415 4573
rect 36538 4564 36544 4616
rect 36596 4613 36602 4616
rect 36596 4607 36625 4613
rect 36613 4573 36625 4607
rect 36596 4567 36625 4573
rect 36596 4564 36602 4567
rect 36722 4564 36728 4616
rect 36780 4564 36786 4616
rect 36814 4564 36820 4616
rect 36872 4564 36878 4616
rect 38028 4613 38056 4644
rect 38013 4607 38071 4613
rect 37476 4576 37872 4604
rect 31386 4536 31392 4548
rect 30616 4508 31392 4536
rect 30616 4496 30622 4508
rect 31386 4496 31392 4508
rect 31444 4496 31450 4548
rect 33134 4496 33140 4548
rect 33192 4496 33198 4548
rect 36449 4539 36507 4545
rect 36449 4505 36461 4539
rect 36495 4505 36507 4539
rect 37476 4536 37504 4576
rect 36449 4499 36507 4505
rect 36740 4508 37504 4536
rect 28994 4428 29000 4480
rect 29052 4428 29058 4480
rect 35986 4428 35992 4480
rect 36044 4428 36050 4480
rect 36464 4468 36492 4499
rect 36740 4468 36768 4508
rect 37550 4496 37556 4548
rect 37608 4496 37614 4548
rect 37737 4539 37795 4545
rect 37737 4505 37749 4539
rect 37783 4505 37795 4539
rect 37844 4536 37872 4576
rect 38013 4573 38025 4607
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 38194 4564 38200 4616
rect 38252 4564 38258 4616
rect 38654 4564 38660 4616
rect 38712 4564 38718 4616
rect 38672 4536 38700 4564
rect 39316 4545 39344 4644
rect 39574 4632 39580 4644
rect 39632 4632 39638 4684
rect 40788 4672 40816 4768
rect 45296 4740 45324 4768
rect 44192 4712 45324 4740
rect 41417 4675 41475 4681
rect 41417 4672 41429 4675
rect 39868 4644 40540 4672
rect 40788 4644 41429 4672
rect 39868 4613 39896 4644
rect 40512 4616 40540 4644
rect 41417 4641 41429 4644
rect 41463 4641 41475 4675
rect 41417 4635 41475 4641
rect 44192 4629 44220 4712
rect 45094 4632 45100 4684
rect 45152 4672 45158 4684
rect 45557 4675 45615 4681
rect 45557 4672 45569 4675
rect 45152 4644 45569 4672
rect 45152 4632 45158 4644
rect 45557 4641 45569 4644
rect 45603 4672 45615 4675
rect 47026 4672 47032 4684
rect 45603 4644 47032 4672
rect 45603 4641 45615 4644
rect 45557 4635 45615 4641
rect 47026 4632 47032 4644
rect 47084 4632 47090 4684
rect 47765 4675 47823 4681
rect 47765 4672 47777 4675
rect 47136 4644 47777 4672
rect 44177 4623 44235 4629
rect 39853 4607 39911 4613
rect 39853 4573 39865 4607
rect 39899 4573 39911 4607
rect 39853 4567 39911 4573
rect 40221 4607 40279 4613
rect 40221 4573 40233 4607
rect 40267 4573 40279 4607
rect 40221 4567 40279 4573
rect 37844 4508 38700 4536
rect 39301 4539 39359 4545
rect 37737 4499 37795 4505
rect 39301 4505 39313 4539
rect 39347 4505 39359 4539
rect 39301 4499 39359 4505
rect 36464 4440 36768 4468
rect 37458 4428 37464 4480
rect 37516 4428 37522 4480
rect 37752 4468 37780 4499
rect 40034 4496 40040 4548
rect 40092 4496 40098 4548
rect 40126 4496 40132 4548
rect 40184 4496 40190 4548
rect 40236 4480 40264 4567
rect 40494 4564 40500 4616
rect 40552 4564 40558 4616
rect 41141 4607 41199 4613
rect 41141 4573 41153 4607
rect 41187 4573 41199 4607
rect 41141 4567 41199 4573
rect 42981 4607 43039 4613
rect 42981 4573 42993 4607
rect 43027 4604 43039 4607
rect 43898 4604 43904 4616
rect 43027 4576 43904 4604
rect 43027 4573 43039 4576
rect 42981 4567 43039 4573
rect 41156 4536 41184 4567
rect 43898 4564 43904 4576
rect 43956 4564 43962 4616
rect 44177 4589 44189 4623
rect 44223 4589 44235 4623
rect 44177 4583 44235 4589
rect 44361 4607 44419 4613
rect 44361 4573 44373 4607
rect 44407 4573 44419 4607
rect 47136 4604 47164 4644
rect 47765 4641 47777 4644
rect 47811 4641 47823 4675
rect 47765 4635 47823 4641
rect 46966 4576 47164 4604
rect 44361 4567 44419 4573
rect 41322 4536 41328 4548
rect 41156 4508 41328 4536
rect 41322 4496 41328 4508
rect 41380 4496 41386 4548
rect 43073 4539 43131 4545
rect 43073 4536 43085 4539
rect 42642 4508 43085 4536
rect 43073 4505 43085 4508
rect 43119 4505 43131 4539
rect 43916 4536 43944 4564
rect 44376 4536 44404 4567
rect 47578 4564 47584 4616
rect 47636 4564 47642 4616
rect 47673 4607 47731 4613
rect 47673 4573 47685 4607
rect 47719 4604 47731 4607
rect 48314 4604 48320 4616
rect 47719 4576 48320 4604
rect 47719 4573 47731 4576
rect 47673 4567 47731 4573
rect 43916 4508 44404 4536
rect 43073 4499 43131 4505
rect 38194 4468 38200 4480
rect 37752 4440 38200 4468
rect 38194 4428 38200 4440
rect 38252 4428 38258 4480
rect 39022 4428 39028 4480
rect 39080 4468 39086 4480
rect 39501 4471 39559 4477
rect 39501 4468 39513 4471
rect 39080 4440 39513 4468
rect 39080 4428 39086 4440
rect 39501 4437 39513 4440
rect 39547 4437 39559 4471
rect 39501 4431 39559 4437
rect 39669 4471 39727 4477
rect 39669 4437 39681 4471
rect 39715 4468 39727 4471
rect 40218 4468 40224 4480
rect 39715 4440 40224 4468
rect 39715 4437 39727 4440
rect 39669 4431 39727 4437
rect 40218 4428 40224 4440
rect 40276 4428 40282 4480
rect 40402 4428 40408 4480
rect 40460 4428 40466 4480
rect 44376 4468 44404 4508
rect 47688 4468 47716 4567
rect 48314 4564 48320 4576
rect 48372 4564 48378 4616
rect 44376 4440 47716 4468
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 27062 4224 27068 4276
rect 27120 4224 27126 4276
rect 28626 4264 28632 4276
rect 28368 4236 28632 4264
rect 28368 4208 28396 4236
rect 28626 4224 28632 4236
rect 28684 4264 28690 4276
rect 31662 4264 31668 4276
rect 28684 4236 31668 4264
rect 28684 4224 28690 4236
rect 28350 4156 28356 4208
rect 28408 4156 28414 4208
rect 28718 4196 28724 4208
rect 28460 4168 28724 4196
rect 26970 4088 26976 4140
rect 27028 4088 27034 4140
rect 26988 4060 27016 4088
rect 28350 4060 28356 4072
rect 26988 4032 28356 4060
rect 28350 4020 28356 4032
rect 28408 4020 28414 4072
rect 28460 4060 28488 4168
rect 28718 4156 28724 4168
rect 28776 4196 28782 4208
rect 30300 4205 30328 4236
rect 31662 4224 31668 4236
rect 31720 4224 31726 4276
rect 35986 4224 35992 4276
rect 36044 4224 36050 4276
rect 36630 4264 36636 4276
rect 36188 4236 36636 4264
rect 30193 4199 30251 4205
rect 30193 4196 30205 4199
rect 28776 4168 30205 4196
rect 28776 4156 28782 4168
rect 30193 4165 30205 4168
rect 30239 4165 30251 4199
rect 30300 4199 30369 4205
rect 30300 4168 30323 4199
rect 30193 4159 30251 4165
rect 30311 4165 30323 4168
rect 30357 4165 30369 4199
rect 31570 4196 31576 4208
rect 30311 4159 30369 4165
rect 30484 4168 31576 4196
rect 28537 4131 28595 4137
rect 28537 4097 28549 4131
rect 28583 4128 28595 4131
rect 29086 4128 29092 4140
rect 28583 4100 29092 4128
rect 28583 4097 28595 4100
rect 28537 4091 28595 4097
rect 29086 4088 29092 4100
rect 29144 4128 29150 4140
rect 29546 4128 29552 4140
rect 29144 4100 29552 4128
rect 29144 4088 29150 4100
rect 29546 4088 29552 4100
rect 29604 4088 29610 4140
rect 30009 4131 30067 4137
rect 30009 4097 30021 4131
rect 30055 4097 30067 4131
rect 30009 4091 30067 4097
rect 28813 4063 28871 4069
rect 28813 4060 28825 4063
rect 28460 4032 28825 4060
rect 28813 4029 28825 4032
rect 28859 4029 28871 4063
rect 30024 4060 30052 4091
rect 30098 4088 30104 4140
rect 30156 4088 30162 4140
rect 30208 4128 30236 4159
rect 30484 4128 30512 4168
rect 31570 4156 31576 4168
rect 31628 4156 31634 4208
rect 34790 4156 34796 4208
rect 34848 4156 34854 4208
rect 30208 4100 30512 4128
rect 32122 4088 32128 4140
rect 32180 4128 32186 4140
rect 32953 4131 33011 4137
rect 32953 4128 32965 4131
rect 32180 4100 32965 4128
rect 32180 4088 32186 4100
rect 32953 4097 32965 4100
rect 32999 4128 33011 4131
rect 33318 4128 33324 4140
rect 32999 4100 33324 4128
rect 32999 4097 33011 4100
rect 32953 4091 33011 4097
rect 33318 4088 33324 4100
rect 33376 4088 33382 4140
rect 33870 4088 33876 4140
rect 33928 4088 33934 4140
rect 36004 4128 36032 4224
rect 36188 4205 36216 4236
rect 36630 4224 36636 4236
rect 36688 4224 36694 4276
rect 36722 4224 36728 4276
rect 36780 4264 36786 4276
rect 38194 4264 38200 4276
rect 36780 4236 38200 4264
rect 36780 4224 36786 4236
rect 38194 4224 38200 4236
rect 38252 4224 38258 4276
rect 38378 4224 38384 4276
rect 38436 4224 38442 4276
rect 38470 4224 38476 4276
rect 38528 4224 38534 4276
rect 38608 4224 38614 4276
rect 38666 4264 38672 4276
rect 39022 4264 39028 4276
rect 38666 4236 39028 4264
rect 38666 4224 38672 4236
rect 39022 4224 39028 4236
rect 39080 4224 39086 4276
rect 39390 4224 39396 4276
rect 39448 4264 39454 4276
rect 39485 4267 39543 4273
rect 39485 4264 39497 4267
rect 39448 4236 39497 4264
rect 39448 4224 39454 4236
rect 39485 4233 39497 4236
rect 39531 4233 39543 4267
rect 39485 4227 39543 4233
rect 40218 4224 40224 4276
rect 40276 4264 40282 4276
rect 40276 4236 40632 4264
rect 40276 4224 40282 4236
rect 36446 4205 36452 4208
rect 36173 4199 36231 4205
rect 36173 4165 36185 4199
rect 36219 4165 36231 4199
rect 36173 4159 36231 4165
rect 36403 4199 36452 4205
rect 36403 4165 36415 4199
rect 36449 4165 36452 4199
rect 36403 4159 36452 4165
rect 36446 4156 36452 4159
rect 36504 4156 36510 4208
rect 37829 4199 37887 4205
rect 37829 4165 37841 4199
rect 37875 4196 37887 4199
rect 38396 4196 38424 4224
rect 40126 4196 40132 4208
rect 37875 4168 38424 4196
rect 38672 4168 39068 4196
rect 37875 4165 37887 4168
rect 37829 4159 37887 4165
rect 36081 4131 36139 4137
rect 36081 4128 36093 4131
rect 36004 4100 36093 4128
rect 36081 4097 36093 4100
rect 36127 4097 36139 4131
rect 36081 4091 36139 4097
rect 36262 4088 36268 4140
rect 36320 4088 36326 4140
rect 36541 4131 36599 4137
rect 36541 4097 36553 4131
rect 36587 4128 36599 4131
rect 37458 4128 37464 4140
rect 36587 4100 37464 4128
rect 36587 4097 36599 4100
rect 36541 4091 36599 4097
rect 37458 4088 37464 4100
rect 37516 4088 37522 4140
rect 37734 4088 37740 4140
rect 37792 4088 37798 4140
rect 37921 4131 37979 4137
rect 37921 4097 37933 4131
rect 37967 4097 37979 4131
rect 38039 4131 38097 4137
rect 38039 4128 38051 4131
rect 37921 4091 37979 4097
rect 38028 4097 38051 4128
rect 38085 4097 38097 4131
rect 38028 4091 38097 4097
rect 30469 4063 30527 4069
rect 30024 4032 30144 4060
rect 28813 4023 28871 4029
rect 28629 3995 28687 4001
rect 28629 3961 28641 3995
rect 28675 3992 28687 3995
rect 28902 3992 28908 4004
rect 28675 3964 28908 3992
rect 28675 3961 28687 3964
rect 28629 3955 28687 3961
rect 28902 3952 28908 3964
rect 28960 3952 28966 4004
rect 28718 3884 28724 3936
rect 28776 3884 28782 3936
rect 29822 3884 29828 3936
rect 29880 3884 29886 3936
rect 30116 3924 30144 4032
rect 30469 4029 30481 4063
rect 30515 4060 30527 4063
rect 30515 4032 30604 4060
rect 30515 4029 30527 4032
rect 30469 4023 30527 4029
rect 30576 3992 30604 4032
rect 30650 4020 30656 4072
rect 30708 4060 30714 4072
rect 30745 4063 30803 4069
rect 30745 4060 30757 4063
rect 30708 4032 30757 4060
rect 30708 4020 30714 4032
rect 30745 4029 30757 4032
rect 30791 4029 30803 4063
rect 30745 4023 30803 4029
rect 33045 4063 33103 4069
rect 33045 4029 33057 4063
rect 33091 4060 33103 4063
rect 33134 4060 33140 4072
rect 33091 4032 33140 4060
rect 33091 4029 33103 4032
rect 33045 4023 33103 4029
rect 33134 4020 33140 4032
rect 33192 4020 33198 4072
rect 34149 4063 34207 4069
rect 34149 4029 34161 4063
rect 34195 4060 34207 4063
rect 35897 4063 35955 4069
rect 35897 4060 35909 4063
rect 34195 4032 35909 4060
rect 34195 4029 34207 4032
rect 34149 4023 34207 4029
rect 35897 4029 35909 4032
rect 35943 4029 35955 4063
rect 36280 4060 36308 4088
rect 37182 4060 37188 4072
rect 36280 4032 37188 4060
rect 35897 4023 35955 4029
rect 37182 4020 37188 4032
rect 37240 4060 37246 4072
rect 37936 4060 37964 4091
rect 37240 4032 37964 4060
rect 37240 4020 37246 4032
rect 31389 3995 31447 4001
rect 31389 3992 31401 3995
rect 30576 3964 31401 3992
rect 31389 3961 31401 3964
rect 31435 3961 31447 3995
rect 31389 3955 31447 3961
rect 35621 3995 35679 4001
rect 35621 3961 35633 3995
rect 35667 3992 35679 3995
rect 36814 3992 36820 4004
rect 35667 3964 36820 3992
rect 35667 3961 35679 3964
rect 35621 3955 35679 3961
rect 36814 3952 36820 3964
rect 36872 3952 36878 4004
rect 38028 3992 38056 4091
rect 38378 4088 38384 4140
rect 38436 4088 38442 4140
rect 38565 4138 38623 4143
rect 38672 4138 38700 4168
rect 38565 4137 38700 4138
rect 38565 4103 38577 4137
rect 38611 4110 38700 4137
rect 38611 4103 38623 4110
rect 38565 4097 38623 4103
rect 38197 4063 38255 4069
rect 38197 4029 38209 4063
rect 38243 4029 38255 4063
rect 38197 4023 38255 4029
rect 38657 4063 38715 4069
rect 38657 4029 38669 4063
rect 38703 4029 38715 4063
rect 39040 4060 39068 4168
rect 39408 4168 40132 4196
rect 39408 4140 39436 4168
rect 40126 4156 40132 4168
rect 40184 4156 40190 4208
rect 40310 4156 40316 4208
rect 40368 4196 40374 4208
rect 40368 4168 40448 4196
rect 40368 4156 40374 4168
rect 39390 4088 39396 4140
rect 39448 4088 39454 4140
rect 40420 4128 40448 4168
rect 40494 4156 40500 4208
rect 40552 4156 40558 4208
rect 40604 4205 40632 4236
rect 40589 4199 40647 4205
rect 40589 4165 40601 4199
rect 40635 4165 40647 4199
rect 40773 4199 40831 4205
rect 40773 4196 40785 4199
rect 40589 4159 40647 4165
rect 40696 4168 40785 4196
rect 40696 4128 40724 4168
rect 40773 4165 40785 4168
rect 40819 4165 40831 4199
rect 40773 4159 40831 4165
rect 40420 4100 40724 4128
rect 41049 4131 41107 4137
rect 41049 4097 41061 4131
rect 41095 4097 41107 4131
rect 41049 4091 41107 4097
rect 39206 4060 39212 4072
rect 39040 4032 39212 4060
rect 38657 4023 38715 4029
rect 37200 3964 38056 3992
rect 30466 3924 30472 3936
rect 30116 3896 30472 3924
rect 30466 3884 30472 3896
rect 30524 3884 30530 3936
rect 36538 3884 36544 3936
rect 36596 3924 36602 3936
rect 37200 3924 37228 3964
rect 38102 3952 38108 4004
rect 38160 3992 38166 4004
rect 38212 3992 38240 4023
rect 38160 3964 38240 3992
rect 38160 3952 38166 3964
rect 38286 3952 38292 4004
rect 38344 3992 38350 4004
rect 38672 3992 38700 4023
rect 39206 4020 39212 4032
rect 39264 4060 39270 4072
rect 39942 4060 39948 4072
rect 39264 4032 39948 4060
rect 39264 4020 39270 4032
rect 39942 4020 39948 4032
rect 40000 4020 40006 4072
rect 40586 4020 40592 4072
rect 40644 4060 40650 4072
rect 41064 4060 41092 4091
rect 40644 4032 41092 4060
rect 40644 4020 40650 4032
rect 38344 3964 38700 3992
rect 39301 3995 39359 4001
rect 38344 3952 38350 3964
rect 39301 3961 39313 3995
rect 39347 3961 39359 3995
rect 39301 3955 39359 3961
rect 36596 3896 37228 3924
rect 36596 3884 36602 3896
rect 37550 3884 37556 3936
rect 37608 3884 37614 3936
rect 38562 3884 38568 3936
rect 38620 3924 38626 3936
rect 39316 3924 39344 3955
rect 38620 3896 39344 3924
rect 38620 3884 38626 3896
rect 40034 3884 40040 3936
rect 40092 3924 40098 3936
rect 40957 3927 41015 3933
rect 40957 3924 40969 3927
rect 40092 3896 40969 3924
rect 40092 3884 40098 3896
rect 40957 3893 40969 3896
rect 41003 3893 41015 3927
rect 40957 3887 41015 3893
rect 41141 3927 41199 3933
rect 41141 3893 41153 3927
rect 41187 3924 41199 3927
rect 41414 3924 41420 3936
rect 41187 3896 41420 3924
rect 41187 3893 41199 3896
rect 41141 3887 41199 3893
rect 41414 3884 41420 3896
rect 41472 3884 41478 3936
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 28718 3680 28724 3732
rect 28776 3680 28782 3732
rect 28902 3680 28908 3732
rect 28960 3680 28966 3732
rect 30098 3680 30104 3732
rect 30156 3680 30162 3732
rect 30742 3680 30748 3732
rect 30800 3680 30806 3732
rect 31278 3723 31336 3729
rect 31278 3720 31290 3723
rect 30852 3692 31290 3720
rect 28736 3652 28764 3680
rect 28368 3624 28764 3652
rect 28368 3525 28396 3624
rect 28626 3544 28632 3596
rect 28684 3584 28690 3596
rect 28721 3587 28779 3593
rect 28721 3584 28733 3587
rect 28684 3556 28733 3584
rect 28684 3544 28690 3556
rect 28721 3553 28733 3556
rect 28767 3553 28779 3587
rect 28721 3547 28779 3553
rect 28261 3519 28319 3525
rect 28261 3485 28273 3519
rect 28307 3485 28319 3519
rect 28261 3479 28319 3485
rect 28353 3519 28411 3525
rect 28353 3485 28365 3519
rect 28399 3485 28411 3519
rect 28353 3479 28411 3485
rect 28813 3519 28871 3525
rect 28813 3485 28825 3519
rect 28859 3485 28871 3519
rect 28920 3516 28948 3680
rect 30285 3655 30343 3661
rect 30285 3621 30297 3655
rect 30331 3652 30343 3655
rect 30852 3652 30880 3692
rect 31278 3689 31290 3692
rect 31324 3689 31336 3723
rect 31278 3683 31336 3689
rect 34790 3680 34796 3732
rect 34848 3680 34854 3732
rect 37734 3680 37740 3732
rect 37792 3720 37798 3732
rect 38289 3723 38347 3729
rect 38289 3720 38301 3723
rect 37792 3692 38301 3720
rect 37792 3680 37798 3692
rect 38289 3689 38301 3692
rect 38335 3689 38347 3723
rect 38289 3683 38347 3689
rect 39390 3680 39396 3732
rect 39448 3680 39454 3732
rect 39942 3680 39948 3732
rect 40000 3720 40006 3732
rect 41785 3723 41843 3729
rect 41785 3720 41797 3723
rect 40000 3692 41797 3720
rect 40000 3680 40006 3692
rect 41785 3689 41797 3692
rect 41831 3689 41843 3723
rect 41785 3683 41843 3689
rect 30331 3624 30880 3652
rect 30929 3655 30987 3661
rect 30331 3621 30343 3624
rect 30285 3615 30343 3621
rect 30929 3621 30941 3655
rect 30975 3621 30987 3655
rect 30929 3615 30987 3621
rect 38197 3655 38255 3661
rect 38197 3621 38209 3655
rect 38243 3652 38255 3655
rect 38378 3652 38384 3664
rect 38243 3624 38384 3652
rect 38243 3621 38255 3624
rect 38197 3615 38255 3621
rect 30944 3584 30972 3615
rect 38378 3612 38384 3624
rect 38436 3652 38442 3664
rect 39408 3652 39436 3680
rect 38436 3624 39436 3652
rect 38436 3612 38442 3624
rect 41414 3612 41420 3664
rect 41472 3612 41478 3664
rect 30024 3556 30972 3584
rect 31021 3587 31079 3593
rect 30024 3525 30052 3556
rect 31021 3553 31033 3587
rect 31067 3584 31079 3587
rect 31846 3584 31852 3596
rect 31067 3556 31852 3584
rect 31067 3553 31079 3556
rect 31021 3547 31079 3553
rect 31846 3544 31852 3556
rect 31904 3544 31910 3596
rect 36541 3587 36599 3593
rect 36541 3553 36553 3587
rect 36587 3584 36599 3587
rect 37366 3584 37372 3596
rect 36587 3556 37372 3584
rect 36587 3553 36599 3556
rect 36541 3547 36599 3553
rect 37366 3544 37372 3556
rect 37424 3544 37430 3596
rect 37645 3587 37703 3593
rect 37645 3553 37657 3587
rect 37691 3584 37703 3587
rect 38286 3584 38292 3596
rect 37691 3556 38292 3584
rect 37691 3553 37703 3556
rect 37645 3547 37703 3553
rect 38286 3544 38292 3556
rect 38344 3584 38350 3596
rect 38749 3587 38807 3593
rect 38749 3584 38761 3587
rect 38344 3556 38761 3584
rect 38344 3544 38350 3556
rect 38749 3553 38761 3556
rect 38795 3553 38807 3587
rect 38749 3547 38807 3553
rect 40034 3544 40040 3596
rect 40092 3584 40098 3596
rect 41322 3584 41328 3596
rect 40092 3556 41328 3584
rect 40092 3544 40098 3556
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 28997 3519 29055 3525
rect 28997 3516 29009 3519
rect 28920 3488 29009 3516
rect 28813 3479 28871 3485
rect 28997 3485 29009 3488
rect 29043 3516 29055 3519
rect 30009 3519 30067 3525
rect 30009 3516 30021 3519
rect 29043 3488 30021 3516
rect 29043 3485 29055 3488
rect 28997 3479 29055 3485
rect 30009 3485 30021 3488
rect 30055 3485 30067 3519
rect 30009 3479 30067 3485
rect 27798 3340 27804 3392
rect 27856 3380 27862 3392
rect 28077 3383 28135 3389
rect 28077 3380 28089 3383
rect 27856 3352 28089 3380
rect 27856 3340 27862 3352
rect 28077 3349 28089 3352
rect 28123 3349 28135 3383
rect 28276 3380 28304 3479
rect 28629 3451 28687 3457
rect 28629 3417 28641 3451
rect 28675 3448 28687 3451
rect 28828 3448 28856 3479
rect 30466 3476 30472 3528
rect 30524 3476 30530 3528
rect 34606 3476 34612 3528
rect 34664 3516 34670 3528
rect 34701 3519 34759 3525
rect 34701 3516 34713 3519
rect 34664 3488 34713 3516
rect 34664 3476 34670 3488
rect 34701 3485 34713 3488
rect 34747 3485 34759 3519
rect 34701 3479 34759 3485
rect 36262 3476 36268 3528
rect 36320 3476 36326 3528
rect 36814 3476 36820 3528
rect 36872 3476 36878 3528
rect 37384 3516 37412 3544
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 37384 3488 38025 3516
rect 38013 3485 38025 3488
rect 38059 3516 38071 3519
rect 38473 3519 38531 3525
rect 38473 3516 38485 3519
rect 38059 3488 38485 3516
rect 38059 3485 38071 3488
rect 38013 3479 38071 3485
rect 38473 3485 38485 3488
rect 38519 3485 38531 3519
rect 38473 3479 38531 3485
rect 38565 3519 38623 3525
rect 38565 3485 38577 3519
rect 38611 3485 38623 3519
rect 38565 3479 38623 3485
rect 38657 3519 38715 3525
rect 38657 3485 38669 3519
rect 38703 3485 38715 3519
rect 38657 3479 38715 3485
rect 39117 3519 39175 3525
rect 39117 3485 39129 3519
rect 39163 3516 39175 3519
rect 39298 3516 39304 3528
rect 39163 3488 39304 3516
rect 39163 3485 39175 3488
rect 39117 3479 39175 3485
rect 29086 3448 29092 3460
rect 28675 3420 29092 3448
rect 28675 3417 28687 3420
rect 28629 3411 28687 3417
rect 29086 3408 29092 3420
rect 29144 3408 29150 3460
rect 30561 3451 30619 3457
rect 30561 3417 30573 3451
rect 30607 3448 30619 3451
rect 30650 3448 30656 3460
rect 30607 3420 30656 3448
rect 30607 3417 30619 3420
rect 30561 3411 30619 3417
rect 30650 3408 30656 3420
rect 30708 3408 30714 3460
rect 30777 3451 30835 3457
rect 30777 3417 30789 3451
rect 30823 3448 30835 3451
rect 31386 3448 31392 3460
rect 30823 3420 31392 3448
rect 30823 3417 30835 3420
rect 30777 3411 30835 3417
rect 31386 3408 31392 3420
rect 31444 3408 31450 3460
rect 32306 3408 32312 3460
rect 32364 3408 32370 3460
rect 33042 3408 33048 3460
rect 33100 3408 33106 3460
rect 36357 3451 36415 3457
rect 36357 3417 36369 3451
rect 36403 3448 36415 3451
rect 36538 3448 36544 3460
rect 36403 3420 36544 3448
rect 36403 3417 36415 3420
rect 36357 3411 36415 3417
rect 36538 3408 36544 3420
rect 36596 3408 36602 3460
rect 36832 3448 36860 3476
rect 37829 3451 37887 3457
rect 37829 3448 37841 3451
rect 36832 3420 37841 3448
rect 37829 3417 37841 3420
rect 37875 3417 37887 3451
rect 37829 3411 37887 3417
rect 37921 3451 37979 3457
rect 37921 3417 37933 3451
rect 37967 3448 37979 3451
rect 38194 3448 38200 3460
rect 37967 3420 38200 3448
rect 37967 3417 37979 3420
rect 37921 3411 37979 3417
rect 28994 3380 29000 3392
rect 28276 3352 29000 3380
rect 28077 3343 28135 3349
rect 28994 3340 29000 3352
rect 29052 3380 29058 3392
rect 29181 3383 29239 3389
rect 29181 3380 29193 3383
rect 29052 3352 29193 3380
rect 29052 3340 29058 3352
rect 29181 3349 29193 3352
rect 29227 3349 29239 3383
rect 29181 3343 29239 3349
rect 35894 3340 35900 3392
rect 35952 3340 35958 3392
rect 37844 3380 37872 3411
rect 38194 3408 38200 3420
rect 38252 3448 38258 3460
rect 38580 3448 38608 3479
rect 38252 3420 38608 3448
rect 38252 3408 38258 3420
rect 38672 3380 38700 3479
rect 39298 3476 39304 3488
rect 39356 3476 39362 3528
rect 41432 3502 41460 3612
rect 68462 3476 68468 3528
rect 68520 3476 68526 3528
rect 40313 3451 40371 3457
rect 40313 3417 40325 3451
rect 40359 3448 40371 3451
rect 40402 3448 40408 3460
rect 40359 3420 40408 3448
rect 40359 3417 40371 3420
rect 40313 3411 40371 3417
rect 40402 3408 40408 3420
rect 40460 3408 40466 3460
rect 37844 3352 38700 3380
rect 39390 3340 39396 3392
rect 39448 3380 39454 3392
rect 39669 3383 39727 3389
rect 39669 3380 39681 3383
rect 39448 3352 39681 3380
rect 39448 3340 39454 3352
rect 39669 3349 39681 3352
rect 39715 3349 39727 3383
rect 39669 3343 39727 3349
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 27430 3136 27436 3188
rect 27488 3176 27494 3188
rect 27488 3148 29408 3176
rect 27488 3136 27494 3148
rect 27448 3049 27476 3136
rect 27709 3111 27767 3117
rect 27709 3077 27721 3111
rect 27755 3108 27767 3111
rect 27798 3108 27804 3120
rect 27755 3080 27804 3108
rect 27755 3077 27767 3080
rect 27709 3071 27767 3077
rect 27798 3068 27804 3080
rect 27856 3068 27862 3120
rect 28442 3068 28448 3120
rect 28500 3068 28506 3120
rect 29380 3049 29408 3148
rect 29822 3136 29828 3188
rect 29880 3136 29886 3188
rect 30466 3136 30472 3188
rect 30524 3176 30530 3188
rect 31205 3179 31263 3185
rect 31205 3176 31217 3179
rect 30524 3148 31217 3176
rect 30524 3136 30530 3148
rect 31205 3145 31217 3148
rect 31251 3145 31263 3179
rect 31205 3139 31263 3145
rect 31570 3136 31576 3188
rect 31628 3136 31634 3188
rect 31662 3136 31668 3188
rect 31720 3136 31726 3188
rect 32217 3179 32275 3185
rect 32217 3145 32229 3179
rect 32263 3176 32275 3179
rect 32306 3176 32312 3188
rect 32263 3148 32312 3176
rect 32263 3145 32275 3148
rect 32217 3139 32275 3145
rect 32306 3136 32312 3148
rect 32364 3136 32370 3188
rect 32858 3136 32864 3188
rect 32916 3136 32922 3188
rect 34698 3136 34704 3188
rect 34756 3176 34762 3188
rect 37366 3176 37372 3188
rect 34756 3148 37044 3176
rect 34756 3136 34762 3148
rect 29641 3111 29699 3117
rect 29641 3077 29653 3111
rect 29687 3108 29699 3111
rect 29840 3108 29868 3136
rect 29687 3080 29868 3108
rect 29687 3077 29699 3080
rect 29641 3071 29699 3077
rect 30374 3068 30380 3120
rect 30432 3068 30438 3120
rect 27433 3043 27491 3049
rect 27433 3009 27445 3043
rect 27479 3009 27491 3043
rect 27433 3003 27491 3009
rect 29365 3043 29423 3049
rect 29365 3009 29377 3043
rect 29411 3009 29423 3043
rect 29365 3003 29423 3009
rect 32122 3000 32128 3052
rect 32180 3000 32186 3052
rect 32677 3043 32735 3049
rect 32677 3009 32689 3043
rect 32723 3040 32735 3043
rect 32876 3040 32904 3136
rect 36354 3068 36360 3120
rect 36412 3068 36418 3120
rect 32723 3012 32904 3040
rect 37016 3040 37044 3148
rect 37108 3148 37372 3176
rect 37108 3117 37136 3148
rect 37366 3136 37372 3148
rect 37424 3136 37430 3188
rect 38286 3136 38292 3188
rect 38344 3176 38350 3188
rect 39025 3179 39083 3185
rect 39025 3176 39037 3179
rect 38344 3148 39037 3176
rect 38344 3136 38350 3148
rect 39025 3145 39037 3148
rect 39071 3145 39083 3179
rect 39025 3139 39083 3145
rect 39224 3148 41414 3176
rect 37093 3111 37151 3117
rect 37093 3077 37105 3111
rect 37139 3077 37151 3111
rect 37642 3108 37648 3120
rect 37093 3071 37151 3077
rect 37292 3080 37648 3108
rect 37292 3040 37320 3080
rect 37642 3068 37648 3080
rect 37700 3068 37706 3120
rect 37016 3012 37320 3040
rect 32723 3009 32735 3012
rect 32677 3003 32735 3009
rect 38654 3000 38660 3052
rect 38712 3000 38718 3052
rect 39022 3000 39028 3052
rect 39080 3040 39086 3052
rect 39117 3043 39175 3049
rect 39117 3040 39129 3043
rect 39080 3012 39129 3040
rect 39080 3000 39086 3012
rect 39117 3009 39129 3012
rect 39163 3009 39175 3043
rect 39117 3003 39175 3009
rect 30650 2932 30656 2984
rect 30708 2972 30714 2984
rect 31113 2975 31171 2981
rect 31113 2972 31125 2975
rect 30708 2944 31125 2972
rect 30708 2932 30714 2944
rect 31113 2941 31125 2944
rect 31159 2941 31171 2975
rect 31113 2935 31171 2941
rect 31386 2932 31392 2984
rect 31444 2972 31450 2984
rect 31757 2975 31815 2981
rect 31757 2972 31769 2975
rect 31444 2944 31769 2972
rect 31444 2932 31450 2944
rect 31757 2941 31769 2944
rect 31803 2972 31815 2975
rect 33042 2972 33048 2984
rect 31803 2944 33048 2972
rect 31803 2941 31815 2944
rect 31757 2935 31815 2941
rect 33042 2932 33048 2944
rect 33100 2932 33106 2984
rect 33870 2932 33876 2984
rect 33928 2972 33934 2984
rect 35069 2975 35127 2981
rect 35069 2972 35081 2975
rect 33928 2944 35081 2972
rect 33928 2932 33934 2944
rect 35069 2941 35081 2944
rect 35115 2941 35127 2975
rect 35069 2935 35127 2941
rect 29086 2864 29092 2916
rect 29144 2904 29150 2916
rect 29181 2907 29239 2913
rect 29181 2904 29193 2907
rect 29144 2876 29193 2904
rect 29144 2864 29150 2876
rect 29181 2873 29193 2876
rect 29227 2873 29239 2907
rect 29181 2867 29239 2873
rect 31846 2864 31852 2916
rect 31904 2904 31910 2916
rect 31904 2876 32904 2904
rect 31904 2864 31910 2876
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 31110 2836 31116 2848
rect 22612 2808 31116 2836
rect 22612 2796 22618 2808
rect 31110 2796 31116 2808
rect 31168 2796 31174 2848
rect 32876 2845 32904 2876
rect 32861 2839 32919 2845
rect 32861 2805 32873 2839
rect 32907 2805 32919 2839
rect 35084 2836 35112 2935
rect 35342 2932 35348 2984
rect 35400 2932 35406 2984
rect 37277 2975 37335 2981
rect 37277 2941 37289 2975
rect 37323 2941 37335 2975
rect 37277 2935 37335 2941
rect 37292 2836 37320 2935
rect 37550 2932 37556 2984
rect 37608 2932 37614 2984
rect 37642 2932 37648 2984
rect 37700 2972 37706 2984
rect 39224 2972 39252 3148
rect 40034 3108 40040 3120
rect 39684 3080 40040 3108
rect 39298 3000 39304 3052
rect 39356 3000 39362 3052
rect 39684 3049 39712 3080
rect 40034 3068 40040 3080
rect 40092 3068 40098 3120
rect 40678 3068 40684 3120
rect 40736 3068 40742 3120
rect 39669 3043 39727 3049
rect 39669 3009 39681 3043
rect 39715 3009 39727 3043
rect 41386 3040 41414 3148
rect 47765 3043 47823 3049
rect 47765 3040 47777 3043
rect 41386 3012 47777 3040
rect 39669 3003 39727 3009
rect 47765 3009 47777 3012
rect 47811 3009 47823 3043
rect 47765 3003 47823 3009
rect 37700 2944 39252 2972
rect 37700 2932 37706 2944
rect 35084 2808 37320 2836
rect 32861 2799 32919 2805
rect 39114 2796 39120 2848
rect 39172 2796 39178 2848
rect 39316 2836 39344 3000
rect 39942 2932 39948 2984
rect 40000 2932 40006 2984
rect 41417 2839 41475 2845
rect 41417 2836 41429 2839
rect 39316 2808 41429 2836
rect 41417 2805 41429 2808
rect 41463 2805 41475 2839
rect 41417 2799 41475 2805
rect 47581 2839 47639 2845
rect 47581 2805 47593 2839
rect 47627 2836 47639 2839
rect 48314 2836 48320 2848
rect 47627 2808 48320 2836
rect 47627 2805 47639 2808
rect 47581 2799 47639 2805
rect 48314 2796 48320 2808
rect 48372 2796 48378 2848
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 28442 2592 28448 2644
rect 28500 2632 28506 2644
rect 28537 2635 28595 2641
rect 28537 2632 28549 2635
rect 28500 2604 28549 2632
rect 28500 2592 28506 2604
rect 28537 2601 28549 2604
rect 28583 2601 28595 2635
rect 28537 2595 28595 2601
rect 30374 2592 30380 2644
rect 30432 2592 30438 2644
rect 32122 2592 32128 2644
rect 32180 2592 32186 2644
rect 34606 2592 34612 2644
rect 34664 2592 34670 2644
rect 35342 2592 35348 2644
rect 35400 2632 35406 2644
rect 35621 2635 35679 2641
rect 35621 2632 35633 2635
rect 35400 2604 35633 2632
rect 35400 2592 35406 2604
rect 35621 2601 35633 2604
rect 35667 2601 35679 2635
rect 35621 2595 35679 2601
rect 36265 2635 36323 2641
rect 36265 2601 36277 2635
rect 36311 2632 36323 2635
rect 36354 2632 36360 2644
rect 36311 2604 36360 2632
rect 36311 2601 36323 2604
rect 36265 2595 36323 2601
rect 36354 2592 36360 2604
rect 36412 2592 36418 2644
rect 38289 2635 38347 2641
rect 38289 2601 38301 2635
rect 38335 2632 38347 2635
rect 38654 2632 38660 2644
rect 38335 2604 38660 2632
rect 38335 2601 38347 2604
rect 38289 2595 38347 2601
rect 38654 2592 38660 2604
rect 38712 2592 38718 2644
rect 39669 2635 39727 2641
rect 39669 2601 39681 2635
rect 39715 2632 39727 2635
rect 39942 2632 39948 2644
rect 39715 2604 39948 2632
rect 39715 2601 39727 2604
rect 39669 2595 39727 2601
rect 39942 2592 39948 2604
rect 40000 2592 40006 2644
rect 40678 2592 40684 2644
rect 40736 2592 40742 2644
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 1857 2567 1915 2573
rect 1857 2564 1869 2567
rect 72 2536 1869 2564
rect 72 2524 78 2536
rect 1857 2533 1869 2536
rect 1903 2533 1915 2567
rect 1857 2527 1915 2533
rect 32140 2496 32168 2592
rect 30300 2468 32168 2496
rect 34624 2496 34652 2592
rect 35802 2524 35808 2576
rect 35860 2564 35866 2576
rect 36081 2567 36139 2573
rect 36081 2564 36093 2567
rect 35860 2536 36093 2564
rect 35860 2524 35866 2536
rect 36081 2533 36093 2536
rect 36127 2533 36139 2567
rect 40586 2564 40592 2576
rect 36081 2527 36139 2533
rect 38212 2536 40592 2564
rect 34624 2468 36216 2496
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 992 2400 1593 2428
rect 992 2388 998 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2225 2431 2283 2437
rect 2225 2428 2237 2431
rect 2004 2400 2237 2428
rect 2004 2388 2010 2400
rect 2225 2397 2237 2400
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7156 2400 7389 2428
rect 7156 2388 7162 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9732 2400 9965 2428
rect 9732 2388 9738 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17460 2400 17693 2428
rect 17460 2388 17466 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 25409 2431 25467 2437
rect 25409 2428 25421 2431
rect 25188 2400 25421 2428
rect 25188 2388 25194 2400
rect 25409 2397 25421 2400
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 30300 2437 30328 2468
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 28408 2400 28457 2428
rect 28408 2388 28414 2400
rect 28445 2397 28457 2400
rect 28491 2428 28503 2431
rect 30285 2431 30343 2437
rect 30285 2428 30297 2431
rect 28491 2400 30297 2428
rect 28491 2397 28503 2400
rect 28445 2391 28503 2397
rect 30285 2397 30297 2400
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 30466 2388 30472 2440
rect 30524 2428 30530 2440
rect 30745 2431 30803 2437
rect 30745 2428 30757 2431
rect 30524 2400 30757 2428
rect 30524 2388 30530 2400
rect 30745 2397 30757 2400
rect 30791 2397 30803 2431
rect 30745 2391 30803 2397
rect 33134 2388 33140 2440
rect 33192 2388 33198 2440
rect 35805 2431 35863 2437
rect 35805 2397 35817 2431
rect 35851 2428 35863 2431
rect 35894 2428 35900 2440
rect 35851 2400 35900 2428
rect 35851 2397 35863 2400
rect 35805 2391 35863 2397
rect 35894 2388 35900 2400
rect 35952 2388 35958 2440
rect 36188 2437 36216 2468
rect 38212 2437 38240 2536
rect 40586 2524 40592 2536
rect 40644 2524 40650 2576
rect 39666 2496 39672 2508
rect 39132 2468 39672 2496
rect 36173 2431 36231 2437
rect 36173 2397 36185 2431
rect 36219 2428 36231 2431
rect 38197 2431 38255 2437
rect 38197 2428 38209 2431
rect 36219 2400 38209 2428
rect 36219 2397 36231 2400
rect 36173 2391 36231 2397
rect 38197 2397 38209 2400
rect 38243 2397 38255 2431
rect 38197 2391 38255 2397
rect 38286 2388 38292 2440
rect 38344 2428 38350 2440
rect 39132 2437 39160 2468
rect 39666 2456 39672 2468
rect 39724 2456 39730 2508
rect 38657 2431 38715 2437
rect 38657 2428 38669 2431
rect 38344 2400 38669 2428
rect 38344 2388 38350 2400
rect 38657 2397 38669 2400
rect 38703 2397 38715 2431
rect 38657 2391 38715 2397
rect 39117 2431 39175 2437
rect 39117 2397 39129 2431
rect 39163 2397 39175 2431
rect 39117 2391 39175 2397
rect 39390 2388 39396 2440
rect 39448 2388 39454 2440
rect 39485 2431 39543 2437
rect 39485 2397 39497 2431
rect 39531 2428 39543 2431
rect 40126 2428 40132 2440
rect 39531 2400 40132 2428
rect 39531 2397 39543 2400
rect 39485 2391 39543 2397
rect 40126 2388 40132 2400
rect 40184 2388 40190 2440
rect 40604 2437 40632 2524
rect 68005 2499 68063 2505
rect 68005 2465 68017 2499
rect 68051 2496 68063 2499
rect 68051 2468 68692 2496
rect 68051 2465 68063 2468
rect 68005 2459 68063 2465
rect 68664 2440 68692 2468
rect 40589 2431 40647 2437
rect 40589 2397 40601 2431
rect 40635 2397 40647 2431
rect 40589 2391 40647 2397
rect 43162 2388 43168 2440
rect 43220 2428 43226 2440
rect 43441 2431 43499 2437
rect 43441 2428 43453 2431
rect 43220 2400 43453 2428
rect 43220 2388 43226 2400
rect 43441 2397 43453 2400
rect 43487 2397 43499 2431
rect 43441 2391 43499 2397
rect 45738 2388 45744 2440
rect 45796 2428 45802 2440
rect 46017 2431 46075 2437
rect 46017 2428 46029 2431
rect 45796 2400 46029 2428
rect 45796 2388 45802 2400
rect 46017 2397 46029 2400
rect 46063 2397 46075 2431
rect 46017 2391 46075 2397
rect 48314 2388 48320 2440
rect 48372 2428 48378 2440
rect 48501 2431 48559 2437
rect 48501 2428 48513 2431
rect 48372 2400 48513 2428
rect 48372 2388 48378 2400
rect 48501 2397 48513 2400
rect 48547 2397 48559 2431
rect 48501 2391 48559 2397
rect 50890 2388 50896 2440
rect 50948 2428 50954 2440
rect 51169 2431 51227 2437
rect 51169 2428 51181 2431
rect 50948 2400 51181 2428
rect 50948 2388 50954 2400
rect 51169 2397 51181 2400
rect 51215 2397 51227 2431
rect 51169 2391 51227 2397
rect 53466 2388 53472 2440
rect 53524 2428 53530 2440
rect 53745 2431 53803 2437
rect 53745 2428 53757 2431
rect 53524 2400 53757 2428
rect 53524 2388 53530 2400
rect 53745 2397 53757 2400
rect 53791 2397 53803 2431
rect 53745 2391 53803 2397
rect 56042 2388 56048 2440
rect 56100 2428 56106 2440
rect 56321 2431 56379 2437
rect 56321 2428 56333 2431
rect 56100 2400 56333 2428
rect 56100 2388 56106 2400
rect 56321 2397 56333 2400
rect 56367 2397 56379 2431
rect 56321 2391 56379 2397
rect 58618 2388 58624 2440
rect 58676 2428 58682 2440
rect 58897 2431 58955 2437
rect 58897 2428 58909 2431
rect 58676 2400 58909 2428
rect 58676 2388 58682 2400
rect 58897 2397 58909 2400
rect 58943 2397 58955 2431
rect 58897 2391 58955 2397
rect 66346 2388 66352 2440
rect 66404 2428 66410 2440
rect 66625 2431 66683 2437
rect 66625 2428 66637 2431
rect 66404 2400 66637 2428
rect 66404 2388 66410 2400
rect 66625 2397 66637 2400
rect 66671 2397 66683 2431
rect 66625 2391 66683 2397
rect 68462 2388 68468 2440
rect 68520 2388 68526 2440
rect 68646 2388 68652 2440
rect 68704 2388 68710 2440
rect 12437 2363 12495 2369
rect 12437 2329 12449 2363
rect 12483 2360 12495 2363
rect 31754 2360 31760 2372
rect 12483 2332 31760 2360
rect 12483 2329 12495 2332
rect 12437 2323 12495 2329
rect 31754 2320 31760 2332
rect 31812 2320 31818 2372
rect 39206 2320 39212 2372
rect 39264 2360 39270 2372
rect 39301 2363 39359 2369
rect 39301 2360 39313 2363
rect 39264 2332 39313 2360
rect 39264 2320 39270 2332
rect 39301 2329 39313 2332
rect 39347 2329 39359 2363
rect 39301 2323 39359 2329
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 12529 2295 12587 2301
rect 12529 2292 12541 2295
rect 12400 2264 12541 2292
rect 12400 2252 12406 2264
rect 12529 2261 12541 2264
rect 12575 2261 12587 2295
rect 12529 2255 12587 2261
rect 48314 2252 48320 2304
rect 48372 2292 48378 2304
rect 48593 2295 48651 2301
rect 48593 2292 48605 2295
rect 48372 2264 48605 2292
rect 48372 2252 48378 2264
rect 48593 2261 48605 2264
rect 48639 2261 48651 2295
rect 48593 2255 48651 2261
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
<< via1 >>
rect 19574 67430 19626 67482
rect 19638 67430 19690 67482
rect 19702 67430 19754 67482
rect 19766 67430 19818 67482
rect 19830 67430 19882 67482
rect 50294 67430 50346 67482
rect 50358 67430 50410 67482
rect 50422 67430 50474 67482
rect 50486 67430 50538 67482
rect 50550 67430 50602 67482
rect 56140 67371 56192 67380
rect 56140 67337 56149 67371
rect 56149 67337 56183 67371
rect 56183 67337 56192 67371
rect 56140 67328 56192 67337
rect 940 67192 992 67244
rect 2228 67235 2280 67244
rect 2228 67201 2237 67235
rect 2237 67201 2271 67235
rect 2271 67201 2280 67235
rect 2228 67192 2280 67201
rect 4804 67235 4856 67244
rect 4804 67201 4813 67235
rect 4813 67201 4847 67235
rect 4847 67201 4856 67235
rect 4804 67192 4856 67201
rect 7380 67235 7432 67244
rect 7380 67201 7389 67235
rect 7389 67201 7423 67235
rect 7423 67201 7432 67235
rect 7380 67192 7432 67201
rect 9956 67235 10008 67244
rect 9956 67201 9965 67235
rect 9965 67201 9999 67235
rect 9999 67201 10008 67235
rect 9956 67192 10008 67201
rect 12440 67192 12492 67244
rect 15108 67235 15160 67244
rect 15108 67201 15117 67235
rect 15117 67201 15151 67235
rect 15151 67201 15160 67235
rect 15108 67192 15160 67201
rect 17684 67235 17736 67244
rect 17684 67201 17693 67235
rect 17693 67201 17727 67235
rect 17727 67201 17736 67235
rect 17684 67192 17736 67201
rect 20260 67235 20312 67244
rect 20260 67201 20269 67235
rect 20269 67201 20303 67235
rect 20303 67201 20312 67235
rect 20260 67192 20312 67201
rect 22836 67235 22888 67244
rect 22836 67201 22845 67235
rect 22845 67201 22879 67235
rect 22879 67201 22888 67235
rect 22836 67192 22888 67201
rect 25412 67235 25464 67244
rect 25412 67201 25421 67235
rect 25421 67201 25455 67235
rect 25455 67201 25464 67235
rect 25412 67192 25464 67201
rect 27988 67235 28040 67244
rect 27988 67201 27997 67235
rect 27997 67201 28031 67235
rect 28031 67201 28040 67235
rect 27988 67192 28040 67201
rect 30380 67192 30432 67244
rect 33140 67235 33192 67244
rect 33140 67201 33149 67235
rect 33149 67201 33183 67235
rect 33183 67201 33192 67235
rect 33140 67192 33192 67201
rect 38292 67235 38344 67244
rect 38292 67201 38301 67235
rect 38301 67201 38335 67235
rect 38335 67201 38344 67235
rect 38292 67192 38344 67201
rect 40868 67235 40920 67244
rect 40868 67201 40877 67235
rect 40877 67201 40911 67235
rect 40911 67201 40920 67235
rect 40868 67192 40920 67201
rect 46020 67235 46072 67244
rect 46020 67201 46029 67235
rect 46029 67201 46063 67235
rect 46063 67201 46072 67235
rect 46020 67192 46072 67201
rect 53748 67235 53800 67244
rect 53748 67201 53757 67235
rect 53757 67201 53791 67235
rect 53791 67201 53800 67235
rect 53748 67192 53800 67201
rect 58900 67235 58952 67244
rect 58900 67201 58909 67235
rect 58909 67201 58943 67235
rect 58943 67201 58952 67235
rect 58900 67192 58952 67201
rect 61476 67235 61528 67244
rect 61476 67201 61485 67235
rect 61485 67201 61519 67235
rect 61519 67201 61528 67235
rect 61476 67192 61528 67201
rect 64052 67235 64104 67244
rect 64052 67201 64061 67235
rect 64061 67201 64095 67235
rect 64095 67201 64104 67235
rect 64052 67192 64104 67201
rect 68928 67192 68980 67244
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 19574 66342 19626 66394
rect 19638 66342 19690 66394
rect 19702 66342 19754 66394
rect 19766 66342 19818 66394
rect 19830 66342 19882 66394
rect 50294 66342 50346 66394
rect 50358 66342 50410 66394
rect 50422 66342 50474 66394
rect 50486 66342 50538 66394
rect 50550 66342 50602 66394
rect 68468 66011 68520 66020
rect 68468 65977 68477 66011
rect 68477 65977 68511 66011
rect 68511 65977 68520 66011
rect 68468 65968 68520 65977
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 19574 65254 19626 65306
rect 19638 65254 19690 65306
rect 19702 65254 19754 65306
rect 19766 65254 19818 65306
rect 19830 65254 19882 65306
rect 50294 65254 50346 65306
rect 50358 65254 50410 65306
rect 50422 65254 50474 65306
rect 50486 65254 50538 65306
rect 50550 65254 50602 65306
rect 1584 64923 1636 64932
rect 1584 64889 1593 64923
rect 1593 64889 1627 64923
rect 1627 64889 1636 64923
rect 1584 64880 1636 64889
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 34934 64710 34986 64762
rect 34998 64710 35050 64762
rect 35062 64710 35114 64762
rect 35126 64710 35178 64762
rect 35190 64710 35242 64762
rect 65654 64710 65706 64762
rect 65718 64710 65770 64762
rect 65782 64710 65834 64762
rect 65846 64710 65898 64762
rect 65910 64710 65962 64762
rect 19574 64166 19626 64218
rect 19638 64166 19690 64218
rect 19702 64166 19754 64218
rect 19766 64166 19818 64218
rect 19830 64166 19882 64218
rect 50294 64166 50346 64218
rect 50358 64166 50410 64218
rect 50422 64166 50474 64218
rect 50486 64166 50538 64218
rect 50550 64166 50602 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 34934 63622 34986 63674
rect 34998 63622 35050 63674
rect 35062 63622 35114 63674
rect 35126 63622 35178 63674
rect 35190 63622 35242 63674
rect 65654 63622 65706 63674
rect 65718 63622 65770 63674
rect 65782 63622 65834 63674
rect 65846 63622 65898 63674
rect 65910 63622 65962 63674
rect 68468 63359 68520 63368
rect 68468 63325 68477 63359
rect 68477 63325 68511 63359
rect 68511 63325 68520 63359
rect 68468 63316 68520 63325
rect 19574 63078 19626 63130
rect 19638 63078 19690 63130
rect 19702 63078 19754 63130
rect 19766 63078 19818 63130
rect 19830 63078 19882 63130
rect 50294 63078 50346 63130
rect 50358 63078 50410 63130
rect 50422 63078 50474 63130
rect 50486 63078 50538 63130
rect 50550 63078 50602 63130
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 34934 62534 34986 62586
rect 34998 62534 35050 62586
rect 35062 62534 35114 62586
rect 35126 62534 35178 62586
rect 35190 62534 35242 62586
rect 65654 62534 65706 62586
rect 65718 62534 65770 62586
rect 65782 62534 65834 62586
rect 65846 62534 65898 62586
rect 65910 62534 65962 62586
rect 19574 61990 19626 62042
rect 19638 61990 19690 62042
rect 19702 61990 19754 62042
rect 19766 61990 19818 62042
rect 19830 61990 19882 62042
rect 50294 61990 50346 62042
rect 50358 61990 50410 62042
rect 50422 61990 50474 62042
rect 50486 61990 50538 62042
rect 50550 61990 50602 62042
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 65654 61446 65706 61498
rect 65718 61446 65770 61498
rect 65782 61446 65834 61498
rect 65846 61446 65898 61498
rect 65910 61446 65962 61498
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 68192 60707 68244 60716
rect 68192 60673 68201 60707
rect 68201 60673 68235 60707
rect 68235 60673 68244 60707
rect 68192 60664 68244 60673
rect 68376 60571 68428 60580
rect 68376 60537 68385 60571
rect 68385 60537 68419 60571
rect 68419 60537 68428 60571
rect 68376 60528 68428 60537
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 65654 60358 65706 60410
rect 65718 60358 65770 60410
rect 65782 60358 65834 60410
rect 65846 60358 65898 60410
rect 65910 60358 65962 60410
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 1584 59415 1636 59424
rect 1584 59381 1593 59415
rect 1593 59381 1627 59415
rect 1627 59381 1636 59415
rect 1584 59372 1636 59381
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 65654 59270 65706 59322
rect 65718 59270 65770 59322
rect 65782 59270 65834 59322
rect 65846 59270 65898 59322
rect 65910 59270 65962 59322
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 65654 58182 65706 58234
rect 65718 58182 65770 58234
rect 65782 58182 65834 58234
rect 65846 58182 65898 58234
rect 65910 58182 65962 58234
rect 68468 57919 68520 57928
rect 68468 57885 68477 57919
rect 68477 57885 68511 57919
rect 68511 57885 68520 57919
rect 68468 57876 68520 57885
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 1584 56831 1636 56840
rect 1584 56797 1593 56831
rect 1593 56797 1627 56831
rect 1627 56797 1636 56831
rect 1584 56788 1636 56797
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 68468 55131 68520 55140
rect 68468 55097 68477 55131
rect 68477 55097 68511 55131
rect 68511 55097 68520 55131
rect 68468 55088 68520 55097
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 68468 52479 68520 52488
rect 68468 52445 68477 52479
rect 68477 52445 68511 52479
rect 68511 52445 68520 52479
rect 68468 52436 68520 52445
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 940 51348 992 51400
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 68468 49759 68520 49768
rect 68468 49725 68477 49759
rect 68477 49725 68511 49759
rect 68511 49725 68520 49759
rect 68468 49716 68520 49725
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 940 48492 992 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 68468 47039 68520 47048
rect 68468 47005 68477 47039
rect 68477 47005 68511 47039
rect 68511 47005 68520 47039
rect 68468 46996 68520 47005
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 940 45908 992 45960
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 68468 44251 68520 44260
rect 68468 44217 68477 44251
rect 68477 44217 68511 44251
rect 68511 44217 68520 44251
rect 68468 44208 68520 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 940 43052 992 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 68468 41599 68520 41608
rect 68468 41565 68477 41599
rect 68477 41565 68511 41599
rect 68511 41565 68520 41599
rect 68468 41556 68520 41565
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 940 37612 992 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 68468 36159 68520 36168
rect 68468 36125 68477 36159
rect 68477 36125 68511 36159
rect 68511 36125 68520 36159
rect 68468 36116 68520 36125
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 940 35028 992 35080
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 68744 33464 68796 33516
rect 68376 33303 68428 33312
rect 68376 33269 68385 33303
rect 68385 33269 68419 33303
rect 68419 33269 68428 33303
rect 68376 33260 68428 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 940 32172 992 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 68468 30719 68520 30728
rect 68468 30685 68477 30719
rect 68477 30685 68511 30719
rect 68511 30685 68520 30719
rect 68468 30676 68520 30685
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 940 29588 992 29640
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 68468 27931 68520 27940
rect 68468 27897 68477 27931
rect 68477 27897 68511 27931
rect 68511 27897 68520 27931
rect 68468 27888 68520 27897
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 940 26732 992 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 28908 25279 28960 25288
rect 28908 25245 28917 25279
rect 28917 25245 28951 25279
rect 28951 25245 28960 25279
rect 28908 25236 28960 25245
rect 31208 25279 31260 25288
rect 31208 25245 31217 25279
rect 31217 25245 31251 25279
rect 31251 25245 31260 25279
rect 31208 25236 31260 25245
rect 68468 25279 68520 25288
rect 68468 25245 68477 25279
rect 68477 25245 68511 25279
rect 68511 25245 68520 25279
rect 68468 25236 68520 25245
rect 29552 25168 29604 25220
rect 28816 25143 28868 25152
rect 28816 25109 28825 25143
rect 28825 25109 28859 25143
rect 28859 25109 28868 25143
rect 28816 25100 28868 25109
rect 30932 25100 30984 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 31208 24896 31260 24948
rect 31668 24896 31720 24948
rect 28816 24828 28868 24880
rect 30288 24803 30340 24812
rect 30288 24769 30322 24803
rect 30322 24769 30340 24803
rect 30288 24760 30340 24769
rect 31852 24760 31904 24812
rect 32496 24760 32548 24812
rect 34060 24828 34112 24880
rect 34244 24803 34296 24812
rect 34244 24769 34278 24803
rect 34278 24769 34296 24803
rect 34244 24760 34296 24769
rect 36084 24760 36136 24812
rect 30012 24735 30064 24744
rect 30012 24701 30021 24735
rect 30021 24701 30055 24735
rect 30055 24701 30064 24735
rect 30012 24692 30064 24701
rect 29460 24556 29512 24608
rect 35348 24599 35400 24608
rect 35348 24565 35357 24599
rect 35357 24565 35391 24599
rect 35391 24565 35400 24599
rect 35348 24556 35400 24565
rect 36820 24599 36872 24608
rect 36820 24565 36829 24599
rect 36829 24565 36863 24599
rect 36863 24565 36872 24599
rect 36820 24556 36872 24565
rect 37004 24556 37056 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 28908 24352 28960 24404
rect 29552 24352 29604 24404
rect 31208 24352 31260 24404
rect 31576 24352 31628 24404
rect 940 24148 992 24200
rect 30564 24284 30616 24336
rect 35348 24352 35400 24404
rect 37004 24352 37056 24404
rect 31024 24216 31076 24268
rect 31852 24259 31904 24268
rect 31852 24225 31861 24259
rect 31861 24225 31895 24259
rect 31895 24225 31904 24259
rect 31852 24216 31904 24225
rect 35532 24284 35584 24336
rect 35900 24216 35952 24268
rect 29460 24148 29512 24200
rect 29552 24191 29604 24200
rect 29552 24157 29561 24191
rect 29561 24157 29595 24191
rect 29595 24157 29604 24191
rect 29552 24148 29604 24157
rect 30564 24191 30616 24200
rect 30564 24157 30573 24191
rect 30573 24157 30607 24191
rect 30607 24157 30616 24191
rect 30564 24148 30616 24157
rect 31392 24148 31444 24200
rect 29920 24012 29972 24064
rect 31300 24080 31352 24132
rect 31484 24012 31536 24064
rect 31760 24055 31812 24064
rect 31760 24021 31769 24055
rect 31769 24021 31803 24055
rect 31803 24021 31812 24055
rect 31760 24012 31812 24021
rect 36268 24216 36320 24268
rect 36544 24148 36596 24200
rect 36728 24191 36780 24200
rect 36728 24157 36737 24191
rect 36737 24157 36771 24191
rect 36771 24157 36780 24191
rect 36728 24148 36780 24157
rect 36452 24080 36504 24132
rect 37740 24080 37792 24132
rect 35900 24012 35952 24064
rect 36360 24055 36412 24064
rect 36360 24021 36369 24055
rect 36369 24021 36403 24055
rect 36403 24021 36412 24055
rect 36360 24012 36412 24021
rect 37556 24012 37608 24064
rect 37832 24012 37884 24064
rect 38292 24012 38344 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 30288 23808 30340 23860
rect 27160 23715 27212 23724
rect 27160 23681 27169 23715
rect 27169 23681 27203 23715
rect 27203 23681 27212 23715
rect 27160 23672 27212 23681
rect 28448 23715 28500 23724
rect 28448 23681 28457 23715
rect 28457 23681 28491 23715
rect 28491 23681 28500 23715
rect 28448 23672 28500 23681
rect 29092 23740 29144 23792
rect 29552 23783 29604 23792
rect 29552 23749 29561 23783
rect 29561 23749 29595 23783
rect 29595 23749 29604 23783
rect 29552 23740 29604 23749
rect 28908 23604 28960 23656
rect 29184 23715 29236 23724
rect 29184 23681 29193 23715
rect 29193 23681 29227 23715
rect 29227 23681 29236 23715
rect 29184 23672 29236 23681
rect 29460 23672 29512 23724
rect 32220 23808 32272 23860
rect 31300 23783 31352 23792
rect 31300 23749 31309 23783
rect 31309 23749 31343 23783
rect 31343 23749 31352 23783
rect 31300 23740 31352 23749
rect 31576 23740 31628 23792
rect 35348 23808 35400 23860
rect 30932 23604 30984 23656
rect 31760 23715 31812 23724
rect 31760 23681 31769 23715
rect 31769 23681 31803 23715
rect 31803 23681 31812 23715
rect 31760 23672 31812 23681
rect 32220 23672 32272 23724
rect 34704 23740 34756 23792
rect 32404 23672 32456 23724
rect 31944 23604 31996 23656
rect 32956 23604 33008 23656
rect 26976 23511 27028 23520
rect 26976 23477 26985 23511
rect 26985 23477 27019 23511
rect 27019 23477 27028 23511
rect 26976 23468 27028 23477
rect 28080 23511 28132 23520
rect 28080 23477 28089 23511
rect 28089 23477 28123 23511
rect 28123 23477 28132 23511
rect 28080 23468 28132 23477
rect 30196 23468 30248 23520
rect 34244 23536 34296 23588
rect 35532 23672 35584 23724
rect 35624 23647 35676 23656
rect 35624 23613 35633 23647
rect 35633 23613 35667 23647
rect 35667 23613 35676 23647
rect 35624 23604 35676 23613
rect 35348 23536 35400 23588
rect 35808 23647 35860 23656
rect 35808 23613 35817 23647
rect 35817 23613 35851 23647
rect 35851 23613 35860 23647
rect 35808 23604 35860 23613
rect 35900 23647 35952 23656
rect 35900 23613 35909 23647
rect 35909 23613 35943 23647
rect 35943 23613 35952 23647
rect 35900 23604 35952 23613
rect 36084 23808 36136 23860
rect 36360 23808 36412 23860
rect 36452 23808 36504 23860
rect 36544 23740 36596 23792
rect 36820 23715 36872 23724
rect 36820 23681 36829 23715
rect 36829 23681 36863 23715
rect 36863 23681 36872 23715
rect 36820 23672 36872 23681
rect 37188 23672 37240 23724
rect 38568 23740 38620 23792
rect 39304 23672 39356 23724
rect 45560 23672 45612 23724
rect 46848 23672 46900 23724
rect 36820 23536 36872 23588
rect 37832 23604 37884 23656
rect 47032 23604 47084 23656
rect 35440 23468 35492 23520
rect 37372 23468 37424 23520
rect 37464 23468 37516 23520
rect 38292 23536 38344 23588
rect 38384 23511 38436 23520
rect 38384 23477 38393 23511
rect 38393 23477 38427 23511
rect 38427 23477 38436 23511
rect 38384 23468 38436 23477
rect 38568 23468 38620 23520
rect 46112 23468 46164 23520
rect 46940 23468 46992 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 28448 23264 28500 23316
rect 30196 23264 30248 23316
rect 31024 23307 31076 23316
rect 31024 23273 31033 23307
rect 31033 23273 31067 23307
rect 31067 23273 31076 23307
rect 31024 23264 31076 23273
rect 32680 23264 32732 23316
rect 33048 23264 33100 23316
rect 34520 23264 34572 23316
rect 34704 23264 34756 23316
rect 35348 23264 35400 23316
rect 36544 23264 36596 23316
rect 36728 23264 36780 23316
rect 37096 23264 37148 23316
rect 37740 23307 37792 23316
rect 37740 23273 37749 23307
rect 37749 23273 37783 23307
rect 37783 23273 37792 23307
rect 37740 23264 37792 23273
rect 26608 23103 26660 23112
rect 26608 23069 26617 23103
rect 26617 23069 26651 23103
rect 26651 23069 26660 23103
rect 26608 23060 26660 23069
rect 29184 23128 29236 23180
rect 29460 23128 29512 23180
rect 28908 23103 28960 23112
rect 28908 23069 28917 23103
rect 28917 23069 28951 23103
rect 28951 23069 28960 23103
rect 28908 23060 28960 23069
rect 29092 23103 29144 23112
rect 29092 23069 29101 23103
rect 29101 23069 29135 23103
rect 29135 23069 29144 23103
rect 29092 23060 29144 23069
rect 29920 23128 29972 23180
rect 31116 23128 31168 23180
rect 26976 22992 27028 23044
rect 28540 22967 28592 22976
rect 28540 22933 28549 22967
rect 28549 22933 28583 22967
rect 28583 22933 28592 22967
rect 28540 22924 28592 22933
rect 29276 22924 29328 22976
rect 31852 23171 31904 23180
rect 31852 23137 31861 23171
rect 31861 23137 31895 23171
rect 31895 23137 31904 23171
rect 31852 23128 31904 23137
rect 31668 23103 31720 23112
rect 31668 23069 31677 23103
rect 31677 23069 31711 23103
rect 31711 23069 31720 23103
rect 31300 23035 31352 23044
rect 31300 23001 31309 23035
rect 31309 23001 31343 23035
rect 31343 23001 31352 23035
rect 31300 22992 31352 23001
rect 31668 23060 31720 23069
rect 32312 23103 32364 23112
rect 32312 23069 32321 23103
rect 32321 23069 32355 23103
rect 32355 23069 32364 23103
rect 32312 23060 32364 23069
rect 32496 23060 32548 23112
rect 35624 23196 35676 23248
rect 37556 23196 37608 23248
rect 34520 23103 34572 23112
rect 34520 23069 34529 23103
rect 34529 23069 34563 23103
rect 34563 23069 34572 23103
rect 34520 23060 34572 23069
rect 35440 23103 35492 23112
rect 35440 23069 35449 23103
rect 35449 23069 35483 23103
rect 35483 23069 35492 23103
rect 36452 23128 36504 23180
rect 35440 23060 35492 23069
rect 36544 23060 36596 23112
rect 30196 22924 30248 22976
rect 30380 22967 30432 22976
rect 30380 22933 30389 22967
rect 30389 22933 30423 22967
rect 30423 22933 30432 22967
rect 30380 22924 30432 22933
rect 31024 22924 31076 22976
rect 31484 22924 31536 22976
rect 32036 23035 32088 23044
rect 32036 23001 32045 23035
rect 32045 23001 32079 23035
rect 32079 23001 32088 23035
rect 32036 22992 32088 23001
rect 32128 22992 32180 23044
rect 32680 23035 32732 23044
rect 32680 23001 32714 23035
rect 32714 23001 32732 23035
rect 32680 22992 32732 23001
rect 32496 22924 32548 22976
rect 34796 22924 34848 22976
rect 35348 22924 35400 22976
rect 37188 23128 37240 23180
rect 37372 23128 37424 23180
rect 38384 23196 38436 23248
rect 37464 23060 37516 23112
rect 38568 23171 38620 23180
rect 38568 23137 38577 23171
rect 38577 23137 38611 23171
rect 38611 23137 38620 23171
rect 38568 23128 38620 23137
rect 39304 23307 39356 23316
rect 39304 23273 39313 23307
rect 39313 23273 39347 23307
rect 39347 23273 39356 23307
rect 39304 23264 39356 23273
rect 46848 23196 46900 23248
rect 48044 23128 48096 23180
rect 38016 23035 38068 23044
rect 38016 23001 38025 23035
rect 38025 23001 38059 23035
rect 38059 23001 38068 23035
rect 38016 22992 38068 23001
rect 36820 22924 36872 22976
rect 37740 22924 37792 22976
rect 38292 22992 38344 23044
rect 45468 23060 45520 23112
rect 46940 23060 46992 23112
rect 49516 23103 49568 23112
rect 49516 23069 49525 23103
rect 49525 23069 49559 23103
rect 49559 23069 49568 23103
rect 49516 23060 49568 23069
rect 46112 22992 46164 23044
rect 47952 23035 48004 23044
rect 47952 23001 47961 23035
rect 47961 23001 47995 23035
rect 47995 23001 48004 23035
rect 47952 22992 48004 23001
rect 44456 22924 44508 22976
rect 45100 22967 45152 22976
rect 45100 22933 45109 22967
rect 45109 22933 45143 22967
rect 45143 22933 45152 22967
rect 45100 22924 45152 22933
rect 47584 22924 47636 22976
rect 49424 22967 49476 22976
rect 49424 22933 49433 22967
rect 49433 22933 49467 22967
rect 49467 22933 49476 22967
rect 49424 22924 49476 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 27160 22720 27212 22772
rect 28080 22720 28132 22772
rect 30288 22720 30340 22772
rect 31208 22720 31260 22772
rect 32128 22720 32180 22772
rect 31484 22695 31536 22704
rect 30840 22584 30892 22636
rect 31484 22661 31493 22695
rect 31493 22661 31527 22695
rect 31527 22661 31536 22695
rect 31484 22652 31536 22661
rect 32496 22652 32548 22704
rect 34796 22720 34848 22772
rect 35440 22763 35492 22772
rect 35440 22729 35449 22763
rect 35449 22729 35483 22763
rect 35483 22729 35492 22763
rect 35440 22720 35492 22729
rect 35624 22720 35676 22772
rect 36268 22720 36320 22772
rect 38292 22720 38344 22772
rect 45008 22720 45060 22772
rect 47124 22720 47176 22772
rect 34060 22627 34112 22636
rect 34060 22593 34069 22627
rect 34069 22593 34103 22627
rect 34103 22593 34112 22627
rect 34060 22584 34112 22593
rect 37372 22652 37424 22704
rect 38016 22652 38068 22704
rect 44088 22652 44140 22704
rect 45100 22652 45152 22704
rect 47308 22652 47360 22704
rect 26700 22516 26752 22568
rect 31300 22516 31352 22568
rect 31576 22516 31628 22568
rect 31668 22516 31720 22568
rect 32036 22516 32088 22568
rect 33324 22559 33376 22568
rect 33324 22525 33333 22559
rect 33333 22525 33367 22559
rect 33367 22525 33376 22559
rect 33324 22516 33376 22525
rect 37464 22516 37516 22568
rect 43628 22516 43680 22568
rect 44364 22559 44416 22568
rect 44364 22525 44373 22559
rect 44373 22525 44407 22559
rect 44407 22525 44416 22559
rect 44364 22516 44416 22525
rect 30472 22380 30524 22432
rect 30748 22423 30800 22432
rect 30748 22389 30757 22423
rect 30757 22389 30791 22423
rect 30791 22389 30800 22423
rect 30748 22380 30800 22389
rect 39028 22448 39080 22500
rect 46572 22584 46624 22636
rect 46848 22627 46900 22636
rect 46848 22593 46857 22627
rect 46857 22593 46891 22627
rect 46891 22593 46900 22627
rect 46848 22584 46900 22593
rect 48872 22627 48924 22636
rect 48872 22593 48881 22627
rect 48881 22593 48915 22627
rect 48915 22593 48924 22627
rect 48872 22584 48924 22593
rect 49424 22584 49476 22636
rect 47584 22559 47636 22568
rect 47584 22525 47593 22559
rect 47593 22525 47627 22559
rect 47627 22525 47636 22559
rect 47584 22516 47636 22525
rect 68468 22491 68520 22500
rect 68468 22457 68477 22491
rect 68477 22457 68511 22491
rect 68511 22457 68520 22491
rect 68468 22448 68520 22457
rect 32404 22380 32456 22432
rect 38752 22423 38804 22432
rect 38752 22389 38761 22423
rect 38761 22389 38795 22423
rect 38795 22389 38804 22423
rect 38752 22380 38804 22389
rect 46664 22380 46716 22432
rect 47400 22380 47452 22432
rect 48320 22380 48372 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 29092 22176 29144 22228
rect 31576 22219 31628 22228
rect 31576 22185 31585 22219
rect 31585 22185 31619 22219
rect 31619 22185 31628 22219
rect 31576 22176 31628 22185
rect 37464 22219 37516 22228
rect 37464 22185 37473 22219
rect 37473 22185 37507 22219
rect 37507 22185 37516 22219
rect 37464 22176 37516 22185
rect 44364 22176 44416 22228
rect 47308 22219 47360 22228
rect 47308 22185 47317 22219
rect 47317 22185 47351 22219
rect 47351 22185 47360 22219
rect 47308 22176 47360 22185
rect 47952 22176 48004 22228
rect 48136 22176 48188 22228
rect 29092 22040 29144 22092
rect 28080 21972 28132 22024
rect 33232 22108 33284 22160
rect 34060 22108 34112 22160
rect 34704 22108 34756 22160
rect 35624 22040 35676 22092
rect 46756 22108 46808 22160
rect 48320 22108 48372 22160
rect 37832 22083 37884 22092
rect 37832 22049 37841 22083
rect 37841 22049 37875 22083
rect 37875 22049 37884 22083
rect 37832 22040 37884 22049
rect 30012 21972 30064 22024
rect 30472 22015 30524 22024
rect 30472 21981 30506 22015
rect 30506 21981 30524 22015
rect 30472 21972 30524 21981
rect 35256 22015 35308 22024
rect 35256 21981 35265 22015
rect 35265 21981 35299 22015
rect 35299 21981 35308 22015
rect 35256 21972 35308 21981
rect 37740 22015 37792 22024
rect 30104 21904 30156 21956
rect 27620 21836 27672 21888
rect 28816 21836 28868 21888
rect 37740 21981 37749 22015
rect 37749 21981 37783 22015
rect 37783 21981 37792 22015
rect 37740 21972 37792 21981
rect 38660 21972 38712 22024
rect 44824 22015 44876 22024
rect 44824 21981 44833 22015
rect 44833 21981 44867 22015
rect 44867 21981 44876 22015
rect 44824 21972 44876 21981
rect 45744 22015 45796 22024
rect 45744 21981 45753 22015
rect 45753 21981 45787 22015
rect 45787 21981 45796 22015
rect 45744 21972 45796 21981
rect 37464 21947 37516 21956
rect 37464 21913 37473 21947
rect 37473 21913 37507 21947
rect 37507 21913 37516 21947
rect 37464 21904 37516 21913
rect 36544 21836 36596 21888
rect 37280 21879 37332 21888
rect 37280 21845 37289 21879
rect 37289 21845 37323 21879
rect 37323 21845 37332 21879
rect 37280 21836 37332 21845
rect 39212 21879 39264 21888
rect 39212 21845 39221 21879
rect 39221 21845 39255 21879
rect 39255 21845 39264 21879
rect 39212 21836 39264 21845
rect 46204 21836 46256 21888
rect 46664 22015 46716 22024
rect 46664 21981 46673 22015
rect 46673 21981 46707 22015
rect 46707 21981 46716 22015
rect 46664 21972 46716 21981
rect 47400 22040 47452 22092
rect 48872 22083 48924 22092
rect 48872 22049 48881 22083
rect 48881 22049 48915 22083
rect 48915 22049 48924 22083
rect 48872 22040 48924 22049
rect 48964 22040 49016 22092
rect 46940 21972 46992 22024
rect 47308 21904 47360 21956
rect 47492 22015 47544 22024
rect 47492 21981 47501 22015
rect 47501 21981 47535 22015
rect 47535 21981 47544 22015
rect 47492 21972 47544 21981
rect 47676 22015 47728 22024
rect 47676 21981 47685 22015
rect 47685 21981 47719 22015
rect 47719 21981 47728 22015
rect 47676 21972 47728 21981
rect 48228 22015 48280 22024
rect 48228 21981 48237 22015
rect 48237 21981 48271 22015
rect 48271 21981 48280 22015
rect 48228 21972 48280 21981
rect 48320 22015 48372 22024
rect 48320 21981 48329 22015
rect 48329 21981 48363 22015
rect 48363 21981 48372 22015
rect 48320 21972 48372 21981
rect 49608 22015 49660 22024
rect 49608 21981 49617 22015
rect 49617 21981 49651 22015
rect 49651 21981 49660 22015
rect 49608 21972 49660 21981
rect 49700 21972 49752 22024
rect 48136 21904 48188 21956
rect 48412 21947 48464 21956
rect 48412 21913 48421 21947
rect 48421 21913 48455 21947
rect 48455 21913 48464 21947
rect 48412 21904 48464 21913
rect 47032 21879 47084 21888
rect 47032 21845 47041 21879
rect 47041 21845 47075 21879
rect 47075 21845 47084 21879
rect 47032 21836 47084 21845
rect 47860 21836 47912 21888
rect 48596 21879 48648 21888
rect 48596 21845 48621 21879
rect 48621 21845 48648 21879
rect 48596 21836 48648 21845
rect 49240 21879 49292 21888
rect 49240 21845 49249 21879
rect 49249 21845 49283 21879
rect 49283 21845 49292 21879
rect 49240 21836 49292 21845
rect 49792 21836 49844 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 29092 21675 29144 21684
rect 29092 21641 29101 21675
rect 29101 21641 29135 21675
rect 29135 21641 29144 21675
rect 29092 21632 29144 21641
rect 30748 21632 30800 21684
rect 31024 21675 31076 21684
rect 31024 21641 31033 21675
rect 31033 21641 31067 21675
rect 31067 21641 31076 21675
rect 31024 21632 31076 21641
rect 34060 21632 34112 21684
rect 35256 21632 35308 21684
rect 35348 21632 35400 21684
rect 940 21496 992 21548
rect 24952 21428 25004 21480
rect 26608 21564 26660 21616
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 27436 21539 27488 21548
rect 27436 21505 27445 21539
rect 27445 21505 27479 21539
rect 27479 21505 27488 21539
rect 27436 21496 27488 21505
rect 27620 21539 27672 21548
rect 27620 21505 27629 21539
rect 27629 21505 27663 21539
rect 27663 21505 27672 21539
rect 27620 21496 27672 21505
rect 28908 21564 28960 21616
rect 30012 21564 30064 21616
rect 30656 21607 30708 21616
rect 30656 21573 30665 21607
rect 30665 21573 30699 21607
rect 30699 21573 30708 21607
rect 30656 21564 30708 21573
rect 28724 21496 28776 21548
rect 29092 21496 29144 21548
rect 31760 21496 31812 21548
rect 32588 21539 32640 21548
rect 32588 21505 32622 21539
rect 32622 21505 32640 21539
rect 32588 21496 32640 21505
rect 33508 21496 33560 21548
rect 36544 21539 36596 21548
rect 36544 21505 36553 21539
rect 36553 21505 36587 21539
rect 36587 21505 36596 21539
rect 36544 21496 36596 21505
rect 36636 21539 36688 21548
rect 36636 21505 36645 21539
rect 36645 21505 36679 21539
rect 36679 21505 36688 21539
rect 36636 21496 36688 21505
rect 37464 21632 37516 21684
rect 38292 21564 38344 21616
rect 39212 21632 39264 21684
rect 33692 21403 33744 21412
rect 33692 21369 33701 21403
rect 33701 21369 33735 21403
rect 33735 21369 33744 21403
rect 33692 21360 33744 21369
rect 1768 21335 1820 21344
rect 1768 21301 1777 21335
rect 1777 21301 1811 21335
rect 1811 21301 1820 21335
rect 1768 21292 1820 21301
rect 26884 21292 26936 21344
rect 28080 21292 28132 21344
rect 30104 21335 30156 21344
rect 30104 21301 30113 21335
rect 30113 21301 30147 21335
rect 30147 21301 30156 21335
rect 30104 21292 30156 21301
rect 30380 21292 30432 21344
rect 33416 21292 33468 21344
rect 34796 21292 34848 21344
rect 36084 21292 36136 21344
rect 36912 21292 36964 21344
rect 37740 21428 37792 21480
rect 44548 21564 44600 21616
rect 42432 21539 42484 21548
rect 42432 21505 42441 21539
rect 42441 21505 42475 21539
rect 42475 21505 42484 21539
rect 42432 21496 42484 21505
rect 42708 21496 42760 21548
rect 42800 21496 42852 21548
rect 43628 21539 43680 21548
rect 43628 21505 43637 21539
rect 43637 21505 43671 21539
rect 43671 21505 43680 21539
rect 43628 21496 43680 21505
rect 45744 21564 45796 21616
rect 46204 21564 46256 21616
rect 46480 21607 46532 21616
rect 46480 21573 46489 21607
rect 46489 21573 46523 21607
rect 46523 21573 46532 21607
rect 46480 21564 46532 21573
rect 46572 21607 46624 21616
rect 46572 21573 46581 21607
rect 46581 21573 46615 21607
rect 46615 21573 46624 21607
rect 46572 21564 46624 21573
rect 46296 21496 46348 21548
rect 46388 21539 46440 21548
rect 46388 21505 46397 21539
rect 46397 21505 46431 21539
rect 46431 21505 46440 21539
rect 46388 21496 46440 21505
rect 46756 21632 46808 21684
rect 46940 21632 46992 21684
rect 47032 21675 47084 21684
rect 47032 21641 47041 21675
rect 47041 21641 47075 21675
rect 47075 21641 47084 21675
rect 47032 21632 47084 21641
rect 47032 21496 47084 21548
rect 47308 21564 47360 21616
rect 47860 21675 47912 21684
rect 47860 21641 47869 21675
rect 47869 21641 47903 21675
rect 47903 21641 47912 21675
rect 47860 21632 47912 21641
rect 48596 21632 48648 21684
rect 49240 21632 49292 21684
rect 47768 21539 47820 21548
rect 47768 21505 47777 21539
rect 47777 21505 47811 21539
rect 47811 21505 47820 21539
rect 49792 21564 49844 21616
rect 47768 21496 47820 21505
rect 48964 21496 49016 21548
rect 46480 21428 46532 21480
rect 48228 21428 48280 21480
rect 37280 21292 37332 21344
rect 39028 21292 39080 21344
rect 42524 21335 42576 21344
rect 42524 21301 42533 21335
rect 42533 21301 42567 21335
rect 42567 21301 42576 21335
rect 42524 21292 42576 21301
rect 46388 21292 46440 21344
rect 47492 21292 47544 21344
rect 48872 21335 48924 21344
rect 48872 21301 48881 21335
rect 48881 21301 48915 21335
rect 48915 21301 48924 21335
rect 48872 21292 48924 21301
rect 49332 21471 49384 21480
rect 49332 21437 49341 21471
rect 49341 21437 49375 21471
rect 49375 21437 49384 21471
rect 49332 21428 49384 21437
rect 50068 21292 50120 21344
rect 50712 21292 50764 21344
rect 50804 21335 50856 21344
rect 50804 21301 50813 21335
rect 50813 21301 50847 21335
rect 50847 21301 50856 21335
rect 50804 21292 50856 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 27160 21088 27212 21140
rect 28724 21088 28776 21140
rect 30104 21088 30156 21140
rect 33416 21131 33468 21140
rect 33416 21097 33425 21131
rect 33425 21097 33459 21131
rect 33459 21097 33468 21131
rect 33416 21088 33468 21097
rect 33692 21088 33744 21140
rect 36912 21131 36964 21140
rect 36912 21097 36921 21131
rect 36921 21097 36955 21131
rect 36955 21097 36964 21131
rect 36912 21088 36964 21097
rect 28540 21020 28592 21072
rect 27436 20952 27488 21004
rect 26792 20927 26844 20936
rect 26792 20893 26801 20927
rect 26801 20893 26835 20927
rect 26835 20893 26844 20927
rect 26792 20884 26844 20893
rect 26884 20927 26936 20936
rect 26884 20893 26893 20927
rect 26893 20893 26927 20927
rect 26927 20893 26936 20927
rect 26884 20884 26936 20893
rect 26516 20816 26568 20868
rect 25780 20748 25832 20800
rect 27160 20927 27212 20936
rect 27160 20893 27169 20927
rect 27169 20893 27203 20927
rect 27203 20893 27212 20927
rect 27160 20884 27212 20893
rect 27804 20884 27856 20936
rect 28816 20884 28868 20936
rect 32956 20952 33008 21004
rect 29368 20816 29420 20868
rect 31760 20884 31812 20936
rect 33232 20884 33284 20936
rect 33600 20927 33652 20936
rect 33600 20893 33609 20927
rect 33609 20893 33643 20927
rect 33643 20893 33652 20927
rect 33600 20884 33652 20893
rect 34704 20995 34756 21004
rect 34704 20961 34713 20995
rect 34713 20961 34747 20995
rect 34747 20961 34756 20995
rect 34704 20952 34756 20961
rect 34796 20884 34848 20936
rect 38660 21020 38712 21072
rect 32220 20748 32272 20800
rect 36268 20816 36320 20868
rect 36544 20816 36596 20868
rect 38292 20927 38344 20936
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 38292 20884 38344 20893
rect 39028 20927 39080 20936
rect 39028 20893 39037 20927
rect 39037 20893 39071 20927
rect 39071 20893 39080 20927
rect 39028 20884 39080 20893
rect 40040 21088 40092 21140
rect 42524 21088 42576 21140
rect 44548 21131 44600 21140
rect 44548 21097 44557 21131
rect 44557 21097 44591 21131
rect 44591 21097 44600 21131
rect 44548 21088 44600 21097
rect 45744 21088 45796 21140
rect 46204 21131 46256 21140
rect 46204 21097 46213 21131
rect 46213 21097 46247 21131
rect 46247 21097 46256 21131
rect 46204 21088 46256 21097
rect 39764 21020 39816 21072
rect 38016 20859 38068 20868
rect 38016 20825 38025 20859
rect 38025 20825 38059 20859
rect 38059 20825 38068 20859
rect 38016 20816 38068 20825
rect 33324 20748 33376 20800
rect 33784 20791 33836 20800
rect 33784 20757 33793 20791
rect 33793 20757 33827 20791
rect 33827 20757 33836 20791
rect 33784 20748 33836 20757
rect 34060 20791 34112 20800
rect 34060 20757 34069 20791
rect 34069 20757 34103 20791
rect 34103 20757 34112 20791
rect 34060 20748 34112 20757
rect 36084 20791 36136 20800
rect 36084 20757 36093 20791
rect 36093 20757 36127 20791
rect 36127 20757 36136 20791
rect 36084 20748 36136 20757
rect 37924 20748 37976 20800
rect 38292 20748 38344 20800
rect 38752 20859 38804 20868
rect 38752 20825 38761 20859
rect 38761 20825 38795 20859
rect 38795 20825 38804 20859
rect 38752 20816 38804 20825
rect 38936 20791 38988 20800
rect 38936 20757 38945 20791
rect 38945 20757 38979 20791
rect 38979 20757 38988 20791
rect 38936 20748 38988 20757
rect 39672 20927 39724 20936
rect 39672 20893 39681 20927
rect 39681 20893 39715 20927
rect 39715 20893 39724 20927
rect 39672 20884 39724 20893
rect 46572 21088 46624 21140
rect 47308 21088 47360 21140
rect 41328 20927 41380 20936
rect 41328 20893 41337 20927
rect 41337 20893 41371 20927
rect 41371 20893 41380 20927
rect 41328 20884 41380 20893
rect 42340 20884 42392 20936
rect 44088 20927 44140 20936
rect 44088 20893 44097 20927
rect 44097 20893 44131 20927
rect 44131 20893 44140 20927
rect 44088 20884 44140 20893
rect 44456 20927 44508 20936
rect 44456 20893 44465 20927
rect 44465 20893 44499 20927
rect 44499 20893 44508 20927
rect 44456 20884 44508 20893
rect 45284 20884 45336 20936
rect 46296 20952 46348 21004
rect 46204 20816 46256 20868
rect 47584 20995 47636 21004
rect 46664 20927 46716 20936
rect 46664 20893 46673 20927
rect 46673 20893 46707 20927
rect 46707 20893 46716 20927
rect 46664 20884 46716 20893
rect 47584 20961 47593 20995
rect 47593 20961 47627 20995
rect 47627 20961 47636 20995
rect 47584 20952 47636 20961
rect 48320 21088 48372 21140
rect 48780 21088 48832 21140
rect 48964 21088 49016 21140
rect 49332 21088 49384 21140
rect 50804 21020 50856 21072
rect 48872 20952 48924 21004
rect 49700 20952 49752 21004
rect 50712 20952 50764 21004
rect 39580 20748 39632 20800
rect 40316 20748 40368 20800
rect 40408 20748 40460 20800
rect 42340 20748 42392 20800
rect 44180 20748 44232 20800
rect 48596 20859 48648 20868
rect 48596 20825 48605 20859
rect 48605 20825 48639 20859
rect 48639 20825 48648 20859
rect 48596 20816 48648 20825
rect 46572 20748 46624 20800
rect 46940 20791 46992 20800
rect 46940 20757 46949 20791
rect 46949 20757 46983 20791
rect 46983 20757 46992 20791
rect 46940 20748 46992 20757
rect 47768 20748 47820 20800
rect 47860 20791 47912 20800
rect 47860 20757 47869 20791
rect 47869 20757 47903 20791
rect 47903 20757 47912 20791
rect 47860 20748 47912 20757
rect 48504 20748 48556 20800
rect 48872 20791 48924 20800
rect 48872 20757 48881 20791
rect 48881 20757 48915 20791
rect 48915 20757 48924 20791
rect 48872 20748 48924 20757
rect 49148 20748 49200 20800
rect 50436 20927 50488 20936
rect 50436 20893 50445 20927
rect 50445 20893 50479 20927
rect 50479 20893 50488 20927
rect 50436 20884 50488 20893
rect 49792 20816 49844 20868
rect 49884 20816 49936 20868
rect 49976 20816 50028 20868
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 26792 20587 26844 20596
rect 26792 20553 26801 20587
rect 26801 20553 26835 20587
rect 26835 20553 26844 20587
rect 26792 20544 26844 20553
rect 28080 20587 28132 20596
rect 28080 20553 28089 20587
rect 28089 20553 28123 20587
rect 28123 20553 28132 20587
rect 28080 20544 28132 20553
rect 25780 20476 25832 20528
rect 33232 20544 33284 20596
rect 38752 20544 38804 20596
rect 39856 20544 39908 20596
rect 32036 20476 32088 20528
rect 34704 20476 34756 20528
rect 24952 20451 25004 20460
rect 24952 20417 24961 20451
rect 24961 20417 24995 20451
rect 24995 20417 25004 20451
rect 24952 20408 25004 20417
rect 26608 20451 26660 20460
rect 26608 20417 26617 20451
rect 26617 20417 26651 20451
rect 26651 20417 26660 20451
rect 26608 20408 26660 20417
rect 28540 20451 28592 20460
rect 28540 20417 28549 20451
rect 28549 20417 28583 20451
rect 28583 20417 28592 20451
rect 28540 20408 28592 20417
rect 28724 20451 28776 20460
rect 28724 20417 28733 20451
rect 28733 20417 28767 20451
rect 28767 20417 28776 20451
rect 28724 20408 28776 20417
rect 28908 20408 28960 20460
rect 29092 20451 29144 20460
rect 29092 20417 29126 20451
rect 29126 20417 29144 20451
rect 29092 20408 29144 20417
rect 30564 20451 30616 20460
rect 30564 20417 30598 20451
rect 30598 20417 30616 20451
rect 30564 20408 30616 20417
rect 32220 20451 32272 20460
rect 32220 20417 32229 20451
rect 32229 20417 32263 20451
rect 32263 20417 32272 20451
rect 32220 20408 32272 20417
rect 33324 20451 33376 20460
rect 33324 20417 33333 20451
rect 33333 20417 33367 20451
rect 33367 20417 33376 20451
rect 33324 20408 33376 20417
rect 34520 20408 34572 20460
rect 36084 20408 36136 20460
rect 36268 20451 36320 20460
rect 36268 20417 36277 20451
rect 36277 20417 36311 20451
rect 36311 20417 36320 20451
rect 36268 20408 36320 20417
rect 27160 20340 27212 20392
rect 27620 20340 27672 20392
rect 30012 20340 30064 20392
rect 38660 20408 38712 20460
rect 38936 20476 38988 20528
rect 40408 20476 40460 20528
rect 42340 20544 42392 20596
rect 42708 20544 42760 20596
rect 45284 20587 45336 20596
rect 45284 20553 45293 20587
rect 45293 20553 45327 20587
rect 45327 20553 45336 20587
rect 45284 20544 45336 20553
rect 46756 20544 46808 20596
rect 38016 20340 38068 20392
rect 39764 20408 39816 20460
rect 27620 20247 27672 20256
rect 27620 20213 27629 20247
rect 27629 20213 27663 20247
rect 27663 20213 27672 20247
rect 27620 20204 27672 20213
rect 28080 20247 28132 20256
rect 28080 20213 28089 20247
rect 28089 20213 28123 20247
rect 28123 20213 28132 20247
rect 28080 20204 28132 20213
rect 29736 20204 29788 20256
rect 30012 20204 30064 20256
rect 30196 20247 30248 20256
rect 30196 20213 30205 20247
rect 30205 20213 30239 20247
rect 30239 20213 30248 20247
rect 30196 20204 30248 20213
rect 30656 20204 30708 20256
rect 31668 20247 31720 20256
rect 31668 20213 31677 20247
rect 31677 20213 31711 20247
rect 31711 20213 31720 20247
rect 31668 20204 31720 20213
rect 33324 20204 33376 20256
rect 33600 20272 33652 20324
rect 37372 20272 37424 20324
rect 40040 20340 40092 20392
rect 40500 20408 40552 20460
rect 41328 20476 41380 20528
rect 40868 20451 40920 20460
rect 40868 20417 40877 20451
rect 40877 20417 40911 20451
rect 40911 20417 40920 20451
rect 40868 20408 40920 20417
rect 42432 20408 42484 20460
rect 43536 20476 43588 20528
rect 46112 20408 46164 20460
rect 46480 20408 46532 20460
rect 47308 20476 47360 20528
rect 49148 20544 49200 20596
rect 49976 20544 50028 20596
rect 47768 20408 47820 20460
rect 48320 20408 48372 20460
rect 50160 20476 50212 20528
rect 41604 20383 41656 20392
rect 41604 20349 41613 20383
rect 41613 20349 41647 20383
rect 41647 20349 41656 20383
rect 41604 20340 41656 20349
rect 42800 20383 42852 20392
rect 42800 20349 42809 20383
rect 42809 20349 42843 20383
rect 42843 20349 42852 20383
rect 42800 20340 42852 20349
rect 33876 20204 33928 20256
rect 36268 20204 36320 20256
rect 37924 20204 37976 20256
rect 38660 20204 38712 20256
rect 38844 20204 38896 20256
rect 40684 20247 40736 20256
rect 40684 20213 40693 20247
rect 40693 20213 40727 20247
rect 40727 20213 40736 20247
rect 40684 20204 40736 20213
rect 41512 20247 41564 20256
rect 41512 20213 41521 20247
rect 41521 20213 41555 20247
rect 41555 20213 41564 20247
rect 41512 20204 41564 20213
rect 44272 20247 44324 20256
rect 44272 20213 44281 20247
rect 44281 20213 44315 20247
rect 44315 20213 44324 20247
rect 44272 20204 44324 20213
rect 44456 20204 44508 20256
rect 46940 20247 46992 20256
rect 46940 20213 46949 20247
rect 46949 20213 46983 20247
rect 46983 20213 46992 20247
rect 46940 20204 46992 20213
rect 47032 20204 47084 20256
rect 47492 20204 47544 20256
rect 47860 20272 47912 20324
rect 48504 20340 48556 20392
rect 49148 20408 49200 20460
rect 49884 20408 49936 20460
rect 48780 20383 48832 20392
rect 48780 20349 48789 20383
rect 48789 20349 48823 20383
rect 48823 20349 48832 20383
rect 48780 20340 48832 20349
rect 50804 20408 50856 20460
rect 47952 20247 48004 20256
rect 47952 20213 47961 20247
rect 47961 20213 47995 20247
rect 47995 20213 48004 20247
rect 47952 20204 48004 20213
rect 48596 20204 48648 20256
rect 49608 20204 49660 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 26516 20043 26568 20052
rect 26516 20009 26525 20043
rect 26525 20009 26559 20043
rect 26559 20009 26568 20043
rect 26516 20000 26568 20009
rect 27620 20000 27672 20052
rect 27804 20000 27856 20052
rect 30012 20000 30064 20052
rect 30564 20000 30616 20052
rect 32036 20043 32088 20052
rect 26700 19864 26752 19916
rect 28632 19864 28684 19916
rect 28908 19864 28960 19916
rect 32036 20009 32045 20043
rect 32045 20009 32079 20043
rect 32079 20009 32088 20043
rect 32036 20000 32088 20009
rect 32588 20043 32640 20052
rect 32588 20009 32597 20043
rect 32597 20009 32631 20043
rect 32631 20009 32640 20043
rect 32588 20000 32640 20009
rect 31668 19932 31720 19984
rect 27160 19839 27212 19848
rect 27160 19805 27169 19839
rect 27169 19805 27203 19839
rect 27203 19805 27212 19839
rect 27160 19796 27212 19805
rect 27252 19839 27304 19848
rect 27252 19805 27261 19839
rect 27261 19805 27295 19839
rect 27295 19805 27304 19839
rect 27252 19796 27304 19805
rect 27528 19796 27580 19848
rect 27620 19796 27672 19848
rect 28724 19796 28776 19848
rect 26608 19728 26660 19780
rect 28448 19771 28500 19780
rect 28448 19737 28457 19771
rect 28457 19737 28491 19771
rect 28491 19737 28500 19771
rect 28448 19728 28500 19737
rect 28632 19728 28684 19780
rect 29644 19796 29696 19848
rect 30196 19796 30248 19848
rect 32220 19796 32272 19848
rect 33324 19932 33376 19984
rect 33508 19932 33560 19984
rect 33692 19975 33744 19984
rect 33692 19941 33701 19975
rect 33701 19941 33735 19975
rect 33735 19941 33744 19975
rect 33692 19932 33744 19941
rect 33140 19839 33192 19848
rect 33140 19805 33149 19839
rect 33149 19805 33183 19839
rect 33183 19805 33192 19839
rect 33140 19796 33192 19805
rect 33508 19796 33560 19848
rect 33600 19839 33652 19848
rect 33600 19805 33609 19839
rect 33609 19805 33643 19839
rect 33643 19805 33652 19839
rect 33600 19796 33652 19805
rect 33692 19796 33744 19848
rect 33968 19796 34020 19848
rect 34336 19796 34388 19848
rect 37372 20000 37424 20052
rect 34704 19864 34756 19916
rect 37832 20000 37884 20052
rect 38660 19932 38712 19984
rect 38844 19975 38896 19984
rect 38844 19941 38853 19975
rect 38853 19941 38887 19975
rect 38887 19941 38896 19975
rect 38844 19932 38896 19941
rect 34612 19796 34664 19848
rect 37188 19839 37240 19848
rect 37188 19805 37197 19839
rect 37197 19805 37231 19839
rect 37231 19805 37240 19839
rect 40224 20000 40276 20052
rect 41512 20000 41564 20052
rect 42800 20000 42852 20052
rect 43536 20043 43588 20052
rect 43536 20009 43545 20043
rect 43545 20009 43579 20043
rect 43579 20009 43588 20043
rect 43536 20000 43588 20009
rect 46664 20000 46716 20052
rect 40868 19932 40920 19984
rect 43444 19932 43496 19984
rect 47492 19932 47544 19984
rect 37188 19796 37240 19805
rect 26976 19703 27028 19712
rect 26976 19669 26985 19703
rect 26985 19669 27019 19703
rect 27019 19669 27028 19703
rect 26976 19660 27028 19669
rect 27436 19660 27488 19712
rect 27804 19660 27856 19712
rect 34520 19728 34572 19780
rect 36636 19728 36688 19780
rect 37280 19728 37332 19780
rect 29736 19703 29788 19712
rect 29736 19669 29761 19703
rect 29761 19669 29788 19703
rect 29736 19660 29788 19669
rect 29920 19703 29972 19712
rect 29920 19669 29929 19703
rect 29929 19669 29963 19703
rect 29963 19669 29972 19703
rect 29920 19660 29972 19669
rect 33784 19660 33836 19712
rect 34796 19703 34848 19712
rect 34796 19669 34805 19703
rect 34805 19669 34839 19703
rect 34839 19669 34848 19703
rect 34796 19660 34848 19669
rect 36728 19660 36780 19712
rect 37004 19703 37056 19712
rect 37004 19669 37013 19703
rect 37013 19669 37047 19703
rect 37047 19669 37056 19703
rect 37004 19660 37056 19669
rect 40684 19796 40736 19848
rect 38384 19728 38436 19780
rect 40316 19660 40368 19712
rect 42616 19839 42668 19848
rect 42616 19805 42625 19839
rect 42625 19805 42659 19839
rect 42659 19805 42668 19839
rect 42616 19796 42668 19805
rect 44180 19864 44232 19916
rect 46020 19864 46072 19916
rect 44824 19839 44876 19848
rect 44824 19805 44833 19839
rect 44833 19805 44867 19839
rect 44867 19805 44876 19839
rect 44824 19796 44876 19805
rect 46480 19728 46532 19780
rect 46664 19839 46716 19848
rect 46664 19805 46673 19839
rect 46673 19805 46707 19839
rect 46707 19805 46716 19839
rect 46664 19796 46716 19805
rect 47032 19796 47084 19848
rect 47124 19839 47176 19848
rect 47124 19805 47133 19839
rect 47133 19805 47167 19839
rect 47167 19805 47176 19839
rect 47124 19796 47176 19805
rect 48504 20000 48556 20052
rect 49976 20000 50028 20052
rect 50528 20000 50580 20052
rect 48320 19932 48372 19984
rect 47952 19864 48004 19916
rect 50528 19864 50580 19916
rect 47400 19728 47452 19780
rect 45468 19660 45520 19712
rect 46388 19703 46440 19712
rect 46388 19669 46397 19703
rect 46397 19669 46431 19703
rect 46431 19669 46440 19703
rect 46388 19660 46440 19669
rect 49608 19839 49660 19848
rect 49608 19805 49617 19839
rect 49617 19805 49651 19839
rect 49651 19805 49660 19839
rect 49608 19796 49660 19805
rect 49976 19839 50028 19848
rect 49976 19805 49985 19839
rect 49985 19805 50019 19839
rect 50019 19805 50028 19839
rect 49976 19796 50028 19805
rect 50068 19796 50120 19848
rect 68468 19839 68520 19848
rect 68468 19805 68477 19839
rect 68477 19805 68511 19839
rect 68511 19805 68520 19839
rect 68468 19796 68520 19805
rect 49700 19771 49752 19780
rect 49700 19737 49709 19771
rect 49709 19737 49743 19771
rect 49743 19737 49752 19771
rect 49700 19728 49752 19737
rect 49792 19728 49844 19780
rect 51080 19728 51132 19780
rect 50160 19660 50212 19712
rect 50620 19660 50672 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 26976 19456 27028 19508
rect 27712 19456 27764 19508
rect 29092 19456 29144 19508
rect 32956 19456 33008 19508
rect 33508 19456 33560 19508
rect 34060 19456 34112 19508
rect 34796 19456 34848 19508
rect 27344 19320 27396 19372
rect 31852 19431 31904 19440
rect 31852 19397 31861 19431
rect 31861 19397 31895 19431
rect 31895 19397 31904 19431
rect 31852 19388 31904 19397
rect 32220 19388 32272 19440
rect 33600 19388 33652 19440
rect 33968 19431 34020 19440
rect 33968 19397 33977 19431
rect 33977 19397 34011 19431
rect 34011 19397 34020 19431
rect 33968 19388 34020 19397
rect 27804 19320 27856 19372
rect 28632 19320 28684 19372
rect 28724 19363 28776 19372
rect 28724 19329 28733 19363
rect 28733 19329 28767 19363
rect 28767 19329 28776 19363
rect 28724 19320 28776 19329
rect 29920 19320 29972 19372
rect 31484 19320 31536 19372
rect 31576 19363 31628 19372
rect 31576 19329 31585 19363
rect 31585 19329 31619 19363
rect 31619 19329 31628 19363
rect 31576 19320 31628 19329
rect 31760 19320 31812 19372
rect 28908 19252 28960 19304
rect 33692 19320 33744 19372
rect 34060 19320 34112 19372
rect 36636 19499 36688 19508
rect 36636 19465 36645 19499
rect 36645 19465 36679 19499
rect 36679 19465 36688 19499
rect 36636 19456 36688 19465
rect 40500 19456 40552 19508
rect 27620 19184 27672 19236
rect 28632 19184 28684 19236
rect 26240 19159 26292 19168
rect 26240 19125 26249 19159
rect 26249 19125 26283 19159
rect 26283 19125 26292 19159
rect 26240 19116 26292 19125
rect 27436 19159 27488 19168
rect 27436 19125 27445 19159
rect 27445 19125 27479 19159
rect 27479 19125 27488 19159
rect 27436 19116 27488 19125
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 33324 19184 33376 19236
rect 32864 19116 32916 19168
rect 34152 19159 34204 19168
rect 34152 19125 34161 19159
rect 34161 19125 34195 19159
rect 34195 19125 34204 19159
rect 34152 19116 34204 19125
rect 36084 19295 36136 19304
rect 36084 19261 36093 19295
rect 36093 19261 36127 19295
rect 36127 19261 36136 19295
rect 36084 19252 36136 19261
rect 36912 19252 36964 19304
rect 37464 19252 37516 19304
rect 41236 19388 41288 19440
rect 42616 19456 42668 19508
rect 44456 19456 44508 19508
rect 44824 19456 44876 19508
rect 46664 19456 46716 19508
rect 47032 19456 47084 19508
rect 47308 19456 47360 19508
rect 39856 19320 39908 19372
rect 40408 19320 40460 19372
rect 40868 19320 40920 19372
rect 41328 19363 41380 19372
rect 41328 19329 41337 19363
rect 41337 19329 41371 19363
rect 41371 19329 41380 19363
rect 41328 19320 41380 19329
rect 43444 19388 43496 19440
rect 43628 19388 43680 19440
rect 43720 19320 43772 19372
rect 42524 19295 42576 19304
rect 42524 19261 42533 19295
rect 42533 19261 42567 19295
rect 42567 19261 42576 19295
rect 42524 19252 42576 19261
rect 43536 19295 43588 19304
rect 43536 19261 43545 19295
rect 43545 19261 43579 19295
rect 43579 19261 43588 19295
rect 43536 19252 43588 19261
rect 44088 19252 44140 19304
rect 46848 19320 46900 19372
rect 46940 19363 46992 19372
rect 46940 19329 46949 19363
rect 46949 19329 46983 19363
rect 46983 19329 46992 19363
rect 46940 19320 46992 19329
rect 50160 19499 50212 19508
rect 50160 19465 50169 19499
rect 50169 19465 50203 19499
rect 50203 19465 50212 19499
rect 50160 19456 50212 19465
rect 48780 19388 48832 19440
rect 47308 19363 47360 19372
rect 47308 19329 47317 19363
rect 47317 19329 47351 19363
rect 47351 19329 47360 19363
rect 47308 19320 47360 19329
rect 47768 19363 47820 19372
rect 47768 19329 47777 19363
rect 47777 19329 47811 19363
rect 47811 19329 47820 19363
rect 47768 19320 47820 19329
rect 49792 19320 49844 19372
rect 49976 19320 50028 19372
rect 36360 19184 36412 19236
rect 44272 19184 44324 19236
rect 46388 19252 46440 19304
rect 46572 19252 46624 19304
rect 46204 19184 46256 19236
rect 50804 19252 50856 19304
rect 35348 19116 35400 19168
rect 36176 19116 36228 19168
rect 38292 19116 38344 19168
rect 39764 19159 39816 19168
rect 39764 19125 39773 19159
rect 39773 19125 39807 19159
rect 39807 19125 39816 19159
rect 39764 19116 39816 19125
rect 42616 19159 42668 19168
rect 42616 19125 42625 19159
rect 42625 19125 42659 19159
rect 42659 19125 42668 19159
rect 42616 19116 42668 19125
rect 43536 19116 43588 19168
rect 47216 19159 47268 19168
rect 47216 19125 47225 19159
rect 47225 19125 47259 19159
rect 47259 19125 47268 19159
rect 47216 19116 47268 19125
rect 47400 19116 47452 19168
rect 47952 19159 48004 19168
rect 47952 19125 47961 19159
rect 47961 19125 47995 19159
rect 47995 19125 48004 19159
rect 47952 19116 48004 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 27252 18912 27304 18964
rect 28080 18912 28132 18964
rect 31852 18912 31904 18964
rect 32864 18955 32916 18964
rect 32864 18921 32873 18955
rect 32873 18921 32907 18955
rect 32907 18921 32916 18955
rect 32864 18912 32916 18921
rect 34060 18912 34112 18964
rect 34612 18912 34664 18964
rect 36084 18912 36136 18964
rect 36820 18955 36872 18964
rect 36820 18921 36829 18955
rect 36829 18921 36863 18955
rect 36863 18921 36872 18955
rect 36820 18912 36872 18921
rect 41144 18912 41196 18964
rect 45008 18912 45060 18964
rect 46112 18955 46164 18964
rect 46112 18921 46121 18955
rect 46121 18921 46155 18955
rect 46155 18921 46164 18955
rect 46112 18912 46164 18921
rect 46388 18912 46440 18964
rect 33324 18819 33376 18828
rect 33324 18785 33333 18819
rect 33333 18785 33367 18819
rect 33367 18785 33376 18819
rect 33324 18776 33376 18785
rect 940 18708 992 18760
rect 25228 18708 25280 18760
rect 26240 18708 26292 18760
rect 27160 18708 27212 18760
rect 28448 18683 28500 18692
rect 28448 18649 28457 18683
rect 28457 18649 28491 18683
rect 28491 18649 28500 18683
rect 28448 18640 28500 18649
rect 29184 18683 29236 18692
rect 29184 18649 29193 18683
rect 29193 18649 29227 18683
rect 29227 18649 29236 18683
rect 33140 18751 33192 18760
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 37004 18844 37056 18896
rect 39396 18844 39448 18896
rect 39764 18844 39816 18896
rect 33140 18708 33192 18717
rect 34520 18708 34572 18760
rect 29184 18640 29236 18649
rect 30196 18640 30248 18692
rect 31392 18683 31444 18692
rect 31392 18649 31401 18683
rect 31401 18649 31435 18683
rect 31435 18649 31444 18683
rect 31392 18640 31444 18649
rect 33968 18683 34020 18692
rect 33968 18649 33977 18683
rect 33977 18649 34011 18683
rect 34011 18649 34020 18683
rect 36728 18776 36780 18828
rect 36176 18751 36228 18760
rect 36176 18717 36183 18751
rect 36183 18717 36228 18751
rect 33968 18640 34020 18649
rect 35348 18640 35400 18692
rect 36176 18708 36228 18717
rect 36268 18751 36320 18760
rect 36268 18717 36277 18751
rect 36277 18717 36311 18751
rect 36311 18717 36320 18751
rect 36268 18708 36320 18717
rect 36360 18751 36412 18760
rect 36360 18717 36369 18751
rect 36369 18717 36403 18751
rect 36403 18717 36412 18751
rect 36360 18708 36412 18717
rect 36452 18708 36504 18760
rect 37096 18727 37123 18760
rect 37123 18727 37148 18760
rect 37096 18708 37148 18727
rect 37188 18751 37240 18760
rect 37188 18717 37197 18751
rect 37197 18717 37231 18751
rect 37231 18717 37240 18751
rect 37188 18708 37240 18717
rect 37924 18751 37976 18760
rect 37924 18717 37933 18751
rect 37933 18717 37967 18751
rect 37967 18717 37976 18751
rect 37924 18708 37976 18717
rect 38384 18751 38436 18760
rect 42524 18776 42576 18828
rect 38384 18717 38398 18751
rect 38398 18717 38432 18751
rect 38432 18717 38436 18751
rect 38384 18708 38436 18717
rect 36820 18683 36872 18692
rect 36820 18649 36829 18683
rect 36829 18649 36863 18683
rect 36863 18649 36872 18683
rect 36820 18640 36872 18649
rect 27528 18572 27580 18624
rect 28908 18572 28960 18624
rect 29552 18572 29604 18624
rect 33508 18572 33560 18624
rect 33692 18572 33744 18624
rect 36728 18572 36780 18624
rect 38200 18683 38252 18692
rect 38200 18649 38209 18683
rect 38209 18649 38243 18683
rect 38243 18649 38252 18683
rect 38200 18640 38252 18649
rect 38292 18683 38344 18692
rect 38292 18649 38301 18683
rect 38301 18649 38335 18683
rect 38335 18649 38344 18683
rect 38292 18640 38344 18649
rect 38476 18640 38528 18692
rect 38660 18640 38712 18692
rect 40132 18751 40184 18760
rect 40132 18717 40141 18751
rect 40141 18717 40175 18751
rect 40175 18717 40184 18751
rect 40132 18708 40184 18717
rect 41052 18683 41104 18692
rect 41052 18649 41086 18683
rect 41086 18649 41104 18683
rect 41052 18640 41104 18649
rect 41236 18640 41288 18692
rect 43812 18819 43864 18828
rect 43812 18785 43821 18819
rect 43821 18785 43855 18819
rect 43855 18785 43864 18819
rect 43812 18776 43864 18785
rect 43444 18708 43496 18760
rect 43720 18751 43772 18760
rect 43720 18717 43729 18751
rect 43729 18717 43763 18751
rect 43763 18717 43772 18751
rect 43720 18708 43772 18717
rect 43904 18751 43956 18760
rect 43904 18717 43913 18751
rect 43913 18717 43947 18751
rect 43947 18717 43956 18751
rect 43904 18708 43956 18717
rect 44364 18751 44416 18760
rect 44364 18717 44373 18751
rect 44373 18717 44407 18751
rect 44407 18717 44416 18751
rect 44364 18708 44416 18717
rect 44088 18640 44140 18692
rect 44824 18640 44876 18692
rect 46664 18844 46716 18896
rect 47216 18912 47268 18964
rect 46756 18708 46808 18760
rect 50804 18912 50856 18964
rect 51080 18955 51132 18964
rect 51080 18921 51089 18955
rect 51089 18921 51123 18955
rect 51123 18921 51132 18955
rect 51080 18912 51132 18921
rect 37372 18572 37424 18624
rect 38752 18572 38804 18624
rect 38936 18572 38988 18624
rect 39488 18615 39540 18624
rect 39488 18581 39497 18615
rect 39497 18581 39531 18615
rect 39531 18581 39540 18615
rect 39488 18572 39540 18581
rect 41604 18572 41656 18624
rect 45008 18572 45060 18624
rect 45652 18615 45704 18624
rect 45652 18581 45661 18615
rect 45661 18581 45695 18615
rect 45695 18581 45704 18615
rect 45652 18572 45704 18581
rect 46480 18615 46532 18624
rect 46480 18581 46489 18615
rect 46489 18581 46523 18615
rect 46523 18581 46532 18615
rect 47676 18683 47728 18692
rect 47676 18649 47685 18683
rect 47685 18649 47719 18683
rect 47719 18649 47728 18683
rect 47676 18640 47728 18649
rect 48228 18640 48280 18692
rect 50620 18819 50672 18828
rect 50620 18785 50629 18819
rect 50629 18785 50663 18819
rect 50663 18785 50672 18819
rect 50620 18776 50672 18785
rect 50804 18819 50856 18828
rect 50804 18785 50813 18819
rect 50813 18785 50847 18819
rect 50847 18785 50856 18819
rect 50804 18776 50856 18785
rect 48872 18751 48924 18760
rect 48872 18717 48881 18751
rect 48881 18717 48915 18751
rect 48915 18717 48924 18751
rect 48872 18708 48924 18717
rect 49700 18708 49752 18760
rect 46480 18572 46532 18581
rect 48780 18615 48832 18624
rect 48780 18581 48789 18615
rect 48789 18581 48823 18615
rect 48823 18581 48832 18615
rect 48780 18572 48832 18581
rect 48964 18572 49016 18624
rect 50160 18615 50212 18624
rect 50160 18581 50169 18615
rect 50169 18581 50203 18615
rect 50203 18581 50212 18615
rect 50160 18572 50212 18581
rect 50712 18572 50764 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 26700 18368 26752 18420
rect 31852 18368 31904 18420
rect 27252 18232 27304 18284
rect 29644 18343 29696 18352
rect 29644 18309 29653 18343
rect 29653 18309 29687 18343
rect 29687 18309 29696 18343
rect 29644 18300 29696 18309
rect 30012 18343 30064 18352
rect 30012 18309 30021 18343
rect 30021 18309 30055 18343
rect 30055 18309 30064 18343
rect 30012 18300 30064 18309
rect 30196 18300 30248 18352
rect 31760 18300 31812 18352
rect 29552 18232 29604 18284
rect 27804 18096 27856 18148
rect 28356 18096 28408 18148
rect 27988 18028 28040 18080
rect 31576 18275 31628 18284
rect 31576 18241 31585 18275
rect 31585 18241 31619 18275
rect 31619 18241 31628 18275
rect 31576 18232 31628 18241
rect 32036 18164 32088 18216
rect 32128 18207 32180 18216
rect 32128 18173 32137 18207
rect 32137 18173 32171 18207
rect 32171 18173 32180 18207
rect 32128 18164 32180 18173
rect 33692 18411 33744 18420
rect 33692 18377 33701 18411
rect 33701 18377 33735 18411
rect 33735 18377 33744 18411
rect 33692 18368 33744 18377
rect 34152 18368 34204 18420
rect 32956 18300 33008 18352
rect 33600 18300 33652 18352
rect 32220 18096 32272 18148
rect 31300 18071 31352 18080
rect 31300 18037 31309 18071
rect 31309 18037 31343 18071
rect 31343 18037 31352 18071
rect 31300 18028 31352 18037
rect 31576 18028 31628 18080
rect 32404 18028 32456 18080
rect 32864 18071 32916 18080
rect 32864 18037 32873 18071
rect 32873 18037 32907 18071
rect 32907 18037 32916 18071
rect 32864 18028 32916 18037
rect 33324 18275 33376 18284
rect 33324 18241 33333 18275
rect 33333 18241 33367 18275
rect 33367 18241 33376 18275
rect 33324 18232 33376 18241
rect 35348 18232 35400 18284
rect 35808 18232 35860 18284
rect 38200 18368 38252 18420
rect 38292 18368 38344 18420
rect 37004 18300 37056 18352
rect 37832 18275 37884 18284
rect 34704 18164 34756 18216
rect 37832 18241 37841 18275
rect 37841 18241 37875 18275
rect 37875 18241 37884 18275
rect 37832 18232 37884 18241
rect 37096 18207 37148 18216
rect 37096 18173 37105 18207
rect 37105 18173 37139 18207
rect 37139 18173 37148 18207
rect 37096 18164 37148 18173
rect 37280 18164 37332 18216
rect 34152 18139 34204 18148
rect 34152 18105 34161 18139
rect 34161 18105 34195 18139
rect 34195 18105 34204 18139
rect 34152 18096 34204 18105
rect 37188 18096 37240 18148
rect 38384 18232 38436 18284
rect 38936 18368 38988 18420
rect 41052 18368 41104 18420
rect 42616 18368 42668 18420
rect 44364 18368 44416 18420
rect 39948 18300 40000 18352
rect 38936 18232 38988 18284
rect 41144 18232 41196 18284
rect 41236 18275 41288 18284
rect 41236 18241 41245 18275
rect 41245 18241 41279 18275
rect 41279 18241 41288 18275
rect 41236 18232 41288 18241
rect 41328 18275 41380 18284
rect 41328 18241 41337 18275
rect 41337 18241 41371 18275
rect 41371 18241 41380 18275
rect 41328 18232 41380 18241
rect 44364 18275 44416 18284
rect 44364 18241 44373 18275
rect 44373 18241 44407 18275
rect 44407 18241 44416 18275
rect 44364 18232 44416 18241
rect 44824 18232 44876 18284
rect 45284 18275 45336 18284
rect 45284 18241 45293 18275
rect 45293 18241 45327 18275
rect 45327 18241 45336 18275
rect 45284 18232 45336 18241
rect 36360 18028 36412 18080
rect 36912 18028 36964 18080
rect 37280 18028 37332 18080
rect 38200 18096 38252 18148
rect 38844 18096 38896 18148
rect 38568 18028 38620 18080
rect 43904 18096 43956 18148
rect 45468 18275 45520 18284
rect 45468 18241 45477 18275
rect 45477 18241 45511 18275
rect 45511 18241 45520 18275
rect 45468 18232 45520 18241
rect 45652 18368 45704 18420
rect 46572 18411 46624 18420
rect 46572 18377 46581 18411
rect 46581 18377 46615 18411
rect 46615 18377 46624 18411
rect 46572 18368 46624 18377
rect 46848 18300 46900 18352
rect 47400 18368 47452 18420
rect 47584 18368 47636 18420
rect 46480 18275 46532 18284
rect 45652 18096 45704 18148
rect 44088 18028 44140 18080
rect 46480 18241 46489 18275
rect 46489 18241 46523 18275
rect 46523 18241 46532 18275
rect 46480 18232 46532 18241
rect 46664 18275 46716 18284
rect 46664 18241 46673 18275
rect 46673 18241 46707 18275
rect 46707 18241 46716 18275
rect 46664 18232 46716 18241
rect 46756 18232 46808 18284
rect 47124 18164 47176 18216
rect 47768 18300 47820 18352
rect 47584 18275 47636 18284
rect 47584 18241 47593 18275
rect 47593 18241 47627 18275
rect 47627 18241 47636 18275
rect 47584 18232 47636 18241
rect 48964 18232 49016 18284
rect 50068 18368 50120 18420
rect 50804 18368 50856 18420
rect 51080 18232 51132 18284
rect 47952 18164 48004 18216
rect 48872 18164 48924 18216
rect 49976 18207 50028 18216
rect 49976 18173 49985 18207
rect 49985 18173 50019 18207
rect 50019 18173 50028 18207
rect 49976 18164 50028 18173
rect 46388 18071 46440 18080
rect 46388 18037 46397 18071
rect 46397 18037 46431 18071
rect 46431 18037 46440 18071
rect 46388 18028 46440 18037
rect 46940 18028 46992 18080
rect 47676 18028 47728 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 1768 17824 1820 17876
rect 27252 17824 27304 17876
rect 27804 17731 27856 17740
rect 27804 17697 27813 17731
rect 27813 17697 27847 17731
rect 27847 17697 27856 17731
rect 27804 17688 27856 17697
rect 25228 17620 25280 17672
rect 27988 17620 28040 17672
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 29736 17824 29788 17876
rect 31392 17824 31444 17876
rect 32128 17867 32180 17876
rect 32128 17833 32137 17867
rect 32137 17833 32171 17867
rect 32171 17833 32180 17867
rect 32128 17824 32180 17833
rect 32220 17867 32272 17876
rect 32220 17833 32229 17867
rect 32229 17833 32263 17867
rect 32263 17833 32272 17867
rect 32220 17824 32272 17833
rect 34060 17824 34112 17876
rect 34152 17824 34204 17876
rect 35808 17867 35860 17876
rect 35808 17833 35817 17867
rect 35817 17833 35851 17867
rect 35851 17833 35860 17867
rect 35808 17824 35860 17833
rect 36452 17824 36504 17876
rect 32036 17756 32088 17808
rect 29276 17552 29328 17604
rect 29736 17595 29788 17604
rect 29736 17561 29745 17595
rect 29745 17561 29779 17595
rect 29779 17561 29788 17595
rect 29736 17552 29788 17561
rect 30196 17552 30248 17604
rect 29368 17484 29420 17536
rect 30012 17484 30064 17536
rect 30748 17663 30800 17672
rect 30748 17629 30757 17663
rect 30757 17629 30791 17663
rect 30791 17629 30800 17663
rect 30748 17620 30800 17629
rect 31300 17620 31352 17672
rect 32404 17663 32456 17672
rect 32404 17629 32413 17663
rect 32413 17629 32447 17663
rect 32447 17629 32456 17663
rect 32404 17620 32456 17629
rect 32864 17688 32916 17740
rect 33600 17620 33652 17672
rect 33968 17620 34020 17672
rect 34428 17620 34480 17672
rect 34704 17663 34756 17672
rect 34704 17629 34713 17663
rect 34713 17629 34747 17663
rect 34747 17629 34756 17663
rect 34704 17620 34756 17629
rect 37372 17824 37424 17876
rect 37832 17824 37884 17876
rect 37188 17756 37240 17808
rect 38660 17824 38712 17876
rect 43444 17824 43496 17876
rect 44088 17824 44140 17876
rect 43720 17756 43772 17808
rect 45284 17824 45336 17876
rect 46480 17867 46532 17876
rect 46480 17833 46489 17867
rect 46489 17833 46523 17867
rect 46523 17833 46532 17867
rect 46480 17824 46532 17833
rect 46848 17824 46900 17876
rect 49976 17824 50028 17876
rect 51080 17824 51132 17876
rect 33140 17484 33192 17536
rect 33232 17527 33284 17536
rect 33232 17493 33241 17527
rect 33241 17493 33275 17527
rect 33275 17493 33284 17527
rect 33232 17484 33284 17493
rect 36636 17552 36688 17604
rect 36912 17620 36964 17672
rect 37188 17663 37240 17672
rect 37188 17629 37197 17663
rect 37197 17629 37231 17663
rect 37231 17629 37240 17663
rect 37188 17620 37240 17629
rect 37280 17620 37332 17672
rect 37924 17620 37976 17672
rect 36176 17484 36228 17536
rect 43812 17663 43864 17672
rect 43812 17629 43821 17663
rect 43821 17629 43855 17663
rect 43855 17629 43864 17663
rect 43812 17620 43864 17629
rect 43904 17620 43956 17672
rect 44364 17663 44416 17672
rect 44364 17629 44373 17663
rect 44373 17629 44407 17663
rect 44407 17629 44416 17663
rect 44364 17620 44416 17629
rect 44456 17620 44508 17672
rect 47584 17688 47636 17740
rect 49240 17688 49292 17740
rect 46664 17663 46716 17672
rect 46664 17629 46673 17663
rect 46673 17629 46707 17663
rect 46707 17629 46716 17663
rect 46664 17620 46716 17629
rect 46756 17620 46808 17672
rect 46940 17620 46992 17672
rect 50160 17620 50212 17672
rect 41604 17552 41656 17604
rect 46388 17552 46440 17604
rect 50712 17620 50764 17672
rect 39580 17484 39632 17536
rect 43168 17484 43220 17536
rect 48412 17527 48464 17536
rect 48412 17493 48421 17527
rect 48421 17493 48455 17527
rect 48455 17493 48464 17527
rect 48412 17484 48464 17493
rect 48780 17527 48832 17536
rect 48780 17493 48789 17527
rect 48789 17493 48823 17527
rect 48823 17493 48832 17527
rect 48780 17484 48832 17493
rect 48872 17527 48924 17536
rect 48872 17493 48881 17527
rect 48881 17493 48915 17527
rect 48915 17493 48924 17527
rect 48872 17484 48924 17493
rect 50068 17484 50120 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 26608 17144 26660 17196
rect 27528 17076 27580 17128
rect 29184 17212 29236 17264
rect 31760 17280 31812 17332
rect 33600 17323 33652 17332
rect 33600 17289 33609 17323
rect 33609 17289 33643 17323
rect 33643 17289 33652 17323
rect 33600 17280 33652 17289
rect 34704 17280 34756 17332
rect 36360 17280 36412 17332
rect 38752 17280 38804 17332
rect 38844 17280 38896 17332
rect 28908 17076 28960 17128
rect 31576 17187 31628 17196
rect 31576 17153 31585 17187
rect 31585 17153 31619 17187
rect 31619 17153 31628 17187
rect 31576 17144 31628 17153
rect 32036 17144 32088 17196
rect 33232 17144 33284 17196
rect 35348 17212 35400 17264
rect 37832 17212 37884 17264
rect 33968 17187 34020 17196
rect 33968 17153 34002 17187
rect 34002 17153 34020 17187
rect 33968 17144 34020 17153
rect 31760 17076 31812 17128
rect 31852 17119 31904 17128
rect 31852 17085 31861 17119
rect 31861 17085 31895 17119
rect 31895 17085 31904 17119
rect 35900 17187 35952 17196
rect 35900 17153 35909 17187
rect 35909 17153 35943 17187
rect 35943 17153 35952 17187
rect 35900 17144 35952 17153
rect 36176 17144 36228 17196
rect 36452 17144 36504 17196
rect 39488 17280 39540 17332
rect 41604 17323 41656 17332
rect 41604 17289 41613 17323
rect 41613 17289 41647 17323
rect 41647 17289 41656 17323
rect 41604 17280 41656 17289
rect 44364 17280 44416 17332
rect 46480 17280 46532 17332
rect 47032 17280 47084 17332
rect 39948 17212 40000 17264
rect 39580 17144 39632 17196
rect 43904 17144 43956 17196
rect 45652 17144 45704 17196
rect 46388 17187 46440 17196
rect 46388 17153 46397 17187
rect 46397 17153 46431 17187
rect 46431 17153 46440 17187
rect 46388 17144 46440 17153
rect 50068 17187 50120 17196
rect 31852 17076 31904 17085
rect 32128 17008 32180 17060
rect 38936 17076 38988 17128
rect 40960 17119 41012 17128
rect 40960 17085 40969 17119
rect 40969 17085 41003 17119
rect 41003 17085 41012 17119
rect 40960 17076 41012 17085
rect 42800 17119 42852 17128
rect 42800 17085 42809 17119
rect 42809 17085 42843 17119
rect 42843 17085 42852 17119
rect 42800 17076 42852 17085
rect 25780 16940 25832 16992
rect 28816 16940 28868 16992
rect 30288 16983 30340 16992
rect 30288 16949 30297 16983
rect 30297 16949 30331 16983
rect 30331 16949 30340 16983
rect 30288 16940 30340 16949
rect 30380 16940 30432 16992
rect 35624 16940 35676 16992
rect 41236 17008 41288 17060
rect 40868 16983 40920 16992
rect 40868 16949 40877 16983
rect 40877 16949 40911 16983
rect 40911 16949 40920 16983
rect 47308 17076 47360 17128
rect 48228 17119 48280 17128
rect 48228 17085 48237 17119
rect 48237 17085 48271 17119
rect 48271 17085 48280 17119
rect 48228 17076 48280 17085
rect 48504 17119 48556 17128
rect 48504 17085 48513 17119
rect 48513 17085 48547 17119
rect 48547 17085 48556 17119
rect 48504 17076 48556 17085
rect 50068 17153 50077 17187
rect 50077 17153 50111 17187
rect 50111 17153 50120 17187
rect 50068 17144 50120 17153
rect 46572 17051 46624 17060
rect 46572 17017 46581 17051
rect 46581 17017 46615 17051
rect 46615 17017 46624 17051
rect 46572 17008 46624 17017
rect 49792 17008 49844 17060
rect 68468 17051 68520 17060
rect 68468 17017 68477 17051
rect 68477 17017 68511 17051
rect 68511 17017 68520 17051
rect 68468 17008 68520 17017
rect 40868 16940 40920 16949
rect 44916 16983 44968 16992
rect 44916 16949 44925 16983
rect 44925 16949 44959 16983
rect 44959 16949 44968 16983
rect 44916 16940 44968 16949
rect 45928 16940 45980 16992
rect 46204 16983 46256 16992
rect 46204 16949 46213 16983
rect 46213 16949 46247 16983
rect 46247 16949 46256 16983
rect 46204 16940 46256 16949
rect 49240 16940 49292 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 28724 16736 28776 16788
rect 28816 16736 28868 16788
rect 33048 16736 33100 16788
rect 25228 16532 25280 16584
rect 25780 16575 25832 16584
rect 25780 16541 25814 16575
rect 25814 16541 25832 16575
rect 25780 16532 25832 16541
rect 27988 16575 28040 16584
rect 27988 16541 27997 16575
rect 27997 16541 28031 16575
rect 28031 16541 28040 16575
rect 27988 16532 28040 16541
rect 37832 16779 37884 16788
rect 37832 16745 37841 16779
rect 37841 16745 37875 16779
rect 37875 16745 37884 16779
rect 37832 16736 37884 16745
rect 39396 16736 39448 16788
rect 29184 16600 29236 16652
rect 28724 16532 28776 16584
rect 28908 16464 28960 16516
rect 29460 16532 29512 16584
rect 30288 16532 30340 16584
rect 35624 16575 35676 16584
rect 35624 16541 35658 16575
rect 35658 16541 35676 16575
rect 35624 16532 35676 16541
rect 38200 16507 38252 16516
rect 38200 16473 38209 16507
rect 38209 16473 38243 16507
rect 38243 16473 38252 16507
rect 38200 16464 38252 16473
rect 26884 16439 26936 16448
rect 26884 16405 26893 16439
rect 26893 16405 26927 16439
rect 26927 16405 26936 16439
rect 26884 16396 26936 16405
rect 26976 16439 27028 16448
rect 26976 16405 26985 16439
rect 26985 16405 27019 16439
rect 27019 16405 27028 16439
rect 26976 16396 27028 16405
rect 27344 16439 27396 16448
rect 27344 16405 27353 16439
rect 27353 16405 27387 16439
rect 27387 16405 27396 16439
rect 27344 16396 27396 16405
rect 28632 16396 28684 16448
rect 29368 16396 29420 16448
rect 30288 16396 30340 16448
rect 35348 16396 35400 16448
rect 38016 16396 38068 16448
rect 39028 16439 39080 16448
rect 39028 16405 39037 16439
rect 39037 16405 39071 16439
rect 39071 16405 39080 16439
rect 39028 16396 39080 16405
rect 39488 16439 39540 16448
rect 39488 16405 39497 16439
rect 39497 16405 39531 16439
rect 39531 16405 39540 16439
rect 39488 16396 39540 16405
rect 39948 16464 40000 16516
rect 43168 16668 43220 16720
rect 45928 16736 45980 16788
rect 46204 16736 46256 16788
rect 48504 16736 48556 16788
rect 48780 16736 48832 16788
rect 42616 16600 42668 16652
rect 44088 16600 44140 16652
rect 43812 16532 43864 16584
rect 44272 16575 44324 16584
rect 44272 16541 44281 16575
rect 44281 16541 44315 16575
rect 44315 16541 44324 16575
rect 44272 16532 44324 16541
rect 42892 16464 42944 16516
rect 40224 16396 40276 16448
rect 42248 16439 42300 16448
rect 42248 16405 42257 16439
rect 42257 16405 42291 16439
rect 42291 16405 42300 16439
rect 42248 16396 42300 16405
rect 42524 16439 42576 16448
rect 42524 16405 42539 16439
rect 42539 16405 42573 16439
rect 42573 16405 42576 16439
rect 42524 16396 42576 16405
rect 43444 16439 43496 16448
rect 43444 16405 43453 16439
rect 43453 16405 43487 16439
rect 43487 16405 43496 16439
rect 43444 16396 43496 16405
rect 44272 16396 44324 16448
rect 44548 16507 44600 16516
rect 44548 16473 44557 16507
rect 44557 16473 44591 16507
rect 44591 16473 44600 16507
rect 44548 16464 44600 16473
rect 45008 16507 45060 16516
rect 45008 16473 45017 16507
rect 45017 16473 45051 16507
rect 45051 16473 45060 16507
rect 45008 16464 45060 16473
rect 45376 16575 45428 16584
rect 45376 16541 45385 16575
rect 45385 16541 45419 16575
rect 45419 16541 45428 16575
rect 45376 16532 45428 16541
rect 46664 16600 46716 16652
rect 48780 16600 48832 16652
rect 49240 16643 49292 16652
rect 49240 16609 49249 16643
rect 49249 16609 49283 16643
rect 49283 16609 49292 16643
rect 49240 16600 49292 16609
rect 46756 16575 46808 16584
rect 46756 16541 46765 16575
rect 46765 16541 46799 16575
rect 46799 16541 46808 16575
rect 46756 16532 46808 16541
rect 48412 16575 48464 16584
rect 48412 16541 48421 16575
rect 48421 16541 48455 16575
rect 48455 16541 48464 16575
rect 48412 16532 48464 16541
rect 45652 16464 45704 16516
rect 49792 16464 49844 16516
rect 51816 16575 51868 16584
rect 51816 16541 51825 16575
rect 51825 16541 51859 16575
rect 51859 16541 51868 16575
rect 51816 16532 51868 16541
rect 44640 16396 44692 16448
rect 44732 16396 44784 16448
rect 45192 16439 45244 16448
rect 45192 16405 45201 16439
rect 45201 16405 45235 16439
rect 45235 16405 45244 16439
rect 45192 16396 45244 16405
rect 49700 16396 49752 16448
rect 51448 16396 51500 16448
rect 52368 16439 52420 16448
rect 52368 16405 52377 16439
rect 52377 16405 52411 16439
rect 52411 16405 52420 16439
rect 52368 16396 52420 16405
rect 52736 16396 52788 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 26148 16124 26200 16176
rect 26056 16099 26108 16108
rect 26056 16065 26065 16099
rect 26065 16065 26099 16099
rect 26099 16065 26108 16099
rect 26056 16056 26108 16065
rect 26148 15988 26200 16040
rect 26608 16235 26660 16244
rect 26608 16201 26617 16235
rect 26617 16201 26651 16235
rect 26651 16201 26660 16235
rect 26608 16192 26660 16201
rect 26700 16192 26752 16244
rect 26976 16192 27028 16244
rect 27344 16192 27396 16244
rect 27988 16192 28040 16244
rect 28908 16192 28960 16244
rect 29368 16192 29420 16244
rect 28816 16056 28868 16108
rect 29276 16099 29328 16108
rect 29276 16065 29285 16099
rect 29285 16065 29319 16099
rect 29319 16065 29328 16099
rect 29276 16056 29328 16065
rect 30012 16192 30064 16244
rect 31760 16192 31812 16244
rect 39948 16192 40000 16244
rect 40868 16235 40920 16244
rect 40868 16201 40877 16235
rect 40877 16201 40911 16235
rect 40911 16201 40920 16235
rect 40868 16192 40920 16201
rect 31484 16124 31536 16176
rect 27528 16031 27580 16040
rect 27528 15997 27537 16031
rect 27537 15997 27571 16031
rect 27571 15997 27580 16031
rect 27528 15988 27580 15997
rect 29000 15988 29052 16040
rect 29368 15988 29420 16040
rect 30656 16056 30708 16108
rect 29920 15988 29972 16040
rect 30288 15988 30340 16040
rect 31116 16056 31168 16108
rect 31208 16031 31260 16040
rect 31208 15997 31217 16031
rect 31217 15997 31251 16031
rect 31251 15997 31260 16031
rect 31208 15988 31260 15997
rect 25228 15920 25280 15972
rect 28540 15920 28592 15972
rect 33048 16056 33100 16108
rect 32128 16031 32180 16040
rect 32128 15997 32137 16031
rect 32137 15997 32171 16031
rect 32171 15997 32180 16031
rect 32128 15988 32180 15997
rect 33416 16099 33468 16108
rect 33416 16065 33425 16099
rect 33425 16065 33459 16099
rect 33459 16065 33468 16099
rect 33416 16056 33468 16065
rect 37832 16124 37884 16176
rect 38108 16124 38160 16176
rect 34520 16056 34572 16108
rect 37096 16056 37148 16108
rect 39396 16099 39448 16108
rect 39396 16065 39430 16099
rect 39430 16065 39448 16099
rect 39396 16056 39448 16065
rect 42248 16192 42300 16244
rect 42524 16192 42576 16244
rect 33784 16031 33836 16040
rect 33784 15997 33793 16031
rect 33793 15997 33827 16031
rect 33827 15997 33836 16031
rect 33784 15988 33836 15997
rect 37280 16031 37332 16040
rect 37280 15997 37289 16031
rect 37289 15997 37323 16031
rect 37323 15997 37332 16031
rect 37280 15988 37332 15997
rect 40224 16056 40276 16108
rect 41052 16056 41104 16108
rect 42800 16124 42852 16176
rect 43444 16124 43496 16176
rect 43904 16192 43956 16244
rect 44088 16192 44140 16244
rect 44640 16192 44692 16244
rect 44916 16192 44968 16244
rect 34612 15920 34664 15972
rect 40960 15920 41012 15972
rect 44732 16167 44784 16176
rect 44732 16133 44741 16167
rect 44741 16133 44775 16167
rect 44775 16133 44784 16167
rect 44732 16124 44784 16133
rect 45744 16124 45796 16176
rect 44088 16099 44140 16108
rect 44088 16065 44097 16099
rect 44097 16065 44131 16099
rect 44131 16065 44140 16099
rect 44088 16056 44140 16065
rect 44456 16031 44508 16040
rect 44456 15997 44465 16031
rect 44465 15997 44499 16031
rect 44499 15997 44508 16031
rect 44456 15988 44508 15997
rect 51816 16192 51868 16244
rect 51448 16124 51500 16176
rect 46480 16099 46532 16108
rect 46480 16065 46489 16099
rect 46489 16065 46523 16099
rect 46523 16065 46532 16099
rect 46480 16056 46532 16065
rect 46572 16056 46624 16108
rect 48504 16056 48556 16108
rect 940 15852 992 15904
rect 24860 15852 24912 15904
rect 28724 15852 28776 15904
rect 31852 15895 31904 15904
rect 31852 15861 31861 15895
rect 31861 15861 31895 15895
rect 31895 15861 31904 15895
rect 31852 15852 31904 15861
rect 33140 15895 33192 15904
rect 33140 15861 33149 15895
rect 33149 15861 33183 15895
rect 33183 15861 33192 15895
rect 33140 15852 33192 15861
rect 38660 15852 38712 15904
rect 39488 15852 39540 15904
rect 43812 15895 43864 15904
rect 43812 15861 43821 15895
rect 43821 15861 43855 15895
rect 43855 15861 43864 15895
rect 43812 15852 43864 15861
rect 45744 15852 45796 15904
rect 46296 15895 46348 15904
rect 46296 15861 46305 15895
rect 46305 15861 46339 15895
rect 46339 15861 46348 15895
rect 46296 15852 46348 15861
rect 48228 15852 48280 15904
rect 48964 15852 49016 15904
rect 50436 16031 50488 16040
rect 50436 15997 50445 16031
rect 50445 15997 50479 16031
rect 50479 15997 50488 16031
rect 50436 15988 50488 15997
rect 52276 15852 52328 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 26056 15648 26108 15700
rect 27344 15648 27396 15700
rect 28540 15648 28592 15700
rect 28816 15648 28868 15700
rect 31116 15648 31168 15700
rect 32956 15648 33008 15700
rect 37464 15648 37516 15700
rect 38108 15691 38160 15700
rect 38108 15657 38117 15691
rect 38117 15657 38151 15691
rect 38151 15657 38160 15691
rect 38108 15648 38160 15657
rect 38660 15648 38712 15700
rect 39396 15648 39448 15700
rect 42892 15691 42944 15700
rect 42892 15657 42901 15691
rect 42901 15657 42935 15691
rect 42935 15657 42944 15691
rect 42892 15648 42944 15657
rect 26240 15512 26292 15564
rect 27252 15512 27304 15564
rect 29368 15580 29420 15632
rect 30196 15580 30248 15632
rect 28632 15555 28684 15564
rect 28632 15521 28641 15555
rect 28641 15521 28675 15555
rect 28675 15521 28684 15555
rect 28632 15512 28684 15521
rect 28724 15512 28776 15564
rect 25136 15487 25188 15496
rect 25136 15453 25145 15487
rect 25145 15453 25179 15487
rect 25179 15453 25188 15487
rect 25136 15444 25188 15453
rect 26056 15487 26108 15496
rect 26056 15453 26065 15487
rect 26065 15453 26099 15487
rect 26099 15453 26108 15487
rect 26056 15444 26108 15453
rect 26884 15444 26936 15496
rect 27620 15444 27672 15496
rect 28080 15444 28132 15496
rect 26976 15376 27028 15428
rect 29644 15512 29696 15564
rect 29092 15444 29144 15496
rect 30104 15444 30156 15496
rect 30748 15487 30800 15496
rect 30748 15453 30757 15487
rect 30757 15453 30791 15487
rect 30791 15453 30800 15487
rect 30748 15444 30800 15453
rect 32312 15444 32364 15496
rect 35348 15444 35400 15496
rect 37280 15444 37332 15496
rect 40132 15580 40184 15632
rect 44916 15648 44968 15700
rect 45376 15648 45428 15700
rect 46296 15648 46348 15700
rect 46756 15648 46808 15700
rect 48228 15648 48280 15700
rect 50436 15648 50488 15700
rect 39304 15512 39356 15564
rect 39948 15512 40000 15564
rect 38016 15487 38068 15496
rect 31668 15376 31720 15428
rect 33140 15376 33192 15428
rect 26240 15308 26292 15360
rect 26608 15351 26660 15360
rect 26608 15317 26617 15351
rect 26617 15317 26651 15351
rect 26651 15317 26660 15351
rect 26608 15308 26660 15317
rect 27068 15308 27120 15360
rect 28724 15308 28776 15360
rect 29552 15351 29604 15360
rect 29552 15317 29561 15351
rect 29561 15317 29595 15351
rect 29595 15317 29604 15351
rect 29552 15308 29604 15317
rect 30656 15308 30708 15360
rect 34796 15376 34848 15428
rect 37556 15376 37608 15428
rect 38016 15453 38025 15487
rect 38025 15453 38059 15487
rect 38059 15453 38068 15487
rect 38016 15444 38068 15453
rect 38844 15487 38896 15496
rect 38844 15453 38853 15487
rect 38853 15453 38887 15487
rect 38887 15453 38896 15487
rect 38844 15444 38896 15453
rect 39028 15444 39080 15496
rect 40224 15444 40276 15496
rect 40408 15487 40460 15496
rect 40408 15453 40417 15487
rect 40417 15453 40451 15487
rect 40451 15453 40460 15487
rect 40408 15444 40460 15453
rect 42800 15512 42852 15564
rect 43628 15512 43680 15564
rect 44732 15512 44784 15564
rect 52000 15648 52052 15700
rect 52368 15648 52420 15700
rect 52552 15580 52604 15632
rect 44640 15444 44692 15496
rect 47400 15444 47452 15496
rect 39212 15419 39264 15428
rect 39212 15385 39221 15419
rect 39221 15385 39255 15419
rect 39255 15385 39264 15419
rect 39212 15376 39264 15385
rect 44364 15376 44416 15428
rect 33968 15351 34020 15360
rect 33968 15317 33977 15351
rect 33977 15317 34011 15351
rect 34011 15317 34020 15351
rect 33968 15308 34020 15317
rect 34704 15308 34756 15360
rect 36084 15351 36136 15360
rect 36084 15317 36093 15351
rect 36093 15317 36127 15351
rect 36127 15317 36136 15351
rect 36084 15308 36136 15317
rect 44180 15308 44232 15360
rect 45836 15308 45888 15360
rect 49792 15487 49844 15496
rect 49792 15453 49801 15487
rect 49801 15453 49835 15487
rect 49835 15453 49844 15487
rect 49792 15444 49844 15453
rect 51816 15487 51868 15496
rect 51816 15453 51825 15487
rect 51825 15453 51859 15487
rect 51859 15453 51868 15487
rect 51816 15444 51868 15453
rect 52644 15487 52696 15496
rect 52644 15453 52653 15487
rect 52653 15453 52687 15487
rect 52687 15453 52696 15487
rect 52644 15444 52696 15453
rect 51632 15376 51684 15428
rect 52092 15376 52144 15428
rect 52184 15419 52236 15428
rect 52184 15385 52193 15419
rect 52193 15385 52227 15419
rect 52227 15385 52236 15419
rect 52184 15376 52236 15385
rect 48504 15308 48556 15360
rect 49884 15351 49936 15360
rect 49884 15317 49893 15351
rect 49893 15317 49927 15351
rect 49927 15317 49936 15351
rect 49884 15308 49936 15317
rect 52000 15308 52052 15360
rect 52460 15308 52512 15360
rect 54484 15444 54536 15496
rect 53932 15351 53984 15360
rect 53932 15317 53941 15351
rect 53941 15317 53975 15351
rect 53975 15317 53984 15351
rect 53932 15308 53984 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 26056 15104 26108 15156
rect 24860 14968 24912 15020
rect 27620 15104 27672 15156
rect 27068 14968 27120 15020
rect 27252 14968 27304 15020
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 28080 15011 28132 15020
rect 28080 14977 28089 15011
rect 28089 14977 28123 15011
rect 28123 14977 28132 15011
rect 28080 14968 28132 14977
rect 25228 14943 25280 14952
rect 25228 14909 25237 14943
rect 25237 14909 25271 14943
rect 25271 14909 25280 14943
rect 25228 14900 25280 14909
rect 28908 15104 28960 15156
rect 29092 15147 29144 15156
rect 29092 15113 29101 15147
rect 29101 15113 29135 15147
rect 29135 15113 29144 15147
rect 29092 15104 29144 15113
rect 31208 15104 31260 15156
rect 31668 15147 31720 15156
rect 31668 15113 31677 15147
rect 31677 15113 31711 15147
rect 31711 15113 31720 15147
rect 31668 15104 31720 15113
rect 31852 15104 31904 15156
rect 33784 15104 33836 15156
rect 34428 15147 34480 15156
rect 34428 15113 34437 15147
rect 34437 15113 34471 15147
rect 34471 15113 34480 15147
rect 34428 15104 34480 15113
rect 28724 15011 28776 15020
rect 28724 14977 28733 15011
rect 28733 14977 28767 15011
rect 28767 14977 28776 15011
rect 28724 14968 28776 14977
rect 29552 15036 29604 15088
rect 29460 15011 29512 15020
rect 29460 14977 29469 15011
rect 29469 14977 29503 15011
rect 29503 14977 29512 15011
rect 29460 14968 29512 14977
rect 30748 14968 30800 15020
rect 38660 15104 38712 15156
rect 40408 15104 40460 15156
rect 33140 14968 33192 15020
rect 33416 14968 33468 15020
rect 34704 15036 34756 15088
rect 34520 14968 34572 15020
rect 38844 15036 38896 15088
rect 42616 15104 42668 15156
rect 44364 15104 44416 15156
rect 45192 15104 45244 15156
rect 48964 15104 49016 15156
rect 35348 15011 35400 15020
rect 35348 14977 35364 15011
rect 35364 14977 35398 15011
rect 35398 14977 35400 15011
rect 35348 14968 35400 14977
rect 36452 14968 36504 15020
rect 31024 14943 31076 14952
rect 31024 14909 31033 14943
rect 31033 14909 31067 14943
rect 31067 14909 31076 14943
rect 31024 14900 31076 14909
rect 32312 14943 32364 14952
rect 32312 14909 32321 14943
rect 32321 14909 32355 14943
rect 32355 14909 32364 14943
rect 32312 14900 32364 14909
rect 34244 14900 34296 14952
rect 39488 15011 39540 15020
rect 39488 14977 39497 15011
rect 39497 14977 39531 15011
rect 39531 14977 39540 15011
rect 39488 14968 39540 14977
rect 39212 14900 39264 14952
rect 40408 15011 40460 15020
rect 40408 14977 40417 15011
rect 40417 14977 40451 15011
rect 40451 14977 40460 15011
rect 40408 14968 40460 14977
rect 40500 15011 40552 15020
rect 40500 14977 40509 15011
rect 40509 14977 40543 15011
rect 40543 14977 40552 15011
rect 40500 14968 40552 14977
rect 40776 14968 40828 15020
rect 43812 15036 43864 15088
rect 42800 14968 42852 15020
rect 42892 15011 42944 15020
rect 42892 14977 42901 15011
rect 42901 14977 42935 15011
rect 42935 14977 42944 15011
rect 42892 14968 42944 14977
rect 42248 14900 42300 14952
rect 43812 14943 43864 14952
rect 43812 14909 43821 14943
rect 43821 14909 43855 14943
rect 43855 14909 43864 14943
rect 43812 14900 43864 14909
rect 44088 14900 44140 14952
rect 44272 14900 44324 14952
rect 25136 14807 25188 14816
rect 25136 14773 25145 14807
rect 25145 14773 25179 14807
rect 25179 14773 25188 14807
rect 25136 14764 25188 14773
rect 27896 14807 27948 14816
rect 27896 14773 27905 14807
rect 27905 14773 27939 14807
rect 27939 14773 27948 14807
rect 27896 14764 27948 14773
rect 29276 14807 29328 14816
rect 29276 14773 29285 14807
rect 29285 14773 29319 14807
rect 29319 14773 29328 14807
rect 29276 14764 29328 14773
rect 33600 14764 33652 14816
rect 33692 14764 33744 14816
rect 35256 14764 35308 14816
rect 36360 14764 36412 14816
rect 36544 14764 36596 14816
rect 36728 14807 36780 14816
rect 36728 14773 36737 14807
rect 36737 14773 36771 14807
rect 36771 14773 36780 14807
rect 36728 14764 36780 14773
rect 36820 14807 36872 14816
rect 36820 14773 36829 14807
rect 36829 14773 36863 14807
rect 36863 14773 36872 14807
rect 36820 14764 36872 14773
rect 38936 14764 38988 14816
rect 39580 14807 39632 14816
rect 39580 14773 39589 14807
rect 39589 14773 39623 14807
rect 39623 14773 39632 14807
rect 39580 14764 39632 14773
rect 40132 14807 40184 14816
rect 40132 14773 40141 14807
rect 40141 14773 40175 14807
rect 40175 14773 40184 14807
rect 40132 14764 40184 14773
rect 40684 14764 40736 14816
rect 40960 14764 41012 14816
rect 44180 14764 44232 14816
rect 44732 14968 44784 15020
rect 45652 14968 45704 15020
rect 46572 14968 46624 15020
rect 46756 14968 46808 15020
rect 48780 15036 48832 15088
rect 51724 15104 51776 15156
rect 49884 15036 49936 15088
rect 51264 15079 51316 15088
rect 51264 15045 51273 15079
rect 51273 15045 51307 15079
rect 51307 15045 51316 15079
rect 51264 15036 51316 15045
rect 51632 15036 51684 15088
rect 53932 15104 53984 15156
rect 54484 15147 54536 15156
rect 54484 15113 54493 15147
rect 54493 15113 54527 15147
rect 54527 15113 54536 15147
rect 54484 15104 54536 15113
rect 52276 15036 52328 15088
rect 47584 14943 47636 14952
rect 47584 14909 47593 14943
rect 47593 14909 47627 14943
rect 47627 14909 47636 14943
rect 47584 14900 47636 14909
rect 48596 14900 48648 14952
rect 48688 14943 48740 14952
rect 48688 14909 48697 14943
rect 48697 14909 48731 14943
rect 48731 14909 48740 14943
rect 48688 14900 48740 14909
rect 49148 14943 49200 14952
rect 49148 14909 49157 14943
rect 49157 14909 49191 14943
rect 49191 14909 49200 14943
rect 49148 14900 49200 14909
rect 51448 14900 51500 14952
rect 52092 15011 52144 15020
rect 52092 14977 52101 15011
rect 52101 14977 52135 15011
rect 52135 14977 52144 15011
rect 52092 14968 52144 14977
rect 52460 14968 52512 15020
rect 52552 15011 52604 15020
rect 52552 14977 52561 15011
rect 52561 14977 52595 15011
rect 52595 14977 52604 15011
rect 52552 14968 52604 14977
rect 53472 15036 53524 15088
rect 47492 14764 47544 14816
rect 48320 14764 48372 14816
rect 48688 14764 48740 14816
rect 49792 14764 49844 14816
rect 50712 14764 50764 14816
rect 51540 14764 51592 14816
rect 52000 14764 52052 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 26332 14603 26384 14612
rect 26332 14569 26341 14603
rect 26341 14569 26375 14603
rect 26375 14569 26384 14603
rect 26332 14560 26384 14569
rect 26884 14603 26936 14612
rect 26884 14569 26893 14603
rect 26893 14569 26927 14603
rect 26927 14569 26936 14603
rect 26884 14560 26936 14569
rect 29276 14560 29328 14612
rect 31024 14603 31076 14612
rect 31024 14569 31033 14603
rect 31033 14569 31067 14603
rect 31067 14569 31076 14603
rect 31024 14560 31076 14569
rect 24860 14424 24912 14476
rect 26056 14424 26108 14476
rect 25136 14356 25188 14408
rect 29920 14535 29972 14544
rect 29920 14501 29929 14535
rect 29929 14501 29963 14535
rect 29963 14501 29972 14535
rect 29920 14492 29972 14501
rect 26240 14399 26292 14408
rect 26240 14365 26249 14399
rect 26249 14365 26283 14399
rect 26283 14365 26292 14399
rect 26240 14356 26292 14365
rect 26608 14356 26660 14408
rect 26976 14356 27028 14408
rect 27068 14356 27120 14408
rect 27344 14356 27396 14408
rect 29644 14356 29696 14408
rect 30748 14424 30800 14476
rect 25964 14220 26016 14272
rect 28632 14263 28684 14272
rect 28632 14229 28641 14263
rect 28641 14229 28675 14263
rect 28675 14229 28684 14263
rect 31116 14356 31168 14408
rect 31484 14399 31536 14408
rect 31484 14365 31493 14399
rect 31493 14365 31527 14399
rect 31527 14365 31536 14399
rect 31484 14356 31536 14365
rect 31852 14560 31904 14612
rect 33140 14603 33192 14612
rect 33140 14569 33149 14603
rect 33149 14569 33183 14603
rect 33183 14569 33192 14603
rect 33140 14560 33192 14569
rect 33600 14560 33652 14612
rect 34428 14560 34480 14612
rect 34612 14560 34664 14612
rect 34796 14560 34848 14612
rect 36452 14603 36504 14612
rect 36452 14569 36461 14603
rect 36461 14569 36495 14603
rect 36495 14569 36504 14603
rect 36452 14560 36504 14569
rect 37096 14560 37148 14612
rect 31944 14399 31996 14408
rect 31944 14365 31953 14399
rect 31953 14365 31987 14399
rect 31987 14365 31996 14399
rect 31944 14356 31996 14365
rect 32956 14356 33008 14408
rect 33324 14399 33376 14408
rect 33324 14365 33333 14399
rect 33333 14365 33367 14399
rect 33367 14365 33376 14399
rect 33324 14356 33376 14365
rect 28632 14220 28684 14229
rect 32496 14263 32548 14272
rect 32496 14229 32505 14263
rect 32505 14229 32539 14263
rect 32539 14229 32548 14263
rect 32496 14220 32548 14229
rect 32680 14288 32732 14340
rect 33968 14467 34020 14476
rect 33968 14433 33977 14467
rect 33977 14433 34011 14467
rect 34011 14433 34020 14467
rect 33968 14424 34020 14433
rect 34520 14356 34572 14408
rect 34704 14356 34756 14408
rect 35348 14399 35400 14408
rect 35348 14365 35357 14399
rect 35357 14365 35391 14399
rect 35391 14365 35400 14399
rect 35348 14356 35400 14365
rect 36360 14424 36412 14476
rect 36728 14467 36780 14476
rect 36728 14433 36737 14467
rect 36737 14433 36771 14467
rect 36771 14433 36780 14467
rect 36728 14424 36780 14433
rect 32772 14220 32824 14272
rect 35072 14331 35124 14340
rect 35072 14297 35081 14331
rect 35081 14297 35115 14331
rect 35115 14297 35124 14331
rect 35072 14288 35124 14297
rect 37004 14356 37056 14408
rect 37464 14331 37516 14340
rect 37464 14297 37473 14331
rect 37473 14297 37507 14331
rect 37507 14297 37516 14331
rect 37464 14288 37516 14297
rect 39488 14492 39540 14544
rect 39764 14560 39816 14612
rect 40500 14560 40552 14612
rect 40684 14560 40736 14612
rect 42248 14560 42300 14612
rect 42892 14603 42944 14612
rect 42892 14569 42901 14603
rect 42901 14569 42935 14603
rect 42935 14569 42944 14603
rect 42892 14560 42944 14569
rect 46572 14560 46624 14612
rect 47216 14560 47268 14612
rect 47492 14560 47544 14612
rect 47584 14560 47636 14612
rect 48964 14560 49016 14612
rect 49148 14560 49200 14612
rect 49700 14560 49752 14612
rect 51264 14560 51316 14612
rect 52000 14560 52052 14612
rect 52644 14560 52696 14612
rect 53472 14560 53524 14612
rect 42708 14492 42760 14544
rect 42800 14492 42852 14544
rect 40224 14424 40276 14476
rect 39672 14356 39724 14408
rect 42524 14399 42576 14408
rect 40316 14288 40368 14340
rect 42524 14365 42530 14399
rect 42530 14365 42564 14399
rect 42564 14365 42576 14399
rect 42524 14356 42576 14365
rect 47308 14535 47360 14544
rect 47308 14501 47317 14535
rect 47317 14501 47351 14535
rect 47351 14501 47360 14535
rect 47308 14492 47360 14501
rect 47400 14535 47452 14544
rect 47400 14501 47409 14535
rect 47409 14501 47443 14535
rect 47443 14501 47452 14535
rect 47400 14492 47452 14501
rect 43076 14399 43128 14408
rect 43076 14365 43085 14399
rect 43085 14365 43119 14399
rect 43119 14365 43128 14399
rect 43076 14356 43128 14365
rect 45560 14424 45612 14476
rect 46480 14424 46532 14476
rect 46756 14424 46808 14476
rect 43812 14356 43864 14408
rect 44088 14356 44140 14408
rect 48688 14492 48740 14544
rect 48872 14492 48924 14544
rect 48872 14356 48924 14408
rect 36728 14220 36780 14272
rect 38568 14220 38620 14272
rect 40500 14263 40552 14272
rect 40500 14229 40509 14263
rect 40509 14229 40543 14263
rect 40543 14229 40552 14263
rect 40500 14220 40552 14229
rect 41236 14263 41288 14272
rect 41236 14229 41245 14263
rect 41245 14229 41279 14263
rect 41279 14229 41288 14263
rect 41236 14220 41288 14229
rect 42248 14220 42300 14272
rect 43168 14263 43220 14272
rect 43168 14229 43177 14263
rect 43177 14229 43211 14263
rect 43211 14229 43220 14263
rect 43168 14220 43220 14229
rect 45836 14220 45888 14272
rect 48688 14288 48740 14340
rect 49700 14399 49752 14408
rect 49700 14365 49709 14399
rect 49709 14365 49743 14399
rect 49743 14365 49752 14399
rect 49700 14356 49752 14365
rect 49792 14356 49844 14408
rect 50988 14399 51040 14408
rect 50988 14365 50997 14399
rect 50997 14365 51031 14399
rect 51031 14365 51040 14399
rect 50988 14356 51040 14365
rect 51448 14356 51500 14408
rect 50160 14288 50212 14340
rect 50620 14331 50672 14340
rect 50620 14297 50629 14331
rect 50629 14297 50663 14331
rect 50663 14297 50672 14331
rect 50620 14288 50672 14297
rect 50804 14288 50856 14340
rect 52460 14356 52512 14408
rect 52552 14356 52604 14408
rect 52736 14399 52788 14408
rect 52736 14365 52745 14399
rect 52745 14365 52779 14399
rect 52779 14365 52788 14399
rect 52736 14356 52788 14365
rect 68468 14399 68520 14408
rect 68468 14365 68477 14399
rect 68477 14365 68511 14399
rect 68511 14365 68520 14399
rect 68468 14356 68520 14365
rect 48228 14263 48280 14272
rect 48228 14229 48237 14263
rect 48237 14229 48271 14263
rect 48271 14229 48280 14263
rect 48228 14220 48280 14229
rect 48596 14263 48648 14272
rect 48596 14229 48605 14263
rect 48605 14229 48639 14263
rect 48639 14229 48648 14263
rect 53472 14288 53524 14340
rect 48596 14220 48648 14229
rect 51264 14263 51316 14272
rect 51264 14229 51273 14263
rect 51273 14229 51307 14263
rect 51307 14229 51316 14263
rect 51264 14220 51316 14229
rect 51632 14263 51684 14272
rect 51632 14229 51641 14263
rect 51641 14229 51675 14263
rect 51675 14229 51684 14263
rect 51632 14220 51684 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 27896 14016 27948 14068
rect 28632 14016 28684 14068
rect 31944 14016 31996 14068
rect 23940 13948 23992 14000
rect 29736 13923 29788 13932
rect 29736 13889 29770 13923
rect 29770 13889 29788 13923
rect 22376 13812 22428 13864
rect 23204 13855 23256 13864
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 24860 13812 24912 13864
rect 29736 13880 29788 13889
rect 33048 13948 33100 14000
rect 32220 13880 32272 13932
rect 34612 14016 34664 14068
rect 35348 14016 35400 14068
rect 33784 13923 33836 13932
rect 33784 13889 33793 13923
rect 33793 13889 33827 13923
rect 33827 13889 33836 13923
rect 33784 13880 33836 13889
rect 33968 13880 34020 13932
rect 28172 13855 28224 13864
rect 28172 13821 28181 13855
rect 28181 13821 28215 13855
rect 28215 13821 28224 13855
rect 28172 13812 28224 13821
rect 28356 13812 28408 13864
rect 29000 13812 29052 13864
rect 33232 13812 33284 13864
rect 34244 13923 34296 13932
rect 34244 13889 34253 13923
rect 34253 13889 34287 13923
rect 34287 13889 34296 13923
rect 34244 13880 34296 13889
rect 34152 13812 34204 13864
rect 36084 13880 36136 13932
rect 39028 14016 39080 14068
rect 39764 14016 39816 14068
rect 40224 14059 40276 14068
rect 40224 14025 40233 14059
rect 40233 14025 40267 14059
rect 40267 14025 40276 14059
rect 40224 14016 40276 14025
rect 40500 14016 40552 14068
rect 42248 14059 42300 14068
rect 42248 14025 42257 14059
rect 42257 14025 42291 14059
rect 42291 14025 42300 14059
rect 42248 14016 42300 14025
rect 43168 14016 43220 14068
rect 44732 14059 44784 14068
rect 44732 14025 44741 14059
rect 44741 14025 44775 14059
rect 44775 14025 44784 14059
rect 44732 14016 44784 14025
rect 45652 14016 45704 14068
rect 36820 13948 36872 14000
rect 36912 13948 36964 14000
rect 36728 13923 36780 13932
rect 36728 13889 36737 13923
rect 36737 13889 36771 13923
rect 36771 13889 36780 13923
rect 36728 13880 36780 13889
rect 36544 13812 36596 13864
rect 37280 13923 37332 13932
rect 37280 13889 37289 13923
rect 37289 13889 37323 13923
rect 37323 13889 37332 13923
rect 37280 13880 37332 13889
rect 38660 13880 38712 13932
rect 27804 13719 27856 13728
rect 27804 13685 27813 13719
rect 27813 13685 27847 13719
rect 27847 13685 27856 13719
rect 27804 13676 27856 13685
rect 30104 13676 30156 13728
rect 31116 13676 31168 13728
rect 31668 13676 31720 13728
rect 34336 13744 34388 13796
rect 33876 13719 33928 13728
rect 33876 13685 33885 13719
rect 33885 13685 33919 13719
rect 33919 13685 33928 13719
rect 33876 13676 33928 13685
rect 38844 13855 38896 13864
rect 38844 13821 38853 13855
rect 38853 13821 38887 13855
rect 38887 13821 38896 13855
rect 38844 13812 38896 13821
rect 39856 13812 39908 13864
rect 40960 13880 41012 13932
rect 36912 13787 36964 13796
rect 36912 13753 36921 13787
rect 36921 13753 36955 13787
rect 36955 13753 36964 13787
rect 36912 13744 36964 13753
rect 38752 13676 38804 13728
rect 40776 13676 40828 13728
rect 44824 13855 44876 13864
rect 44824 13821 44833 13855
rect 44833 13821 44867 13855
rect 44867 13821 44876 13855
rect 44824 13812 44876 13821
rect 47216 13880 47268 13932
rect 49608 14016 49660 14068
rect 49700 14016 49752 14068
rect 50804 14016 50856 14068
rect 49792 13948 49844 14000
rect 48412 13880 48464 13932
rect 43812 13787 43864 13796
rect 43812 13753 43821 13787
rect 43821 13753 43855 13787
rect 43855 13753 43864 13787
rect 43812 13744 43864 13753
rect 44548 13744 44600 13796
rect 48136 13855 48188 13864
rect 48136 13821 48145 13855
rect 48145 13821 48179 13855
rect 48179 13821 48188 13855
rect 48136 13812 48188 13821
rect 48688 13880 48740 13932
rect 48872 13880 48924 13932
rect 49148 13880 49200 13932
rect 49240 13923 49292 13932
rect 49240 13889 49249 13923
rect 49249 13889 49283 13923
rect 49283 13889 49292 13923
rect 49240 13880 49292 13889
rect 51264 13948 51316 14000
rect 42800 13676 42852 13728
rect 44364 13719 44416 13728
rect 44364 13685 44373 13719
rect 44373 13685 44407 13719
rect 44407 13685 44416 13719
rect 44364 13676 44416 13685
rect 45192 13719 45244 13728
rect 45192 13685 45201 13719
rect 45201 13685 45235 13719
rect 45235 13685 45244 13719
rect 45192 13676 45244 13685
rect 46388 13719 46440 13728
rect 46388 13685 46397 13719
rect 46397 13685 46431 13719
rect 46431 13685 46440 13719
rect 46388 13676 46440 13685
rect 46480 13719 46532 13728
rect 46480 13685 46489 13719
rect 46489 13685 46523 13719
rect 46523 13685 46532 13719
rect 46480 13676 46532 13685
rect 47032 13676 47084 13728
rect 47952 13676 48004 13728
rect 49424 13812 49476 13864
rect 50252 13880 50304 13932
rect 50712 13812 50764 13864
rect 50160 13744 50212 13796
rect 51172 13855 51224 13864
rect 51172 13821 51181 13855
rect 51181 13821 51215 13855
rect 51215 13821 51224 13855
rect 51172 13812 51224 13821
rect 51816 13812 51868 13864
rect 51724 13744 51776 13796
rect 52552 13880 52604 13932
rect 48780 13676 48832 13728
rect 51356 13676 51408 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 23204 13472 23256 13524
rect 23940 13515 23992 13524
rect 23940 13481 23949 13515
rect 23949 13481 23983 13515
rect 23983 13481 23992 13515
rect 23940 13472 23992 13481
rect 29736 13472 29788 13524
rect 33324 13472 33376 13524
rect 39212 13515 39264 13524
rect 39212 13481 39221 13515
rect 39221 13481 39255 13515
rect 39255 13481 39264 13515
rect 39212 13472 39264 13481
rect 39580 13472 39632 13524
rect 39672 13472 39724 13524
rect 24952 13447 25004 13456
rect 24952 13413 24961 13447
rect 24961 13413 24995 13447
rect 24995 13413 25004 13447
rect 24952 13404 25004 13413
rect 27068 13336 27120 13388
rect 940 13268 992 13320
rect 22376 13268 22428 13320
rect 23572 13311 23624 13320
rect 23572 13277 23581 13311
rect 23581 13277 23615 13311
rect 23615 13277 23624 13311
rect 23572 13268 23624 13277
rect 23848 13311 23900 13320
rect 23848 13277 23857 13311
rect 23857 13277 23891 13311
rect 23891 13277 23900 13311
rect 23848 13268 23900 13277
rect 30104 13336 30156 13388
rect 31484 13336 31536 13388
rect 31668 13336 31720 13388
rect 24860 13243 24912 13252
rect 24860 13209 24869 13243
rect 24869 13209 24903 13243
rect 24903 13209 24912 13243
rect 24860 13200 24912 13209
rect 25044 13243 25096 13252
rect 25044 13209 25053 13243
rect 25053 13209 25087 13243
rect 25087 13209 25096 13243
rect 25044 13200 25096 13209
rect 25320 13200 25372 13252
rect 25780 13243 25832 13252
rect 25780 13209 25789 13243
rect 25789 13209 25823 13243
rect 25823 13209 25832 13243
rect 25780 13200 25832 13209
rect 26516 13200 26568 13252
rect 30012 13311 30064 13320
rect 30012 13277 30021 13311
rect 30021 13277 30055 13311
rect 30055 13277 30064 13311
rect 30012 13268 30064 13277
rect 31944 13336 31996 13388
rect 32220 13311 32272 13320
rect 32220 13277 32229 13311
rect 32229 13277 32263 13311
rect 32263 13277 32272 13311
rect 32220 13268 32272 13277
rect 32404 13311 32456 13320
rect 32404 13277 32413 13311
rect 32413 13277 32447 13311
rect 32447 13277 32456 13311
rect 32404 13268 32456 13277
rect 32496 13268 32548 13320
rect 38844 13336 38896 13388
rect 33048 13268 33100 13320
rect 40500 13472 40552 13524
rect 44824 13472 44876 13524
rect 40868 13404 40920 13456
rect 39856 13311 39908 13320
rect 25504 13132 25556 13184
rect 26700 13132 26752 13184
rect 32864 13200 32916 13252
rect 34060 13200 34112 13252
rect 36268 13200 36320 13252
rect 37648 13200 37700 13252
rect 30564 13175 30616 13184
rect 30564 13141 30573 13175
rect 30573 13141 30607 13175
rect 30607 13141 30616 13175
rect 30564 13132 30616 13141
rect 32128 13132 32180 13184
rect 34428 13132 34480 13184
rect 36452 13175 36504 13184
rect 36452 13141 36461 13175
rect 36461 13141 36495 13175
rect 36495 13141 36504 13175
rect 36452 13132 36504 13141
rect 39856 13277 39865 13311
rect 39865 13277 39899 13311
rect 39899 13277 39908 13311
rect 39856 13268 39908 13277
rect 41052 13200 41104 13252
rect 42524 13336 42576 13388
rect 48228 13472 48280 13524
rect 47216 13447 47268 13456
rect 47216 13413 47225 13447
rect 47225 13413 47259 13447
rect 47259 13413 47268 13447
rect 47216 13404 47268 13413
rect 47952 13404 48004 13456
rect 48136 13404 48188 13456
rect 48780 13515 48832 13524
rect 48780 13481 48789 13515
rect 48789 13481 48823 13515
rect 48823 13481 48832 13515
rect 48780 13472 48832 13481
rect 49792 13515 49844 13524
rect 49792 13481 49801 13515
rect 49801 13481 49835 13515
rect 49835 13481 49844 13515
rect 49792 13472 49844 13481
rect 51448 13472 51500 13524
rect 51724 13472 51776 13524
rect 49148 13404 49200 13456
rect 46112 13336 46164 13388
rect 42248 13268 42300 13320
rect 42340 13311 42392 13320
rect 42340 13277 42349 13311
rect 42349 13277 42383 13311
rect 42383 13277 42392 13311
rect 42340 13268 42392 13277
rect 42984 13311 43036 13320
rect 42984 13277 42993 13311
rect 42993 13277 43027 13311
rect 43027 13277 43036 13311
rect 42984 13268 43036 13277
rect 46756 13268 46808 13320
rect 47952 13311 48004 13320
rect 47952 13277 47961 13311
rect 47961 13277 47995 13311
rect 47995 13277 48004 13311
rect 47952 13268 48004 13277
rect 48228 13311 48280 13320
rect 48228 13277 48237 13311
rect 48237 13277 48271 13311
rect 48271 13277 48280 13311
rect 48228 13268 48280 13277
rect 44548 13200 44600 13252
rect 45744 13243 45796 13252
rect 45744 13209 45753 13243
rect 45753 13209 45787 13243
rect 45787 13209 45796 13243
rect 45744 13200 45796 13209
rect 39948 13132 40000 13184
rect 42432 13132 42484 13184
rect 47308 13132 47360 13184
rect 48320 13200 48372 13252
rect 48596 13311 48648 13320
rect 48596 13277 48605 13311
rect 48605 13277 48639 13311
rect 48639 13277 48648 13311
rect 48596 13268 48648 13277
rect 48872 13311 48924 13320
rect 48872 13277 48881 13311
rect 48881 13277 48915 13311
rect 48915 13277 48924 13311
rect 48872 13268 48924 13277
rect 48780 13132 48832 13184
rect 48964 13132 49016 13184
rect 49240 13268 49292 13320
rect 49332 13268 49384 13320
rect 50988 13404 51040 13456
rect 51632 13404 51684 13456
rect 50620 13336 50672 13388
rect 50896 13379 50948 13388
rect 50896 13345 50905 13379
rect 50905 13345 50939 13379
rect 50939 13345 50948 13379
rect 50896 13336 50948 13345
rect 49700 13200 49752 13252
rect 50252 13268 50304 13320
rect 51172 13268 51224 13320
rect 51356 13311 51408 13320
rect 51356 13277 51365 13311
rect 51365 13277 51399 13311
rect 51399 13277 51408 13311
rect 51356 13268 51408 13277
rect 51540 13311 51592 13320
rect 51540 13277 51549 13311
rect 51549 13277 51583 13311
rect 51583 13277 51592 13311
rect 51540 13268 51592 13277
rect 52000 13311 52052 13320
rect 52000 13277 52009 13311
rect 52009 13277 52043 13311
rect 52043 13277 52052 13311
rect 52000 13268 52052 13277
rect 51448 13200 51500 13252
rect 49976 13132 50028 13184
rect 50068 13132 50120 13184
rect 53564 13200 53616 13252
rect 53748 13175 53800 13184
rect 53748 13141 53757 13175
rect 53757 13141 53791 13175
rect 53791 13141 53800 13175
rect 53748 13132 53800 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 23572 12928 23624 12980
rect 25044 12928 25096 12980
rect 26700 12971 26752 12980
rect 26700 12937 26709 12971
rect 26709 12937 26743 12971
rect 26743 12937 26752 12971
rect 26700 12928 26752 12937
rect 30012 12928 30064 12980
rect 30564 12928 30616 12980
rect 23664 12860 23716 12912
rect 24860 12792 24912 12844
rect 22376 12724 22428 12776
rect 24492 12724 24544 12776
rect 25228 12767 25280 12776
rect 25228 12733 25237 12767
rect 25237 12733 25271 12767
rect 25271 12733 25280 12767
rect 25228 12724 25280 12733
rect 25320 12724 25372 12776
rect 27068 12792 27120 12844
rect 27804 12835 27856 12844
rect 27804 12801 27838 12835
rect 27838 12801 27856 12835
rect 27804 12792 27856 12801
rect 29000 12835 29052 12844
rect 29000 12801 29009 12835
rect 29009 12801 29043 12835
rect 29043 12801 29052 12835
rect 29000 12792 29052 12801
rect 30932 12928 30984 12980
rect 31208 12971 31260 12980
rect 31208 12937 31217 12971
rect 31217 12937 31251 12971
rect 31251 12937 31260 12971
rect 31208 12928 31260 12937
rect 25504 12656 25556 12708
rect 26884 12656 26936 12708
rect 30472 12656 30524 12708
rect 31116 12835 31168 12844
rect 31116 12801 31125 12835
rect 31125 12801 31159 12835
rect 31159 12801 31168 12835
rect 31116 12792 31168 12801
rect 32036 12860 32088 12912
rect 32404 12928 32456 12980
rect 32864 12928 32916 12980
rect 33968 12928 34020 12980
rect 34060 12971 34112 12980
rect 34060 12937 34069 12971
rect 34069 12937 34103 12971
rect 34103 12937 34112 12971
rect 34060 12928 34112 12937
rect 34152 12928 34204 12980
rect 34428 12903 34480 12912
rect 34428 12869 34437 12903
rect 34437 12869 34471 12903
rect 34471 12869 34480 12903
rect 34428 12860 34480 12869
rect 34612 12903 34664 12912
rect 34612 12869 34647 12903
rect 34647 12869 34664 12903
rect 34612 12860 34664 12869
rect 34796 12860 34848 12912
rect 36268 12971 36320 12980
rect 36268 12937 36277 12971
rect 36277 12937 36311 12971
rect 36311 12937 36320 12971
rect 36268 12928 36320 12937
rect 36452 12860 36504 12912
rect 36820 12903 36872 12912
rect 36820 12869 36855 12903
rect 36855 12869 36872 12903
rect 37648 12971 37700 12980
rect 37648 12937 37657 12971
rect 37657 12937 37691 12971
rect 37691 12937 37700 12971
rect 37648 12928 37700 12937
rect 38660 12928 38712 12980
rect 36820 12860 36872 12869
rect 31392 12724 31444 12776
rect 31668 12724 31720 12776
rect 31944 12724 31996 12776
rect 33876 12792 33928 12844
rect 33968 12792 34020 12844
rect 26240 12631 26292 12640
rect 26240 12597 26249 12631
rect 26249 12597 26283 12631
rect 26283 12597 26292 12631
rect 26240 12588 26292 12597
rect 26332 12631 26384 12640
rect 26332 12597 26341 12631
rect 26341 12597 26375 12631
rect 26375 12597 26384 12631
rect 26332 12588 26384 12597
rect 26700 12588 26752 12640
rect 27436 12631 27488 12640
rect 27436 12597 27445 12631
rect 27445 12597 27479 12631
rect 27479 12597 27488 12631
rect 27436 12588 27488 12597
rect 29276 12588 29328 12640
rect 31576 12588 31628 12640
rect 33784 12656 33836 12708
rect 34520 12656 34572 12708
rect 36728 12835 36780 12844
rect 36728 12801 36737 12835
rect 36737 12801 36771 12835
rect 36771 12801 36780 12835
rect 36728 12792 36780 12801
rect 37004 12835 37056 12844
rect 37004 12801 37013 12835
rect 37013 12801 37047 12835
rect 37047 12801 37056 12835
rect 37004 12792 37056 12801
rect 37280 12835 37332 12844
rect 37280 12801 37289 12835
rect 37289 12801 37323 12835
rect 37323 12801 37332 12835
rect 37280 12792 37332 12801
rect 37464 12835 37516 12844
rect 37464 12801 37473 12835
rect 37473 12801 37507 12835
rect 37507 12801 37516 12835
rect 37464 12792 37516 12801
rect 37832 12835 37884 12844
rect 37832 12801 37841 12835
rect 37841 12801 37875 12835
rect 37875 12801 37884 12835
rect 37832 12792 37884 12801
rect 37924 12835 37976 12844
rect 37924 12801 37933 12835
rect 37933 12801 37967 12835
rect 37967 12801 37976 12835
rect 37924 12792 37976 12801
rect 38752 12860 38804 12912
rect 39212 12792 39264 12844
rect 40224 12928 40276 12980
rect 41052 12971 41104 12980
rect 41052 12937 41061 12971
rect 41061 12937 41095 12971
rect 41095 12937 41104 12971
rect 41052 12928 41104 12937
rect 39948 12903 40000 12912
rect 39948 12869 39957 12903
rect 39957 12869 39991 12903
rect 39991 12869 40000 12903
rect 39948 12860 40000 12869
rect 42340 12928 42392 12980
rect 44548 12971 44600 12980
rect 44548 12937 44557 12971
rect 44557 12937 44591 12971
rect 44591 12937 44600 12971
rect 44548 12928 44600 12937
rect 45744 12928 45796 12980
rect 48228 12928 48280 12980
rect 51356 12928 51408 12980
rect 53564 12971 53616 12980
rect 53564 12937 53573 12971
rect 53573 12937 53607 12971
rect 53607 12937 53616 12971
rect 53564 12928 53616 12937
rect 53748 12928 53800 12980
rect 44180 12903 44232 12912
rect 44180 12869 44189 12903
rect 44189 12869 44223 12903
rect 44223 12869 44232 12903
rect 44180 12860 44232 12869
rect 44916 12860 44968 12912
rect 48412 12860 48464 12912
rect 51632 12860 51684 12912
rect 40040 12835 40092 12844
rect 40040 12801 40050 12835
rect 40050 12801 40084 12835
rect 40084 12801 40092 12835
rect 40040 12792 40092 12801
rect 40132 12835 40184 12844
rect 40132 12801 40167 12835
rect 40167 12801 40184 12835
rect 40132 12792 40184 12801
rect 41236 12792 41288 12844
rect 42156 12792 42208 12844
rect 42248 12792 42300 12844
rect 44732 12792 44784 12844
rect 45836 12792 45888 12844
rect 46480 12792 46532 12844
rect 49148 12792 49200 12844
rect 36728 12656 36780 12708
rect 32772 12631 32824 12640
rect 32772 12597 32781 12631
rect 32781 12597 32815 12631
rect 32815 12597 32824 12631
rect 32772 12588 32824 12597
rect 33232 12631 33284 12640
rect 33232 12597 33241 12631
rect 33241 12597 33275 12631
rect 33275 12597 33284 12631
rect 33232 12588 33284 12597
rect 35900 12588 35952 12640
rect 38660 12656 38712 12708
rect 37280 12631 37332 12640
rect 37280 12597 37289 12631
rect 37289 12597 37323 12631
rect 37323 12597 37332 12631
rect 37280 12588 37332 12597
rect 38292 12588 38344 12640
rect 38936 12656 38988 12708
rect 39764 12588 39816 12640
rect 40776 12588 40828 12640
rect 46388 12724 46440 12776
rect 48228 12767 48280 12776
rect 48228 12733 48237 12767
rect 48237 12733 48271 12767
rect 48271 12733 48280 12767
rect 48228 12724 48280 12733
rect 48964 12724 49016 12776
rect 49332 12767 49384 12776
rect 49332 12733 49341 12767
rect 49341 12733 49375 12767
rect 49375 12733 49384 12767
rect 49332 12724 49384 12733
rect 49700 12724 49752 12776
rect 42800 12588 42852 12640
rect 46112 12656 46164 12708
rect 50068 12835 50120 12844
rect 50068 12801 50077 12835
rect 50077 12801 50111 12835
rect 50111 12801 50120 12835
rect 50068 12792 50120 12801
rect 50528 12792 50580 12844
rect 50896 12792 50948 12844
rect 52184 12792 52236 12844
rect 53472 12835 53524 12844
rect 53472 12801 53481 12835
rect 53481 12801 53515 12835
rect 53515 12801 53524 12835
rect 53472 12792 53524 12801
rect 49976 12767 50028 12776
rect 49976 12733 49985 12767
rect 49985 12733 50019 12767
rect 50019 12733 50028 12767
rect 49976 12724 50028 12733
rect 51264 12767 51316 12776
rect 51264 12733 51273 12767
rect 51273 12733 51307 12767
rect 51307 12733 51316 12767
rect 51264 12724 51316 12733
rect 51540 12724 51592 12776
rect 49608 12588 49660 12640
rect 51816 12631 51868 12640
rect 51816 12597 51825 12631
rect 51825 12597 51859 12631
rect 51859 12597 51868 12631
rect 51816 12588 51868 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 23664 12427 23716 12436
rect 23664 12393 23673 12427
rect 23673 12393 23707 12427
rect 23707 12393 23716 12427
rect 23664 12384 23716 12393
rect 24492 12427 24544 12436
rect 24492 12393 24501 12427
rect 24501 12393 24535 12427
rect 24535 12393 24544 12427
rect 24492 12384 24544 12393
rect 26516 12384 26568 12436
rect 29368 12384 29420 12436
rect 23848 12180 23900 12232
rect 26332 12316 26384 12368
rect 24952 12248 25004 12300
rect 26240 12248 26292 12300
rect 29276 12248 29328 12300
rect 25228 12180 25280 12232
rect 24860 12155 24912 12164
rect 24860 12121 24869 12155
rect 24869 12121 24903 12155
rect 24903 12121 24912 12155
rect 24860 12112 24912 12121
rect 23572 12044 23624 12096
rect 27436 12223 27488 12232
rect 27436 12189 27445 12223
rect 27445 12189 27479 12223
rect 27479 12189 27488 12223
rect 27436 12180 27488 12189
rect 32312 12384 32364 12436
rect 32680 12384 32732 12436
rect 32956 12384 33008 12436
rect 34612 12384 34664 12436
rect 37372 12384 37424 12436
rect 38660 12384 38712 12436
rect 31484 12316 31536 12368
rect 30932 12248 30984 12300
rect 31668 12248 31720 12300
rect 33140 12291 33192 12300
rect 33140 12257 33149 12291
rect 33149 12257 33183 12291
rect 33183 12257 33192 12291
rect 33140 12248 33192 12257
rect 37004 12316 37056 12368
rect 38936 12316 38988 12368
rect 48228 12384 48280 12436
rect 51264 12427 51316 12436
rect 51264 12393 51273 12427
rect 51273 12393 51307 12427
rect 51307 12393 51316 12427
rect 51264 12384 51316 12393
rect 51448 12427 51500 12436
rect 51448 12393 51457 12427
rect 51457 12393 51491 12427
rect 51491 12393 51500 12427
rect 51448 12384 51500 12393
rect 40592 12316 40644 12368
rect 28632 12112 28684 12164
rect 30380 12223 30432 12232
rect 30380 12189 30389 12223
rect 30389 12189 30423 12223
rect 30423 12189 30432 12223
rect 30380 12180 30432 12189
rect 30840 12180 30892 12232
rect 32404 12180 32456 12232
rect 32864 12223 32916 12232
rect 32864 12189 32873 12223
rect 32873 12189 32907 12223
rect 32907 12189 32916 12223
rect 32864 12180 32916 12189
rect 32956 12223 33008 12232
rect 32956 12189 32965 12223
rect 32965 12189 32999 12223
rect 32999 12189 33008 12223
rect 32956 12180 33008 12189
rect 33600 12223 33652 12232
rect 33600 12189 33609 12223
rect 33609 12189 33643 12223
rect 33643 12189 33652 12223
rect 33600 12180 33652 12189
rect 37280 12248 37332 12300
rect 37464 12248 37516 12300
rect 39396 12248 39448 12300
rect 43076 12291 43128 12300
rect 43076 12257 43085 12291
rect 43085 12257 43119 12291
rect 43119 12257 43128 12291
rect 43076 12248 43128 12257
rect 46112 12248 46164 12300
rect 47124 12248 47176 12300
rect 27436 12044 27488 12096
rect 29276 12087 29328 12096
rect 29276 12053 29285 12087
rect 29285 12053 29319 12087
rect 29319 12053 29328 12087
rect 29276 12044 29328 12053
rect 30196 12087 30248 12096
rect 30196 12053 30205 12087
rect 30205 12053 30239 12087
rect 30239 12053 30248 12087
rect 30196 12044 30248 12053
rect 31668 12087 31720 12096
rect 31668 12053 31677 12087
rect 31677 12053 31711 12087
rect 31711 12053 31720 12087
rect 31668 12044 31720 12053
rect 32680 12087 32732 12096
rect 32680 12053 32689 12087
rect 32689 12053 32723 12087
rect 32723 12053 32732 12087
rect 32680 12044 32732 12053
rect 32864 12044 32916 12096
rect 33692 12087 33744 12096
rect 33692 12053 33701 12087
rect 33701 12053 33735 12087
rect 33735 12053 33744 12087
rect 33692 12044 33744 12053
rect 34796 12180 34848 12232
rect 50528 12291 50580 12300
rect 50528 12257 50537 12291
rect 50537 12257 50571 12291
rect 50571 12257 50580 12291
rect 50528 12248 50580 12257
rect 51448 12248 51500 12300
rect 35072 12112 35124 12164
rect 35164 12044 35216 12096
rect 35900 12044 35952 12096
rect 37832 12223 37884 12232
rect 37832 12189 37841 12223
rect 37841 12189 37875 12223
rect 37875 12189 37884 12223
rect 37832 12180 37884 12189
rect 36360 12112 36412 12164
rect 38016 12112 38068 12164
rect 38844 12180 38896 12232
rect 38936 12180 38988 12232
rect 40224 12180 40276 12232
rect 40684 12223 40736 12232
rect 40684 12189 40693 12223
rect 40693 12189 40727 12223
rect 40727 12189 40736 12223
rect 40684 12180 40736 12189
rect 40868 12223 40920 12232
rect 40868 12189 40877 12223
rect 40877 12189 40911 12223
rect 40911 12189 40920 12223
rect 40868 12180 40920 12189
rect 41236 12180 41288 12232
rect 42248 12180 42300 12232
rect 44916 12180 44968 12232
rect 49976 12180 50028 12232
rect 36912 12087 36964 12096
rect 36912 12053 36921 12087
rect 36921 12053 36955 12087
rect 36955 12053 36964 12087
rect 36912 12044 36964 12053
rect 38752 12044 38804 12096
rect 40408 12087 40460 12096
rect 40408 12053 40423 12087
rect 40423 12053 40457 12087
rect 40457 12053 40460 12087
rect 40408 12044 40460 12053
rect 40592 12044 40644 12096
rect 40776 12087 40828 12096
rect 40776 12053 40785 12087
rect 40785 12053 40819 12087
rect 40819 12053 40828 12087
rect 40776 12044 40828 12053
rect 41604 12087 41656 12096
rect 41604 12053 41613 12087
rect 41613 12053 41647 12087
rect 41647 12053 41656 12087
rect 41604 12044 41656 12053
rect 43352 12155 43404 12164
rect 43352 12121 43361 12155
rect 43361 12121 43395 12155
rect 43395 12121 43404 12155
rect 43352 12112 43404 12121
rect 47124 12112 47176 12164
rect 49332 12112 49384 12164
rect 50988 12112 51040 12164
rect 44732 12044 44784 12096
rect 44824 12087 44876 12096
rect 44824 12053 44833 12087
rect 44833 12053 44867 12087
rect 44867 12053 44876 12087
rect 44824 12044 44876 12053
rect 50160 12087 50212 12096
rect 50160 12053 50169 12087
rect 50169 12053 50203 12087
rect 50203 12053 50212 12087
rect 50160 12044 50212 12053
rect 50620 12044 50672 12096
rect 52092 12112 52144 12164
rect 51448 12044 51500 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 25780 11840 25832 11892
rect 27160 11840 27212 11892
rect 29276 11840 29328 11892
rect 30380 11840 30432 11892
rect 31668 11840 31720 11892
rect 32312 11840 32364 11892
rect 33692 11840 33744 11892
rect 35072 11840 35124 11892
rect 25688 11704 25740 11756
rect 26700 11772 26752 11824
rect 26884 11772 26936 11824
rect 30932 11815 30984 11824
rect 30932 11781 30941 11815
rect 30941 11781 30975 11815
rect 30975 11781 30984 11815
rect 30932 11772 30984 11781
rect 31392 11772 31444 11824
rect 26424 11747 26476 11756
rect 26424 11713 26459 11747
rect 26459 11713 26476 11747
rect 26424 11704 26476 11713
rect 28080 11747 28132 11756
rect 28080 11713 28089 11747
rect 28089 11713 28123 11747
rect 28123 11713 28132 11747
rect 28080 11704 28132 11713
rect 31208 11747 31260 11756
rect 31208 11713 31217 11747
rect 31217 11713 31251 11747
rect 31251 11713 31260 11747
rect 31208 11704 31260 11713
rect 29000 11636 29052 11688
rect 31484 11747 31536 11756
rect 31484 11713 31493 11747
rect 31493 11713 31527 11747
rect 31527 11713 31536 11747
rect 31484 11704 31536 11713
rect 32680 11704 32732 11756
rect 36360 11840 36412 11892
rect 36912 11840 36964 11892
rect 34612 11704 34664 11756
rect 35164 11704 35216 11756
rect 35808 11704 35860 11756
rect 36084 11747 36136 11756
rect 36084 11713 36093 11747
rect 36093 11713 36127 11747
rect 36127 11713 36136 11747
rect 36084 11704 36136 11713
rect 37740 11840 37792 11892
rect 37832 11840 37884 11892
rect 41604 11840 41656 11892
rect 42156 11883 42208 11892
rect 42156 11849 42165 11883
rect 42165 11849 42199 11883
rect 42199 11849 42208 11883
rect 42156 11840 42208 11849
rect 43352 11840 43404 11892
rect 47124 11883 47176 11892
rect 47124 11849 47133 11883
rect 47133 11849 47167 11883
rect 47167 11849 47176 11883
rect 47124 11840 47176 11849
rect 49332 11883 49384 11892
rect 49332 11849 49341 11883
rect 49341 11849 49375 11883
rect 49375 11849 49384 11883
rect 49332 11840 49384 11849
rect 40592 11772 40644 11824
rect 38752 11704 38804 11756
rect 38844 11747 38896 11756
rect 38844 11713 38853 11747
rect 38853 11713 38887 11747
rect 38887 11713 38896 11747
rect 38844 11704 38896 11713
rect 39120 11747 39172 11756
rect 39120 11713 39154 11747
rect 39154 11713 39172 11747
rect 39120 11704 39172 11713
rect 40408 11747 40460 11756
rect 40408 11713 40417 11747
rect 40417 11713 40451 11747
rect 40451 11713 40460 11747
rect 40408 11704 40460 11713
rect 44732 11772 44784 11824
rect 32220 11636 32272 11688
rect 32588 11636 32640 11688
rect 33048 11679 33100 11688
rect 33048 11645 33057 11679
rect 33057 11645 33091 11679
rect 33091 11645 33100 11679
rect 33048 11636 33100 11645
rect 24860 11543 24912 11552
rect 24860 11509 24869 11543
rect 24869 11509 24903 11543
rect 24903 11509 24912 11543
rect 24860 11500 24912 11509
rect 25228 11500 25280 11552
rect 26424 11500 26476 11552
rect 26608 11500 26660 11552
rect 28908 11500 28960 11552
rect 32772 11568 32824 11620
rect 30564 11500 30616 11552
rect 30840 11543 30892 11552
rect 30840 11509 30849 11543
rect 30849 11509 30883 11543
rect 30883 11509 30892 11543
rect 30840 11500 30892 11509
rect 31300 11543 31352 11552
rect 31300 11509 31309 11543
rect 31309 11509 31343 11543
rect 31343 11509 31352 11543
rect 31300 11500 31352 11509
rect 32680 11500 32732 11552
rect 33968 11500 34020 11552
rect 35808 11543 35860 11552
rect 35808 11509 35817 11543
rect 35817 11509 35851 11543
rect 35851 11509 35860 11543
rect 35808 11500 35860 11509
rect 36452 11679 36504 11688
rect 36452 11645 36461 11679
rect 36461 11645 36495 11679
rect 36495 11645 36504 11679
rect 36452 11636 36504 11645
rect 40776 11636 40828 11688
rect 41144 11636 41196 11688
rect 44456 11704 44508 11756
rect 44916 11747 44968 11756
rect 44916 11713 44925 11747
rect 44925 11713 44959 11747
rect 44959 11713 44968 11747
rect 44916 11704 44968 11713
rect 42432 11679 42484 11688
rect 42432 11645 42441 11679
rect 42441 11645 42475 11679
rect 42475 11645 42484 11679
rect 42432 11636 42484 11645
rect 36452 11500 36504 11552
rect 37004 11543 37056 11552
rect 37004 11509 37013 11543
rect 37013 11509 37047 11543
rect 37047 11509 37056 11543
rect 37004 11500 37056 11509
rect 38292 11500 38344 11552
rect 39212 11500 39264 11552
rect 44824 11636 44876 11688
rect 45100 11636 45152 11688
rect 46112 11704 46164 11756
rect 47768 11772 47820 11824
rect 50160 11840 50212 11892
rect 47216 11704 47268 11756
rect 49884 11815 49936 11824
rect 49884 11781 49893 11815
rect 49893 11781 49927 11815
rect 49927 11781 49936 11815
rect 49884 11772 49936 11781
rect 50344 11772 50396 11824
rect 50528 11772 50580 11824
rect 50988 11772 51040 11824
rect 47584 11679 47636 11688
rect 47584 11645 47593 11679
rect 47593 11645 47627 11679
rect 47627 11645 47636 11679
rect 47584 11636 47636 11645
rect 47860 11679 47912 11688
rect 47860 11645 47869 11679
rect 47869 11645 47903 11679
rect 47903 11645 47912 11679
rect 47860 11636 47912 11645
rect 49608 11568 49660 11620
rect 50436 11636 50488 11688
rect 51448 11840 51500 11892
rect 52184 11840 52236 11892
rect 52092 11772 52144 11824
rect 51540 11747 51592 11756
rect 51540 11713 51549 11747
rect 51549 11713 51583 11747
rect 51583 11713 51592 11747
rect 51540 11704 51592 11713
rect 51908 11747 51960 11756
rect 51908 11713 51917 11747
rect 51917 11713 51951 11747
rect 51951 11713 51960 11747
rect 51908 11704 51960 11713
rect 52276 11704 52328 11756
rect 41696 11543 41748 11552
rect 41696 11509 41705 11543
rect 41705 11509 41739 11543
rect 41739 11509 41748 11543
rect 41696 11500 41748 11509
rect 41880 11500 41932 11552
rect 49516 11543 49568 11552
rect 49516 11509 49525 11543
rect 49525 11509 49559 11543
rect 49559 11509 49568 11543
rect 49516 11500 49568 11509
rect 51264 11543 51316 11552
rect 51264 11509 51273 11543
rect 51273 11509 51307 11543
rect 51307 11509 51316 11543
rect 51264 11500 51316 11509
rect 51724 11568 51776 11620
rect 68468 11611 68520 11620
rect 68468 11577 68477 11611
rect 68477 11577 68511 11611
rect 68511 11577 68520 11611
rect 68468 11568 68520 11577
rect 51816 11500 51868 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 22376 11203 22428 11212
rect 22376 11169 22385 11203
rect 22385 11169 22419 11203
rect 22419 11169 22428 11203
rect 22376 11160 22428 11169
rect 24400 11160 24452 11212
rect 25504 11160 25556 11212
rect 25964 11160 26016 11212
rect 26516 11296 26568 11348
rect 26608 11339 26660 11348
rect 26608 11305 26617 11339
rect 26617 11305 26651 11339
rect 26651 11305 26660 11339
rect 26608 11296 26660 11305
rect 27160 11339 27212 11348
rect 27160 11305 27169 11339
rect 27169 11305 27203 11339
rect 27203 11305 27212 11339
rect 27160 11296 27212 11305
rect 28080 11296 28132 11348
rect 28356 11339 28408 11348
rect 28356 11305 28365 11339
rect 28365 11305 28399 11339
rect 28399 11305 28408 11339
rect 28356 11296 28408 11305
rect 28632 11296 28684 11348
rect 23664 11024 23716 11076
rect 25136 11092 25188 11144
rect 25320 11092 25372 11144
rect 25780 11135 25832 11144
rect 25780 11101 25789 11135
rect 25789 11101 25823 11135
rect 25823 11101 25832 11135
rect 25780 11092 25832 11101
rect 25872 11135 25924 11144
rect 25872 11101 25881 11135
rect 25881 11101 25915 11135
rect 25915 11101 25924 11135
rect 25872 11092 25924 11101
rect 26056 11135 26108 11144
rect 26056 11101 26065 11135
rect 26065 11101 26099 11135
rect 26099 11101 26108 11135
rect 26056 11092 26108 11101
rect 26240 11203 26292 11212
rect 26240 11169 26249 11203
rect 26249 11169 26283 11203
rect 26283 11169 26292 11203
rect 26240 11160 26292 11169
rect 26424 11135 26476 11144
rect 26424 11101 26433 11135
rect 26433 11101 26467 11135
rect 26467 11101 26476 11135
rect 26424 11092 26476 11101
rect 25504 11024 25556 11076
rect 26792 11024 26844 11076
rect 25044 10956 25096 11008
rect 25412 10999 25464 11008
rect 25412 10965 25421 10999
rect 25421 10965 25455 10999
rect 25455 10965 25464 10999
rect 25412 10956 25464 10965
rect 25780 10956 25832 11008
rect 26240 10956 26292 11008
rect 27344 11135 27396 11144
rect 27344 11101 27353 11135
rect 27353 11101 27387 11135
rect 27387 11101 27396 11135
rect 27344 11092 27396 11101
rect 27436 11135 27488 11144
rect 27436 11101 27445 11135
rect 27445 11101 27479 11135
rect 27479 11101 27488 11135
rect 27436 11092 27488 11101
rect 28080 11092 28132 11144
rect 28356 11092 28408 11144
rect 28540 11135 28592 11144
rect 28540 11101 28549 11135
rect 28549 11101 28583 11135
rect 28583 11101 28592 11135
rect 28540 11092 28592 11101
rect 30012 11092 30064 11144
rect 30564 11228 30616 11280
rect 32680 11228 32732 11280
rect 30564 11135 30616 11144
rect 30564 11101 30573 11135
rect 30573 11101 30607 11135
rect 30607 11101 30616 11135
rect 30564 11092 30616 11101
rect 31392 11092 31444 11144
rect 32588 11092 32640 11144
rect 28172 10956 28224 11008
rect 30656 11024 30708 11076
rect 30748 11024 30800 11076
rect 35808 11296 35860 11348
rect 35900 11296 35952 11348
rect 38936 11296 38988 11348
rect 39120 11296 39172 11348
rect 39764 11296 39816 11348
rect 41236 11339 41288 11348
rect 41236 11305 41245 11339
rect 41245 11305 41279 11339
rect 41279 11305 41288 11339
rect 41236 11296 41288 11305
rect 47860 11296 47912 11348
rect 50620 11296 50672 11348
rect 51264 11296 51316 11348
rect 51356 11296 51408 11348
rect 47032 11228 47084 11280
rect 47768 11271 47820 11280
rect 47768 11237 47777 11271
rect 47777 11237 47811 11271
rect 47811 11237 47820 11271
rect 47768 11228 47820 11237
rect 34796 11135 34848 11144
rect 34796 11101 34805 11135
rect 34805 11101 34839 11135
rect 34839 11101 34848 11135
rect 34796 11092 34848 11101
rect 38844 11160 38896 11212
rect 39856 11203 39908 11212
rect 39856 11169 39865 11203
rect 39865 11169 39899 11203
rect 39899 11169 39908 11203
rect 39856 11160 39908 11169
rect 37464 11092 37516 11144
rect 37924 11135 37976 11144
rect 37924 11101 37933 11135
rect 37933 11101 37967 11135
rect 37967 11101 37976 11135
rect 37924 11092 37976 11101
rect 37372 11024 37424 11076
rect 38108 11135 38160 11144
rect 38108 11101 38117 11135
rect 38117 11101 38151 11135
rect 38151 11101 38160 11135
rect 38108 11092 38160 11101
rect 38292 11092 38344 11144
rect 39212 11135 39264 11144
rect 39212 11101 39221 11135
rect 39221 11101 39255 11135
rect 39255 11101 39264 11135
rect 39212 11092 39264 11101
rect 39396 11135 39448 11144
rect 39396 11101 39405 11135
rect 39405 11101 39439 11135
rect 39439 11101 39448 11135
rect 39396 11092 39448 11101
rect 41328 11092 41380 11144
rect 45560 11160 45612 11212
rect 46020 11160 46072 11212
rect 46388 11135 46440 11144
rect 46388 11101 46397 11135
rect 46397 11101 46431 11135
rect 46431 11101 46440 11135
rect 46388 11092 46440 11101
rect 48320 11160 48372 11212
rect 49976 11160 50028 11212
rect 32772 10956 32824 11008
rect 32864 10956 32916 11008
rect 37096 10956 37148 11008
rect 40132 11067 40184 11076
rect 40132 11033 40166 11067
rect 40166 11033 40184 11067
rect 40132 11024 40184 11033
rect 41696 11024 41748 11076
rect 43076 11024 43128 11076
rect 45836 11024 45888 11076
rect 47216 11024 47268 11076
rect 49332 11092 49384 11144
rect 52000 11160 52052 11212
rect 52276 11160 52328 11212
rect 49608 11024 49660 11076
rect 37648 10999 37700 11008
rect 37648 10965 37657 10999
rect 37657 10965 37691 10999
rect 37691 10965 37700 10999
rect 37648 10956 37700 10965
rect 42524 10956 42576 11008
rect 43168 10999 43220 11008
rect 43168 10965 43177 10999
rect 43177 10965 43211 10999
rect 43211 10965 43220 10999
rect 43168 10956 43220 10965
rect 49240 10956 49292 11008
rect 51448 11024 51500 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 23664 10752 23716 10804
rect 24400 10795 24452 10804
rect 24400 10761 24409 10795
rect 24409 10761 24443 10795
rect 24443 10761 24452 10795
rect 24400 10752 24452 10761
rect 24860 10752 24912 10804
rect 25320 10795 25372 10804
rect 25320 10761 25329 10795
rect 25329 10761 25363 10795
rect 25363 10761 25372 10795
rect 25320 10752 25372 10761
rect 25504 10795 25556 10804
rect 25504 10761 25513 10795
rect 25513 10761 25547 10795
rect 25547 10761 25556 10795
rect 25504 10752 25556 10761
rect 25688 10795 25740 10804
rect 25688 10761 25697 10795
rect 25697 10761 25731 10795
rect 25731 10761 25740 10795
rect 25688 10752 25740 10761
rect 26424 10752 26476 10804
rect 26792 10795 26844 10804
rect 26792 10761 26801 10795
rect 26801 10761 26835 10795
rect 26835 10761 26844 10795
rect 26792 10752 26844 10761
rect 27344 10795 27396 10804
rect 27344 10761 27353 10795
rect 27353 10761 27387 10795
rect 27387 10761 27396 10795
rect 27344 10752 27396 10761
rect 28448 10752 28500 10804
rect 33600 10752 33652 10804
rect 38568 10752 38620 10804
rect 41144 10752 41196 10804
rect 25228 10684 25280 10736
rect 25964 10684 26016 10736
rect 26056 10684 26108 10736
rect 26332 10684 26384 10736
rect 23664 10616 23716 10668
rect 940 10412 992 10464
rect 24768 10659 24820 10668
rect 24768 10625 24777 10659
rect 24777 10625 24811 10659
rect 24811 10625 24820 10659
rect 24768 10616 24820 10625
rect 25780 10659 25832 10668
rect 25780 10625 25789 10659
rect 25789 10625 25823 10659
rect 25823 10625 25832 10659
rect 25780 10616 25832 10625
rect 25872 10616 25924 10668
rect 25044 10591 25096 10600
rect 25044 10557 25053 10591
rect 25053 10557 25087 10591
rect 25087 10557 25096 10591
rect 25044 10548 25096 10557
rect 25136 10591 25188 10600
rect 25136 10557 25145 10591
rect 25145 10557 25179 10591
rect 25179 10557 25188 10591
rect 25136 10548 25188 10557
rect 25412 10480 25464 10532
rect 25504 10412 25556 10464
rect 27528 10727 27580 10736
rect 27528 10693 27537 10727
rect 27537 10693 27571 10727
rect 27571 10693 27580 10727
rect 27528 10684 27580 10693
rect 28172 10684 28224 10736
rect 29000 10684 29052 10736
rect 30196 10684 30248 10736
rect 28540 10616 28592 10668
rect 27344 10591 27396 10600
rect 27344 10557 27353 10591
rect 27353 10557 27387 10591
rect 27387 10557 27396 10591
rect 27344 10548 27396 10557
rect 28908 10548 28960 10600
rect 29276 10591 29328 10600
rect 29276 10557 29285 10591
rect 29285 10557 29319 10591
rect 29319 10557 29328 10591
rect 29276 10548 29328 10557
rect 33048 10659 33100 10668
rect 33048 10625 33057 10659
rect 33057 10625 33091 10659
rect 33091 10625 33100 10659
rect 33048 10616 33100 10625
rect 30564 10548 30616 10600
rect 34520 10616 34572 10668
rect 37004 10684 37056 10736
rect 34060 10591 34112 10600
rect 34060 10557 34069 10591
rect 34069 10557 34103 10591
rect 34103 10557 34112 10591
rect 34060 10548 34112 10557
rect 32772 10480 32824 10532
rect 35256 10548 35308 10600
rect 35808 10591 35860 10600
rect 35808 10557 35817 10591
rect 35817 10557 35851 10591
rect 35851 10557 35860 10591
rect 35808 10548 35860 10557
rect 38108 10684 38160 10736
rect 37372 10659 37424 10668
rect 37372 10625 37381 10659
rect 37381 10625 37415 10659
rect 37415 10625 37424 10659
rect 37372 10616 37424 10625
rect 37740 10616 37792 10668
rect 37832 10616 37884 10668
rect 40776 10727 40828 10736
rect 40776 10693 40785 10727
rect 40785 10693 40819 10727
rect 40819 10693 40828 10727
rect 40776 10684 40828 10693
rect 41328 10684 41380 10736
rect 43076 10795 43128 10804
rect 43076 10761 43085 10795
rect 43085 10761 43119 10795
rect 43119 10761 43128 10795
rect 43076 10752 43128 10761
rect 44364 10752 44416 10804
rect 44916 10752 44968 10804
rect 45192 10752 45244 10804
rect 50988 10795 51040 10804
rect 50988 10761 50997 10795
rect 50997 10761 51031 10795
rect 51031 10761 51040 10795
rect 50988 10752 51040 10761
rect 51448 10795 51500 10804
rect 51448 10761 51457 10795
rect 51457 10761 51491 10795
rect 51491 10761 51500 10795
rect 51448 10752 51500 10761
rect 49516 10727 49568 10736
rect 49516 10693 49525 10727
rect 49525 10693 49559 10727
rect 49559 10693 49568 10727
rect 49516 10684 49568 10693
rect 41604 10616 41656 10668
rect 41880 10659 41932 10668
rect 41880 10625 41889 10659
rect 41889 10625 41923 10659
rect 41923 10625 41932 10659
rect 41880 10616 41932 10625
rect 47584 10616 47636 10668
rect 49240 10659 49292 10668
rect 49240 10625 49249 10659
rect 49249 10625 49283 10659
rect 49283 10625 49292 10659
rect 49240 10616 49292 10625
rect 51080 10659 51132 10668
rect 51080 10625 51089 10659
rect 51089 10625 51123 10659
rect 51123 10625 51132 10659
rect 51080 10616 51132 10625
rect 39764 10548 39816 10600
rect 41328 10548 41380 10600
rect 42248 10548 42300 10600
rect 37648 10480 37700 10532
rect 37740 10480 37792 10532
rect 38292 10480 38344 10532
rect 40132 10480 40184 10532
rect 45100 10591 45152 10600
rect 45100 10557 45109 10591
rect 45109 10557 45143 10591
rect 45143 10557 45152 10591
rect 45100 10548 45152 10557
rect 45560 10548 45612 10600
rect 28356 10412 28408 10464
rect 29552 10455 29604 10464
rect 29552 10421 29561 10455
rect 29561 10421 29595 10455
rect 29595 10421 29604 10455
rect 29552 10412 29604 10421
rect 33232 10455 33284 10464
rect 33232 10421 33241 10455
rect 33241 10421 33275 10455
rect 33275 10421 33284 10455
rect 33232 10412 33284 10421
rect 33508 10412 33560 10464
rect 33692 10412 33744 10464
rect 35348 10455 35400 10464
rect 35348 10421 35357 10455
rect 35357 10421 35391 10455
rect 35391 10421 35400 10455
rect 35348 10412 35400 10421
rect 36636 10412 36688 10464
rect 38844 10412 38896 10464
rect 42156 10455 42208 10464
rect 42156 10421 42165 10455
rect 42165 10421 42199 10455
rect 42199 10421 42208 10455
rect 42156 10412 42208 10421
rect 43812 10455 43864 10464
rect 43812 10421 43821 10455
rect 43821 10421 43855 10455
rect 43855 10421 43864 10455
rect 43812 10412 43864 10421
rect 44640 10455 44692 10464
rect 44640 10421 44649 10455
rect 44649 10421 44683 10455
rect 44683 10421 44692 10455
rect 44640 10412 44692 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 26424 10208 26476 10260
rect 25780 10072 25832 10124
rect 25596 10004 25648 10056
rect 26056 10004 26108 10056
rect 27344 10208 27396 10260
rect 33048 10208 33100 10260
rect 33232 10208 33284 10260
rect 34060 10208 34112 10260
rect 42248 10208 42300 10260
rect 26792 10140 26844 10192
rect 29276 10140 29328 10192
rect 35624 10140 35676 10192
rect 26884 10047 26936 10056
rect 26884 10013 26893 10047
rect 26893 10013 26927 10047
rect 26927 10013 26936 10047
rect 26884 10004 26936 10013
rect 24860 9936 24912 9988
rect 25504 9979 25556 9988
rect 25504 9945 25513 9979
rect 25513 9945 25547 9979
rect 25547 9945 25556 9979
rect 25504 9936 25556 9945
rect 27528 10047 27580 10056
rect 27528 10013 27537 10047
rect 27537 10013 27571 10047
rect 27571 10013 27580 10047
rect 27528 10004 27580 10013
rect 30748 10072 30800 10124
rect 30932 10072 30984 10124
rect 28264 9979 28316 9988
rect 28264 9945 28273 9979
rect 28273 9945 28307 9979
rect 28307 9945 28316 9979
rect 28264 9936 28316 9945
rect 30564 10004 30616 10056
rect 31392 10004 31444 10056
rect 32772 10004 32824 10056
rect 28908 9936 28960 9988
rect 32220 9936 32272 9988
rect 33508 10047 33560 10056
rect 33508 10013 33517 10047
rect 33517 10013 33551 10047
rect 33551 10013 33560 10047
rect 33508 10004 33560 10013
rect 33600 10047 33652 10056
rect 33600 10013 33609 10047
rect 33609 10013 33643 10047
rect 33643 10013 33652 10047
rect 33600 10004 33652 10013
rect 35440 10072 35492 10124
rect 34796 10004 34848 10056
rect 37648 10004 37700 10056
rect 40592 10140 40644 10192
rect 43168 10208 43220 10260
rect 38292 10072 38344 10124
rect 39028 10072 39080 10124
rect 40040 10072 40092 10124
rect 23480 9868 23532 9920
rect 25688 9911 25740 9920
rect 25688 9877 25713 9911
rect 25713 9877 25740 9911
rect 25688 9868 25740 9877
rect 26148 9868 26200 9920
rect 26516 9868 26568 9920
rect 27436 9868 27488 9920
rect 31024 9911 31076 9920
rect 31024 9877 31033 9911
rect 31033 9877 31067 9911
rect 31067 9877 31076 9911
rect 31024 9868 31076 9877
rect 31116 9868 31168 9920
rect 34520 9936 34572 9988
rect 36728 9936 36780 9988
rect 33048 9911 33100 9920
rect 33048 9877 33057 9911
rect 33057 9877 33091 9911
rect 33091 9877 33100 9911
rect 33048 9868 33100 9877
rect 37188 9911 37240 9920
rect 37188 9877 37197 9911
rect 37197 9877 37231 9911
rect 37231 9877 37240 9911
rect 37188 9868 37240 9877
rect 37372 9911 37424 9920
rect 37372 9877 37381 9911
rect 37381 9877 37415 9911
rect 37415 9877 37424 9911
rect 37372 9868 37424 9877
rect 39580 10004 39632 10056
rect 40684 10004 40736 10056
rect 42064 10072 42116 10124
rect 42432 10183 42484 10192
rect 42432 10149 42441 10183
rect 42441 10149 42475 10183
rect 42475 10149 42484 10183
rect 42432 10140 42484 10149
rect 44916 10208 44968 10260
rect 45560 10208 45612 10260
rect 46388 10208 46440 10260
rect 41328 10047 41380 10056
rect 41328 10013 41337 10047
rect 41337 10013 41371 10047
rect 41371 10013 41380 10047
rect 41328 10004 41380 10013
rect 42248 10047 42300 10056
rect 42248 10013 42257 10047
rect 42257 10013 42291 10047
rect 42291 10013 42300 10047
rect 42248 10004 42300 10013
rect 42524 10047 42576 10056
rect 42524 10013 42533 10047
rect 42533 10013 42567 10047
rect 42567 10013 42576 10047
rect 42524 10004 42576 10013
rect 42800 10072 42852 10124
rect 38936 9868 38988 9920
rect 39120 9911 39172 9920
rect 39120 9877 39129 9911
rect 39129 9877 39163 9911
rect 39163 9877 39172 9911
rect 39120 9868 39172 9877
rect 40592 9911 40644 9920
rect 40592 9877 40601 9911
rect 40601 9877 40635 9911
rect 40635 9877 40644 9911
rect 40592 9868 40644 9877
rect 43812 10072 43864 10124
rect 43352 10047 43404 10056
rect 43352 10013 43361 10047
rect 43361 10013 43395 10047
rect 43395 10013 43404 10047
rect 43352 10004 43404 10013
rect 43904 9936 43956 9988
rect 45560 10115 45612 10124
rect 45560 10081 45569 10115
rect 45569 10081 45603 10115
rect 45603 10081 45612 10115
rect 45560 10072 45612 10081
rect 46020 10004 46072 10056
rect 47584 10072 47636 10124
rect 50160 10047 50212 10056
rect 50160 10013 50169 10047
rect 50169 10013 50203 10047
rect 50203 10013 50212 10047
rect 50160 10004 50212 10013
rect 46940 9936 46992 9988
rect 48044 9979 48096 9988
rect 48044 9945 48053 9979
rect 48053 9945 48087 9979
rect 48087 9945 48096 9979
rect 48044 9936 48096 9945
rect 45928 9868 45980 9920
rect 46480 9868 46532 9920
rect 50068 9868 50120 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 23572 9596 23624 9648
rect 24768 9664 24820 9716
rect 26148 9664 26200 9716
rect 26332 9664 26384 9716
rect 30748 9707 30800 9716
rect 30748 9673 30757 9707
rect 30757 9673 30791 9707
rect 30791 9673 30800 9707
rect 30748 9664 30800 9673
rect 30932 9707 30984 9716
rect 30932 9673 30941 9707
rect 30941 9673 30975 9707
rect 30975 9673 30984 9707
rect 30932 9664 30984 9673
rect 31024 9664 31076 9716
rect 31392 9664 31444 9716
rect 25688 9639 25740 9648
rect 25688 9605 25697 9639
rect 25697 9605 25731 9639
rect 25731 9605 25740 9639
rect 25688 9596 25740 9605
rect 25780 9596 25832 9648
rect 26056 9596 26108 9648
rect 23480 9460 23532 9512
rect 24768 9571 24820 9580
rect 24768 9537 24777 9571
rect 24777 9537 24811 9571
rect 24811 9537 24820 9571
rect 24768 9528 24820 9537
rect 24860 9571 24912 9580
rect 24860 9537 24869 9571
rect 24869 9537 24903 9571
rect 24903 9537 24912 9571
rect 24860 9528 24912 9537
rect 25228 9528 25280 9580
rect 26608 9639 26660 9648
rect 26608 9605 26617 9639
rect 26617 9605 26651 9639
rect 26651 9605 26660 9639
rect 26608 9596 26660 9605
rect 24676 9460 24728 9512
rect 25780 9460 25832 9512
rect 23204 9324 23256 9376
rect 23480 9324 23532 9376
rect 26056 9435 26108 9444
rect 26056 9401 26065 9435
rect 26065 9401 26099 9435
rect 26099 9401 26108 9435
rect 26976 9528 27028 9580
rect 29552 9596 29604 9648
rect 27436 9571 27488 9580
rect 27436 9537 27445 9571
rect 27445 9537 27479 9571
rect 27479 9537 27488 9571
rect 27436 9528 27488 9537
rect 26792 9460 26844 9512
rect 27620 9460 27672 9512
rect 28264 9460 28316 9512
rect 30932 9528 30984 9580
rect 34520 9707 34572 9716
rect 34520 9673 34529 9707
rect 34529 9673 34563 9707
rect 34563 9673 34572 9707
rect 34520 9664 34572 9673
rect 32680 9596 32732 9648
rect 33048 9639 33100 9648
rect 33048 9605 33057 9639
rect 33057 9605 33091 9639
rect 33091 9605 33100 9639
rect 33048 9596 33100 9605
rect 34428 9596 34480 9648
rect 35808 9664 35860 9716
rect 36728 9707 36780 9716
rect 36728 9673 36737 9707
rect 36737 9673 36771 9707
rect 36771 9673 36780 9707
rect 36728 9664 36780 9673
rect 26056 9392 26108 9401
rect 26332 9324 26384 9376
rect 27252 9367 27304 9376
rect 27252 9333 27261 9367
rect 27261 9333 27295 9367
rect 27295 9333 27304 9367
rect 27252 9324 27304 9333
rect 27712 9367 27764 9376
rect 27712 9333 27721 9367
rect 27721 9333 27755 9367
rect 27755 9333 27764 9367
rect 27712 9324 27764 9333
rect 30012 9324 30064 9376
rect 31576 9460 31628 9512
rect 32220 9571 32272 9580
rect 32220 9537 32229 9571
rect 32229 9537 32263 9571
rect 32263 9537 32272 9571
rect 32220 9528 32272 9537
rect 32496 9528 32548 9580
rect 35716 9571 35768 9580
rect 35716 9537 35725 9571
rect 35725 9537 35759 9571
rect 35759 9537 35768 9571
rect 35716 9528 35768 9537
rect 35900 9528 35952 9580
rect 37924 9596 37976 9648
rect 38016 9571 38068 9580
rect 38016 9537 38025 9571
rect 38025 9537 38059 9571
rect 38059 9537 38068 9571
rect 38016 9528 38068 9537
rect 38936 9571 38988 9580
rect 38936 9537 38945 9571
rect 38945 9537 38979 9571
rect 38979 9537 38988 9571
rect 38936 9528 38988 9537
rect 39120 9528 39172 9580
rect 43352 9707 43404 9716
rect 43352 9673 43361 9707
rect 43361 9673 43395 9707
rect 43395 9673 43404 9707
rect 43352 9664 43404 9673
rect 43904 9664 43956 9716
rect 46020 9664 46072 9716
rect 39304 9528 39356 9580
rect 39580 9571 39632 9580
rect 39580 9537 39589 9571
rect 39589 9537 39623 9571
rect 39623 9537 39632 9571
rect 39580 9528 39632 9537
rect 40592 9596 40644 9648
rect 34796 9392 34848 9444
rect 36084 9503 36136 9512
rect 36084 9469 36093 9503
rect 36093 9469 36127 9503
rect 36127 9469 36136 9503
rect 36084 9460 36136 9469
rect 38200 9503 38252 9512
rect 38200 9469 38209 9503
rect 38209 9469 38243 9503
rect 38243 9469 38252 9503
rect 38200 9460 38252 9469
rect 40132 9460 40184 9512
rect 33508 9324 33560 9376
rect 35532 9367 35584 9376
rect 35532 9333 35541 9367
rect 35541 9333 35575 9367
rect 35575 9333 35584 9367
rect 35532 9324 35584 9333
rect 39028 9367 39080 9376
rect 39028 9333 39037 9367
rect 39037 9333 39071 9367
rect 39071 9333 39080 9367
rect 39028 9324 39080 9333
rect 40040 9324 40092 9376
rect 41604 9528 41656 9580
rect 41696 9571 41748 9580
rect 41696 9537 41705 9571
rect 41705 9537 41739 9571
rect 41739 9537 41748 9571
rect 41696 9528 41748 9537
rect 45560 9596 45612 9648
rect 43904 9571 43956 9580
rect 41880 9460 41932 9512
rect 42156 9460 42208 9512
rect 43904 9537 43913 9571
rect 43913 9537 43947 9571
rect 43947 9537 43956 9571
rect 43904 9528 43956 9537
rect 44272 9503 44324 9512
rect 44272 9469 44281 9503
rect 44281 9469 44315 9503
rect 44315 9469 44324 9503
rect 44272 9460 44324 9469
rect 41512 9324 41564 9376
rect 41788 9324 41840 9376
rect 41880 9324 41932 9376
rect 43260 9324 43312 9376
rect 44456 9324 44508 9376
rect 45100 9571 45152 9580
rect 45100 9537 45109 9571
rect 45109 9537 45143 9571
rect 45143 9537 45152 9571
rect 45100 9528 45152 9537
rect 46756 9596 46808 9648
rect 50160 9664 50212 9716
rect 48964 9596 49016 9648
rect 46480 9571 46532 9580
rect 46480 9537 46489 9571
rect 46489 9537 46523 9571
rect 46523 9537 46532 9571
rect 46480 9528 46532 9537
rect 46572 9571 46624 9580
rect 46572 9537 46581 9571
rect 46581 9537 46615 9571
rect 46615 9537 46624 9571
rect 46572 9528 46624 9537
rect 47216 9571 47268 9580
rect 47216 9537 47225 9571
rect 47225 9537 47259 9571
rect 47259 9537 47268 9571
rect 47216 9528 47268 9537
rect 47860 9571 47912 9580
rect 47860 9537 47869 9571
rect 47869 9537 47903 9571
rect 47903 9537 47912 9571
rect 47860 9528 47912 9537
rect 47952 9571 48004 9580
rect 47952 9537 47961 9571
rect 47961 9537 47995 9571
rect 47995 9537 48004 9571
rect 47952 9528 48004 9537
rect 49240 9571 49292 9580
rect 49240 9537 49249 9571
rect 49249 9537 49283 9571
rect 49283 9537 49292 9571
rect 49240 9528 49292 9537
rect 51080 9571 51132 9580
rect 51080 9537 51089 9571
rect 51089 9537 51123 9571
rect 51123 9537 51132 9571
rect 51080 9528 51132 9537
rect 45652 9460 45704 9512
rect 45468 9392 45520 9444
rect 46756 9435 46808 9444
rect 46756 9401 46765 9435
rect 46765 9401 46799 9435
rect 46799 9401 46808 9435
rect 46756 9392 46808 9401
rect 48044 9460 48096 9512
rect 51448 9460 51500 9512
rect 45192 9324 45244 9376
rect 46664 9324 46716 9376
rect 47308 9367 47360 9376
rect 47308 9333 47317 9367
rect 47317 9333 47351 9367
rect 47351 9333 47360 9367
rect 47308 9324 47360 9333
rect 47676 9367 47728 9376
rect 47676 9333 47685 9367
rect 47685 9333 47719 9367
rect 47719 9333 47728 9367
rect 47676 9324 47728 9333
rect 49148 9324 49200 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 23572 9120 23624 9172
rect 24768 9120 24820 9172
rect 26056 9120 26108 9172
rect 26148 9163 26200 9172
rect 26148 9129 26157 9163
rect 26157 9129 26191 9163
rect 26191 9129 26200 9163
rect 26148 9120 26200 9129
rect 26608 9120 26660 9172
rect 26792 9163 26844 9172
rect 26792 9129 26801 9163
rect 26801 9129 26835 9163
rect 26835 9129 26844 9163
rect 26792 9120 26844 9129
rect 27252 9120 27304 9172
rect 27712 9120 27764 9172
rect 34428 9163 34480 9172
rect 34428 9129 34437 9163
rect 34437 9129 34471 9163
rect 34471 9129 34480 9163
rect 34428 9120 34480 9129
rect 34796 9120 34848 9172
rect 36084 9163 36136 9172
rect 36084 9129 36093 9163
rect 36093 9129 36127 9163
rect 36127 9129 36136 9163
rect 36084 9120 36136 9129
rect 39028 9120 39080 9172
rect 40684 9120 40736 9172
rect 24952 9027 25004 9036
rect 24952 8993 24961 9027
rect 24961 8993 24995 9027
rect 24995 8993 25004 9027
rect 24952 8984 25004 8993
rect 25596 8984 25648 9036
rect 23664 8848 23716 8900
rect 24400 8848 24452 8900
rect 24676 8848 24728 8900
rect 26516 8916 26568 8968
rect 26608 8823 26660 8832
rect 26608 8789 26617 8823
rect 26617 8789 26651 8823
rect 26651 8789 26660 8823
rect 26608 8780 26660 8789
rect 26700 8780 26752 8832
rect 35808 9052 35860 9104
rect 27620 8959 27672 8968
rect 27620 8925 27629 8959
rect 27629 8925 27663 8959
rect 27663 8925 27672 8959
rect 27620 8916 27672 8925
rect 30012 8916 30064 8968
rect 30380 8916 30432 8968
rect 31300 8916 31352 8968
rect 33600 8916 33652 8968
rect 35808 8916 35860 8968
rect 36452 9095 36504 9104
rect 36452 9061 36461 9095
rect 36461 9061 36495 9095
rect 36495 9061 36504 9095
rect 36452 9052 36504 9061
rect 39120 9052 39172 9104
rect 40132 8984 40184 9036
rect 41328 8984 41380 9036
rect 43260 9120 43312 9172
rect 47676 9120 47728 9172
rect 47860 9120 47912 9172
rect 48044 9120 48096 9172
rect 48228 9120 48280 9172
rect 49056 9120 49108 9172
rect 49148 9163 49200 9172
rect 49148 9129 49157 9163
rect 49157 9129 49191 9163
rect 49191 9129 49200 9163
rect 49148 9120 49200 9129
rect 34428 8848 34480 8900
rect 35348 8848 35400 8900
rect 35900 8848 35952 8900
rect 29368 8823 29420 8832
rect 29368 8789 29377 8823
rect 29377 8789 29411 8823
rect 29411 8789 29420 8823
rect 29368 8780 29420 8789
rect 32772 8823 32824 8832
rect 32772 8789 32781 8823
rect 32781 8789 32815 8823
rect 32815 8789 32824 8823
rect 32772 8780 32824 8789
rect 35716 8780 35768 8832
rect 37096 8916 37148 8968
rect 37372 8916 37424 8968
rect 37464 8959 37516 8968
rect 37464 8925 37473 8959
rect 37473 8925 37507 8959
rect 37507 8925 37516 8959
rect 37464 8916 37516 8925
rect 37832 8959 37884 8968
rect 37832 8925 37841 8959
rect 37841 8925 37875 8959
rect 37875 8925 37884 8959
rect 37832 8916 37884 8925
rect 44272 8984 44324 9036
rect 45652 8984 45704 9036
rect 47032 8984 47084 9036
rect 45100 8959 45152 8968
rect 45100 8925 45109 8959
rect 45109 8925 45143 8959
rect 45143 8925 45152 8959
rect 45100 8916 45152 8925
rect 45192 8916 45244 8968
rect 45560 8959 45612 8968
rect 45560 8925 45569 8959
rect 45569 8925 45603 8959
rect 45603 8925 45612 8959
rect 45560 8916 45612 8925
rect 38384 8848 38436 8900
rect 40684 8848 40736 8900
rect 37188 8780 37240 8832
rect 37372 8780 37424 8832
rect 39580 8780 39632 8832
rect 41972 8780 42024 8832
rect 42984 8848 43036 8900
rect 48596 8959 48648 8968
rect 48596 8925 48605 8959
rect 48605 8925 48639 8959
rect 48639 8925 48648 8959
rect 48596 8916 48648 8925
rect 48780 8959 48832 8968
rect 48780 8925 48789 8959
rect 48789 8925 48823 8959
rect 48823 8925 48832 8959
rect 48780 8916 48832 8925
rect 48872 8959 48924 8968
rect 48872 8925 48881 8959
rect 48881 8925 48915 8959
rect 48915 8925 48924 8959
rect 48872 8916 48924 8925
rect 48964 8959 49016 8968
rect 48964 8925 48973 8959
rect 48973 8925 49007 8959
rect 49007 8925 49016 8959
rect 48964 8916 49016 8925
rect 49792 8916 49844 8968
rect 46756 8848 46808 8900
rect 47308 8848 47360 8900
rect 49056 8848 49108 8900
rect 50068 8916 50120 8968
rect 68468 8959 68520 8968
rect 68468 8925 68477 8959
rect 68477 8925 68511 8959
rect 68511 8925 68520 8959
rect 68468 8916 68520 8925
rect 45376 8780 45428 8832
rect 48228 8780 48280 8832
rect 48964 8780 49016 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 23204 8576 23256 8628
rect 25596 8576 25648 8628
rect 26148 8576 26200 8628
rect 23480 8551 23532 8560
rect 23480 8517 23489 8551
rect 23489 8517 23523 8551
rect 23523 8517 23532 8551
rect 23480 8508 23532 8517
rect 24492 8508 24544 8560
rect 29368 8576 29420 8628
rect 32404 8576 32456 8628
rect 32772 8576 32824 8628
rect 33968 8576 34020 8628
rect 35532 8576 35584 8628
rect 37832 8576 37884 8628
rect 38384 8576 38436 8628
rect 40684 8619 40736 8628
rect 40684 8585 40693 8619
rect 40693 8585 40727 8619
rect 40727 8585 40736 8619
rect 40684 8576 40736 8585
rect 28080 8551 28132 8560
rect 28080 8517 28089 8551
rect 28089 8517 28123 8551
rect 28123 8517 28132 8551
rect 28080 8508 28132 8517
rect 26700 8483 26752 8492
rect 26700 8449 26709 8483
rect 26709 8449 26743 8483
rect 26743 8449 26752 8483
rect 26700 8440 26752 8449
rect 26976 8483 27028 8492
rect 26976 8449 26985 8483
rect 26985 8449 27019 8483
rect 27019 8449 27028 8483
rect 26976 8440 27028 8449
rect 24952 8347 25004 8356
rect 24952 8313 24961 8347
rect 24961 8313 24995 8347
rect 24995 8313 25004 8347
rect 24952 8304 25004 8313
rect 32772 8415 32824 8424
rect 32772 8381 32781 8415
rect 32781 8381 32815 8415
rect 32815 8381 32824 8415
rect 32772 8372 32824 8381
rect 34244 8372 34296 8424
rect 33232 8304 33284 8356
rect 34704 8483 34756 8492
rect 34704 8449 34738 8483
rect 34738 8449 34756 8483
rect 34704 8440 34756 8449
rect 34428 8415 34480 8424
rect 34428 8381 34437 8415
rect 34437 8381 34471 8415
rect 34471 8381 34480 8415
rect 34428 8372 34480 8381
rect 36268 8440 36320 8492
rect 36636 8483 36688 8492
rect 36636 8449 36645 8483
rect 36645 8449 36679 8483
rect 36679 8449 36688 8483
rect 36636 8440 36688 8449
rect 37556 8508 37608 8560
rect 37924 8440 37976 8492
rect 40776 8508 40828 8560
rect 41972 8551 42024 8560
rect 41972 8517 41981 8551
rect 41981 8517 42015 8551
rect 42015 8517 42024 8551
rect 41972 8508 42024 8517
rect 46940 8576 46992 8628
rect 47952 8576 48004 8628
rect 48596 8619 48648 8628
rect 48596 8585 48605 8619
rect 48605 8585 48639 8619
rect 48639 8585 48648 8619
rect 48596 8576 48648 8585
rect 48780 8619 48832 8628
rect 48780 8585 48789 8619
rect 48789 8585 48823 8619
rect 48823 8585 48832 8619
rect 48780 8576 48832 8585
rect 49332 8576 49384 8628
rect 38200 8440 38252 8492
rect 38660 8372 38712 8424
rect 39948 8372 40000 8424
rect 35808 8347 35860 8356
rect 35808 8313 35817 8347
rect 35817 8313 35851 8347
rect 35851 8313 35860 8347
rect 35808 8304 35860 8313
rect 26240 8279 26292 8288
rect 26240 8245 26249 8279
rect 26249 8245 26283 8279
rect 26283 8245 26292 8279
rect 26240 8236 26292 8245
rect 30748 8236 30800 8288
rect 33324 8279 33376 8288
rect 33324 8245 33333 8279
rect 33333 8245 33367 8279
rect 33367 8245 33376 8279
rect 33324 8236 33376 8245
rect 34796 8236 34848 8288
rect 36636 8279 36688 8288
rect 36636 8245 36645 8279
rect 36645 8245 36679 8279
rect 36679 8245 36688 8279
rect 36636 8236 36688 8245
rect 41880 8483 41932 8492
rect 41880 8449 41889 8483
rect 41889 8449 41923 8483
rect 41923 8449 41932 8483
rect 41880 8440 41932 8449
rect 42064 8483 42116 8492
rect 42064 8449 42073 8483
rect 42073 8449 42107 8483
rect 42107 8449 42116 8483
rect 42064 8440 42116 8449
rect 41328 8372 41380 8424
rect 46572 8508 46624 8560
rect 48044 8508 48096 8560
rect 42984 8440 43036 8492
rect 44732 8440 44784 8492
rect 45468 8440 45520 8492
rect 45744 8440 45796 8492
rect 46020 8483 46072 8492
rect 46020 8449 46029 8483
rect 46029 8449 46063 8483
rect 46063 8449 46072 8483
rect 46020 8440 46072 8449
rect 46204 8440 46256 8492
rect 46756 8440 46808 8492
rect 49700 8508 49752 8560
rect 48872 8483 48924 8492
rect 48872 8449 48881 8483
rect 48881 8449 48915 8483
rect 48915 8449 48924 8483
rect 48872 8440 48924 8449
rect 51448 8483 51500 8492
rect 51448 8449 51457 8483
rect 51457 8449 51491 8483
rect 51491 8449 51500 8483
rect 51448 8440 51500 8449
rect 47032 8372 47084 8424
rect 49792 8415 49844 8424
rect 49792 8381 49801 8415
rect 49801 8381 49835 8415
rect 49835 8381 49844 8415
rect 49792 8372 49844 8381
rect 45560 8304 45612 8356
rect 46020 8304 46072 8356
rect 44732 8236 44784 8288
rect 49332 8236 49384 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 24492 8075 24544 8084
rect 24492 8041 24501 8075
rect 24501 8041 24535 8075
rect 24535 8041 24544 8075
rect 24492 8032 24544 8041
rect 26976 8032 27028 8084
rect 32220 8032 32272 8084
rect 32772 8032 32824 8084
rect 34520 8032 34572 8084
rect 34704 8075 34756 8084
rect 34704 8041 34713 8075
rect 34713 8041 34747 8075
rect 34747 8041 34756 8075
rect 34704 8032 34756 8041
rect 36268 7964 36320 8016
rect 25596 7896 25648 7948
rect 27620 7939 27672 7948
rect 27620 7905 27629 7939
rect 27629 7905 27663 7939
rect 27663 7905 27672 7939
rect 27620 7896 27672 7905
rect 29920 7896 29972 7948
rect 30380 7939 30432 7948
rect 30380 7905 30389 7939
rect 30389 7905 30423 7939
rect 30423 7905 30432 7939
rect 30380 7896 30432 7905
rect 32772 7896 32824 7948
rect 37924 7896 37976 7948
rect 38568 7896 38620 7948
rect 940 7828 992 7880
rect 24400 7871 24452 7880
rect 24400 7837 24409 7871
rect 24409 7837 24443 7871
rect 24443 7837 24452 7871
rect 24400 7828 24452 7837
rect 29828 7871 29880 7880
rect 29828 7837 29837 7871
rect 29837 7837 29871 7871
rect 29871 7837 29880 7871
rect 29828 7828 29880 7837
rect 24768 7760 24820 7812
rect 26332 7760 26384 7812
rect 27896 7803 27948 7812
rect 27896 7769 27905 7803
rect 27905 7769 27939 7803
rect 27939 7769 27948 7803
rect 27896 7760 27948 7769
rect 29276 7760 29328 7812
rect 31944 7828 31996 7880
rect 34428 7828 34480 7880
rect 34520 7828 34572 7880
rect 34796 7828 34848 7880
rect 30380 7760 30432 7812
rect 30748 7760 30800 7812
rect 31668 7760 31720 7812
rect 33324 7760 33376 7812
rect 35256 7871 35308 7880
rect 35256 7837 35265 7871
rect 35265 7837 35299 7871
rect 35299 7837 35308 7871
rect 35256 7828 35308 7837
rect 36636 7871 36688 7880
rect 36636 7837 36670 7871
rect 36670 7837 36688 7871
rect 36636 7828 36688 7837
rect 26240 7692 26292 7744
rect 29552 7692 29604 7744
rect 30012 7692 30064 7744
rect 33416 7692 33468 7744
rect 35900 7692 35952 7744
rect 35992 7735 36044 7744
rect 35992 7701 36001 7735
rect 36001 7701 36035 7735
rect 36035 7701 36044 7735
rect 35992 7692 36044 7701
rect 45744 8032 45796 8084
rect 45836 8075 45888 8084
rect 45836 8041 45845 8075
rect 45845 8041 45879 8075
rect 45879 8041 45888 8075
rect 45836 8032 45888 8041
rect 46112 7964 46164 8016
rect 41788 7828 41840 7880
rect 42156 7828 42208 7880
rect 42432 7871 42484 7880
rect 42432 7837 42441 7871
rect 42441 7837 42475 7871
rect 42475 7837 42484 7871
rect 42432 7828 42484 7837
rect 43536 7871 43588 7880
rect 43536 7837 43545 7871
rect 43545 7837 43579 7871
rect 43579 7837 43588 7871
rect 43536 7828 43588 7837
rect 46388 7871 46440 7880
rect 46388 7837 46397 7871
rect 46397 7837 46431 7871
rect 46431 7837 46440 7871
rect 46388 7828 46440 7837
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 41144 7735 41196 7744
rect 41144 7701 41153 7735
rect 41153 7701 41187 7735
rect 41187 7701 41196 7735
rect 41144 7692 41196 7701
rect 41420 7760 41472 7812
rect 46204 7760 46256 7812
rect 46664 7828 46716 7880
rect 47952 8032 48004 8084
rect 49792 8032 49844 8084
rect 47768 7939 47820 7948
rect 47768 7905 47777 7939
rect 47777 7905 47811 7939
rect 47811 7905 47820 7939
rect 47768 7896 47820 7905
rect 47676 7828 47728 7880
rect 49332 7939 49384 7948
rect 49332 7905 49341 7939
rect 49341 7905 49375 7939
rect 49375 7905 49384 7939
rect 49332 7896 49384 7905
rect 42064 7692 42116 7744
rect 42800 7692 42852 7744
rect 46020 7735 46072 7744
rect 46020 7701 46029 7735
rect 46029 7701 46063 7735
rect 46063 7701 46072 7735
rect 46020 7692 46072 7701
rect 48412 7803 48464 7812
rect 48412 7769 48437 7803
rect 48437 7769 48464 7803
rect 48412 7760 48464 7769
rect 47768 7692 47820 7744
rect 48136 7692 48188 7744
rect 48320 7692 48372 7744
rect 49516 7760 49568 7812
rect 48596 7735 48648 7744
rect 48596 7701 48605 7735
rect 48605 7701 48639 7735
rect 48639 7701 48648 7735
rect 48596 7692 48648 7701
rect 49148 7735 49200 7744
rect 49148 7701 49157 7735
rect 49157 7701 49191 7735
rect 49191 7701 49200 7735
rect 49148 7692 49200 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 26332 7531 26384 7540
rect 26332 7497 26341 7531
rect 26341 7497 26375 7531
rect 26375 7497 26384 7531
rect 26332 7488 26384 7497
rect 27896 7488 27948 7540
rect 29276 7531 29328 7540
rect 29276 7497 29285 7531
rect 29285 7497 29319 7531
rect 29319 7497 29328 7531
rect 29276 7488 29328 7497
rect 24768 7420 24820 7472
rect 29000 7352 29052 7404
rect 29552 7420 29604 7472
rect 31116 7420 31168 7472
rect 28540 7327 28592 7336
rect 28540 7293 28549 7327
rect 28549 7293 28583 7327
rect 28583 7293 28592 7327
rect 28540 7284 28592 7293
rect 28632 7284 28684 7336
rect 28816 7284 28868 7336
rect 28448 7216 28500 7268
rect 30104 7352 30156 7404
rect 31668 7488 31720 7540
rect 31944 7531 31996 7540
rect 31944 7497 31953 7531
rect 31953 7497 31987 7531
rect 31987 7497 31996 7531
rect 31944 7488 31996 7497
rect 30380 7216 30432 7268
rect 28632 7148 28684 7200
rect 29920 7148 29972 7200
rect 31576 7352 31628 7404
rect 31668 7352 31720 7404
rect 32404 7420 32456 7472
rect 33416 7531 33468 7540
rect 33416 7497 33425 7531
rect 33425 7497 33459 7531
rect 33459 7497 33468 7531
rect 33416 7488 33468 7497
rect 33692 7488 33744 7540
rect 35992 7488 36044 7540
rect 39396 7488 39448 7540
rect 34428 7352 34480 7404
rect 32220 7327 32272 7336
rect 32220 7293 32229 7327
rect 32229 7293 32263 7327
rect 32263 7293 32272 7327
rect 32220 7284 32272 7293
rect 32772 7284 32824 7336
rect 33232 7284 33284 7336
rect 34244 7284 34296 7336
rect 37464 7352 37516 7404
rect 40040 7395 40092 7404
rect 40040 7361 40049 7395
rect 40049 7361 40083 7395
rect 40083 7361 40092 7395
rect 40040 7352 40092 7361
rect 40132 7352 40184 7404
rect 41328 7420 41380 7472
rect 42432 7488 42484 7540
rect 43536 7488 43588 7540
rect 46020 7488 46072 7540
rect 45928 7463 45980 7472
rect 45928 7429 45937 7463
rect 45937 7429 45971 7463
rect 45971 7429 45980 7463
rect 45928 7420 45980 7429
rect 41144 7395 41196 7404
rect 41144 7361 41178 7395
rect 41178 7361 41196 7395
rect 41144 7352 41196 7361
rect 42432 7395 42484 7404
rect 42432 7361 42441 7395
rect 42441 7361 42475 7395
rect 42475 7361 42484 7395
rect 42432 7352 42484 7361
rect 42524 7352 42576 7404
rect 47676 7488 47728 7540
rect 48320 7488 48372 7540
rect 48412 7488 48464 7540
rect 48596 7488 48648 7540
rect 49148 7488 49200 7540
rect 48136 7463 48188 7472
rect 48136 7429 48145 7463
rect 48145 7429 48179 7463
rect 48179 7429 48188 7463
rect 48136 7420 48188 7429
rect 46756 7352 46808 7404
rect 48044 7352 48096 7404
rect 49516 7420 49568 7472
rect 47768 7284 47820 7336
rect 49700 7352 49752 7404
rect 49792 7216 49844 7268
rect 32864 7148 32916 7200
rect 33968 7148 34020 7200
rect 36268 7191 36320 7200
rect 36268 7157 36277 7191
rect 36277 7157 36311 7191
rect 36311 7157 36320 7191
rect 36268 7148 36320 7157
rect 37004 7191 37056 7200
rect 37004 7157 37013 7191
rect 37013 7157 37047 7191
rect 37047 7157 37056 7191
rect 37004 7148 37056 7157
rect 39948 7191 40000 7200
rect 39948 7157 39957 7191
rect 39957 7157 39991 7191
rect 39991 7157 40000 7191
rect 39948 7148 40000 7157
rect 46112 7191 46164 7200
rect 46112 7157 46121 7191
rect 46121 7157 46155 7191
rect 46155 7157 46164 7191
rect 46112 7148 46164 7157
rect 46480 7191 46532 7200
rect 46480 7157 46489 7191
rect 46489 7157 46523 7191
rect 46523 7157 46532 7191
rect 46480 7148 46532 7157
rect 46664 7191 46716 7200
rect 46664 7157 46673 7191
rect 46673 7157 46707 7191
rect 46707 7157 46716 7191
rect 46664 7148 46716 7157
rect 46848 7148 46900 7200
rect 49056 7191 49108 7200
rect 49056 7157 49065 7191
rect 49065 7157 49099 7191
rect 49099 7157 49108 7191
rect 49056 7148 49108 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 29552 6944 29604 6996
rect 35900 6944 35952 6996
rect 37924 6944 37976 6996
rect 39120 6944 39172 6996
rect 42524 6944 42576 6996
rect 28540 6876 28592 6928
rect 33416 6876 33468 6928
rect 33508 6876 33560 6928
rect 27896 6851 27948 6860
rect 25596 6783 25648 6792
rect 25596 6749 25605 6783
rect 25605 6749 25639 6783
rect 25639 6749 25648 6783
rect 25596 6740 25648 6749
rect 27896 6817 27905 6851
rect 27905 6817 27939 6851
rect 27939 6817 27948 6851
rect 27896 6808 27948 6817
rect 28908 6808 28960 6860
rect 28448 6740 28500 6792
rect 28816 6783 28868 6792
rect 28816 6749 28825 6783
rect 28825 6749 28859 6783
rect 28859 6749 28868 6783
rect 28816 6740 28868 6749
rect 26608 6672 26660 6724
rect 27436 6715 27488 6724
rect 27436 6681 27445 6715
rect 27445 6681 27479 6715
rect 27479 6681 27488 6715
rect 27436 6672 27488 6681
rect 27528 6647 27580 6656
rect 27528 6613 27543 6647
rect 27543 6613 27577 6647
rect 27577 6613 27580 6647
rect 27528 6604 27580 6613
rect 28908 6715 28960 6724
rect 28908 6681 28917 6715
rect 28917 6681 28951 6715
rect 28951 6681 28960 6715
rect 28908 6672 28960 6681
rect 32220 6808 32272 6860
rect 31760 6783 31812 6792
rect 31760 6749 31769 6783
rect 31769 6749 31803 6783
rect 31803 6749 31812 6783
rect 31760 6740 31812 6749
rect 32496 6740 32548 6792
rect 34244 6808 34296 6860
rect 34060 6740 34112 6792
rect 36084 6740 36136 6792
rect 37004 6740 37056 6792
rect 37188 6740 37240 6792
rect 37464 6783 37516 6792
rect 33232 6672 33284 6724
rect 37464 6749 37473 6783
rect 37473 6749 37507 6783
rect 37507 6749 37516 6783
rect 37464 6740 37516 6749
rect 39580 6876 39632 6928
rect 38200 6740 38252 6792
rect 39580 6740 39632 6792
rect 39948 6783 40000 6792
rect 39948 6749 39957 6783
rect 39957 6749 39991 6783
rect 39991 6749 40000 6783
rect 39948 6740 40000 6749
rect 42064 6876 42116 6928
rect 42432 6808 42484 6860
rect 45928 6944 45980 6996
rect 42156 6783 42208 6792
rect 42156 6749 42165 6783
rect 42165 6749 42199 6783
rect 42199 6749 42208 6783
rect 42156 6740 42208 6749
rect 42800 6740 42852 6792
rect 46480 6876 46532 6928
rect 49056 6944 49108 6996
rect 49792 6987 49844 6996
rect 49792 6953 49801 6987
rect 49801 6953 49835 6987
rect 49835 6953 49844 6987
rect 49792 6944 49844 6953
rect 29736 6604 29788 6656
rect 30104 6647 30156 6656
rect 30104 6613 30113 6647
rect 30113 6613 30147 6647
rect 30147 6613 30156 6647
rect 30104 6604 30156 6613
rect 30840 6604 30892 6656
rect 32588 6604 32640 6656
rect 33692 6647 33744 6656
rect 33692 6613 33701 6647
rect 33701 6613 33735 6647
rect 33735 6613 33744 6647
rect 33692 6604 33744 6613
rect 33784 6604 33836 6656
rect 34520 6604 34572 6656
rect 34704 6647 34756 6656
rect 34704 6613 34713 6647
rect 34713 6613 34747 6647
rect 34747 6613 34756 6647
rect 34704 6604 34756 6613
rect 35624 6604 35676 6656
rect 37280 6647 37332 6656
rect 37280 6613 37289 6647
rect 37289 6613 37323 6647
rect 37323 6613 37332 6647
rect 37280 6604 37332 6613
rect 38660 6604 38712 6656
rect 40224 6647 40276 6656
rect 40224 6613 40233 6647
rect 40233 6613 40267 6647
rect 40267 6613 40276 6647
rect 40224 6604 40276 6613
rect 44272 6672 44324 6724
rect 40592 6604 40644 6656
rect 45928 6740 45980 6792
rect 46112 6740 46164 6792
rect 46756 6783 46808 6792
rect 46756 6749 46765 6783
rect 46765 6749 46799 6783
rect 46799 6749 46808 6783
rect 46756 6740 46808 6749
rect 45376 6715 45428 6724
rect 45376 6681 45385 6715
rect 45385 6681 45419 6715
rect 45419 6681 45428 6715
rect 45376 6672 45428 6681
rect 46020 6672 46072 6724
rect 46204 6672 46256 6724
rect 47032 6740 47084 6792
rect 48780 6672 48832 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 26608 6400 26660 6452
rect 27528 6400 27580 6452
rect 28632 6400 28684 6452
rect 28816 6443 28868 6452
rect 28816 6409 28825 6443
rect 28825 6409 28859 6443
rect 28859 6409 28868 6443
rect 28816 6400 28868 6409
rect 29000 6400 29052 6452
rect 29828 6400 29880 6452
rect 30104 6400 30156 6452
rect 26976 6264 27028 6316
rect 27896 6264 27948 6316
rect 28356 6264 28408 6316
rect 28816 6264 28868 6316
rect 28448 6196 28500 6248
rect 28908 6196 28960 6248
rect 27988 6128 28040 6180
rect 28724 6128 28776 6180
rect 29552 6307 29604 6316
rect 29552 6273 29561 6307
rect 29561 6273 29595 6307
rect 29595 6273 29604 6307
rect 29552 6264 29604 6273
rect 29920 6307 29972 6316
rect 29920 6273 29929 6307
rect 29929 6273 29963 6307
rect 29963 6273 29972 6307
rect 29920 6264 29972 6273
rect 30012 6196 30064 6248
rect 30472 6307 30524 6316
rect 30472 6273 30481 6307
rect 30481 6273 30515 6307
rect 30515 6273 30524 6307
rect 30472 6264 30524 6273
rect 30564 6264 30616 6316
rect 30656 6307 30708 6316
rect 30656 6273 30665 6307
rect 30665 6273 30699 6307
rect 30699 6273 30708 6307
rect 30656 6264 30708 6273
rect 31760 6400 31812 6452
rect 31668 6332 31720 6384
rect 33784 6332 33836 6384
rect 36268 6332 36320 6384
rect 32772 6239 32824 6248
rect 32772 6205 32781 6239
rect 32781 6205 32815 6239
rect 32815 6205 32824 6239
rect 32772 6196 32824 6205
rect 33048 6239 33100 6248
rect 33048 6205 33057 6239
rect 33057 6205 33091 6239
rect 33091 6205 33100 6239
rect 33048 6196 33100 6205
rect 32496 6128 32548 6180
rect 30104 6060 30156 6112
rect 30288 6060 30340 6112
rect 31024 6103 31076 6112
rect 31024 6069 31033 6103
rect 31033 6069 31067 6103
rect 31067 6069 31076 6103
rect 31024 6060 31076 6069
rect 31576 6060 31628 6112
rect 34520 6103 34572 6112
rect 34520 6069 34529 6103
rect 34529 6069 34563 6103
rect 34563 6069 34572 6103
rect 34520 6060 34572 6069
rect 35808 6307 35860 6316
rect 35808 6273 35817 6307
rect 35817 6273 35851 6307
rect 35851 6273 35860 6307
rect 35808 6264 35860 6273
rect 36360 6307 36412 6316
rect 36360 6273 36369 6307
rect 36369 6273 36403 6307
rect 36403 6273 36412 6307
rect 36360 6264 36412 6273
rect 38844 6443 38896 6452
rect 38844 6409 38853 6443
rect 38853 6409 38887 6443
rect 38887 6409 38896 6443
rect 38844 6400 38896 6409
rect 39120 6443 39172 6452
rect 39120 6409 39129 6443
rect 39129 6409 39163 6443
rect 39163 6409 39172 6443
rect 39120 6400 39172 6409
rect 41512 6400 41564 6452
rect 44272 6443 44324 6452
rect 44272 6409 44281 6443
rect 44281 6409 44315 6443
rect 44315 6409 44324 6443
rect 44272 6400 44324 6409
rect 38292 6332 38344 6384
rect 43904 6332 43956 6384
rect 36084 6239 36136 6248
rect 36084 6205 36093 6239
rect 36093 6205 36127 6239
rect 36127 6205 36136 6239
rect 36084 6196 36136 6205
rect 36176 6196 36228 6248
rect 37096 6264 37148 6316
rect 37372 6264 37424 6316
rect 38292 6196 38344 6248
rect 38936 6307 38988 6316
rect 38936 6273 38945 6307
rect 38945 6273 38979 6307
rect 38979 6273 38988 6307
rect 38936 6264 38988 6273
rect 39304 6264 39356 6316
rect 40408 6307 40460 6316
rect 40408 6273 40417 6307
rect 40417 6273 40451 6307
rect 40451 6273 40460 6307
rect 40408 6264 40460 6273
rect 40592 6307 40644 6316
rect 40592 6273 40601 6307
rect 40601 6273 40635 6307
rect 40635 6273 40644 6307
rect 40592 6264 40644 6273
rect 46112 6332 46164 6384
rect 46204 6332 46256 6384
rect 48780 6443 48832 6452
rect 48780 6409 48789 6443
rect 48789 6409 48823 6443
rect 48823 6409 48832 6443
rect 48780 6400 48832 6409
rect 46664 6332 46716 6384
rect 41236 6239 41288 6248
rect 41236 6205 41245 6239
rect 41245 6205 41279 6239
rect 41279 6205 41288 6239
rect 41236 6196 41288 6205
rect 41420 6239 41472 6248
rect 41420 6205 41429 6239
rect 41429 6205 41463 6239
rect 41463 6205 41472 6239
rect 41420 6196 41472 6205
rect 45836 6196 45888 6248
rect 46572 6307 46624 6316
rect 46572 6273 46581 6307
rect 46581 6273 46615 6307
rect 46615 6273 46624 6307
rect 46572 6264 46624 6273
rect 46756 6196 46808 6248
rect 46020 6128 46072 6180
rect 46572 6128 46624 6180
rect 47952 6264 48004 6316
rect 48320 6264 48372 6316
rect 68468 6171 68520 6180
rect 68468 6137 68477 6171
rect 68477 6137 68511 6171
rect 68511 6137 68520 6171
rect 68468 6128 68520 6137
rect 37004 6103 37056 6112
rect 37004 6069 37013 6103
rect 37013 6069 37047 6103
rect 37047 6069 37056 6103
rect 37004 6060 37056 6069
rect 37832 6103 37884 6112
rect 37832 6069 37841 6103
rect 37841 6069 37875 6103
rect 37875 6069 37884 6103
rect 37832 6060 37884 6069
rect 38568 6103 38620 6112
rect 38568 6069 38577 6103
rect 38577 6069 38611 6103
rect 38611 6069 38620 6103
rect 38568 6060 38620 6069
rect 40868 6060 40920 6112
rect 46204 6103 46256 6112
rect 46204 6069 46213 6103
rect 46213 6069 46247 6103
rect 46247 6069 46256 6103
rect 46204 6060 46256 6069
rect 47400 6060 47452 6112
rect 48872 6060 48924 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 27436 5856 27488 5908
rect 29552 5856 29604 5908
rect 30288 5856 30340 5908
rect 30380 5899 30432 5908
rect 30380 5865 30389 5899
rect 30389 5865 30423 5899
rect 30423 5865 30432 5899
rect 30380 5856 30432 5865
rect 27988 5720 28040 5772
rect 28080 5695 28132 5704
rect 28080 5661 28089 5695
rect 28089 5661 28123 5695
rect 28123 5661 28132 5695
rect 28080 5652 28132 5661
rect 29920 5763 29972 5772
rect 29920 5729 29929 5763
rect 29929 5729 29963 5763
rect 29963 5729 29972 5763
rect 29920 5720 29972 5729
rect 30564 5763 30616 5772
rect 30564 5729 30573 5763
rect 30573 5729 30607 5763
rect 30607 5729 30616 5763
rect 30564 5720 30616 5729
rect 30748 5763 30800 5772
rect 30748 5729 30757 5763
rect 30757 5729 30791 5763
rect 30791 5729 30800 5763
rect 30748 5720 30800 5729
rect 31944 5856 31996 5908
rect 31668 5720 31720 5772
rect 33048 5899 33100 5908
rect 33048 5865 33057 5899
rect 33057 5865 33091 5899
rect 33091 5865 33100 5899
rect 33048 5856 33100 5865
rect 33692 5856 33744 5908
rect 36176 5899 36228 5908
rect 36176 5865 36185 5899
rect 36185 5865 36219 5899
rect 36219 5865 36228 5899
rect 36176 5856 36228 5865
rect 37004 5856 37056 5908
rect 37280 5899 37332 5908
rect 37280 5865 37289 5899
rect 37289 5865 37323 5899
rect 37323 5865 37332 5899
rect 37280 5856 37332 5865
rect 37464 5856 37516 5908
rect 25596 5584 25648 5636
rect 25688 5627 25740 5636
rect 25688 5593 25697 5627
rect 25697 5593 25731 5627
rect 25731 5593 25740 5627
rect 25688 5584 25740 5593
rect 26424 5584 26476 5636
rect 27252 5559 27304 5568
rect 27252 5525 27261 5559
rect 27261 5525 27295 5559
rect 27295 5525 27304 5559
rect 27252 5516 27304 5525
rect 27712 5559 27764 5568
rect 27712 5525 27721 5559
rect 27721 5525 27755 5559
rect 27755 5525 27764 5559
rect 27712 5516 27764 5525
rect 28540 5695 28592 5704
rect 28540 5661 28549 5695
rect 28549 5661 28583 5695
rect 28583 5661 28592 5695
rect 28540 5652 28592 5661
rect 28632 5652 28684 5704
rect 29828 5695 29880 5704
rect 29828 5661 29837 5695
rect 29837 5661 29871 5695
rect 29871 5661 29880 5695
rect 29828 5652 29880 5661
rect 30012 5652 30064 5704
rect 30104 5652 30156 5704
rect 30380 5652 30432 5704
rect 30840 5695 30892 5704
rect 30840 5661 30849 5695
rect 30849 5661 30883 5695
rect 30883 5661 30892 5695
rect 30840 5652 30892 5661
rect 31576 5695 31628 5704
rect 28448 5516 28500 5568
rect 28816 5516 28868 5568
rect 31208 5584 31260 5636
rect 31576 5661 31585 5695
rect 31585 5661 31619 5695
rect 31619 5661 31628 5695
rect 31576 5652 31628 5661
rect 31944 5652 31996 5704
rect 32312 5695 32364 5704
rect 32312 5661 32321 5695
rect 32321 5661 32355 5695
rect 32355 5661 32364 5695
rect 32312 5652 32364 5661
rect 32496 5695 32548 5704
rect 32496 5661 32505 5695
rect 32505 5661 32539 5695
rect 32539 5661 32548 5695
rect 32496 5652 32548 5661
rect 32588 5695 32640 5704
rect 32588 5661 32623 5695
rect 32623 5661 32640 5695
rect 32588 5652 32640 5661
rect 33140 5652 33192 5704
rect 33416 5652 33468 5704
rect 34520 5652 34572 5704
rect 37096 5788 37148 5840
rect 37740 5720 37792 5772
rect 37832 5720 37884 5772
rect 38568 5856 38620 5908
rect 38936 5856 38988 5908
rect 40500 5856 40552 5908
rect 40868 5856 40920 5908
rect 46204 5856 46256 5908
rect 46388 5899 46440 5908
rect 46388 5865 46397 5899
rect 46397 5865 46431 5899
rect 46431 5865 46440 5899
rect 46388 5856 46440 5865
rect 46756 5899 46808 5908
rect 46756 5865 46765 5899
rect 46765 5865 46799 5899
rect 46799 5865 46808 5899
rect 48872 5899 48924 5908
rect 46756 5856 46808 5865
rect 48872 5865 48881 5899
rect 48881 5865 48915 5899
rect 48915 5865 48924 5899
rect 48872 5856 48924 5865
rect 38200 5652 38252 5704
rect 41236 5788 41288 5840
rect 46112 5788 46164 5840
rect 31484 5559 31536 5568
rect 31484 5525 31493 5559
rect 31493 5525 31527 5559
rect 31527 5525 31536 5559
rect 31484 5516 31536 5525
rect 31576 5516 31628 5568
rect 32128 5559 32180 5568
rect 32128 5525 32137 5559
rect 32137 5525 32171 5559
rect 32171 5525 32180 5559
rect 32128 5516 32180 5525
rect 36176 5516 36228 5568
rect 36452 5559 36504 5568
rect 36452 5525 36461 5559
rect 36461 5525 36495 5559
rect 36495 5525 36504 5559
rect 36452 5516 36504 5525
rect 36820 5516 36872 5568
rect 37188 5516 37240 5568
rect 39396 5695 39448 5704
rect 39396 5661 39405 5695
rect 39405 5661 39439 5695
rect 39439 5661 39448 5695
rect 39396 5652 39448 5661
rect 40408 5720 40460 5772
rect 41328 5720 41380 5772
rect 45836 5720 45888 5772
rect 40224 5695 40276 5704
rect 40224 5661 40233 5695
rect 40233 5661 40267 5695
rect 40267 5661 40276 5695
rect 40224 5652 40276 5661
rect 43904 5652 43956 5704
rect 46296 5720 46348 5772
rect 46940 5720 46992 5772
rect 47400 5763 47452 5772
rect 47400 5729 47409 5763
rect 47409 5729 47443 5763
rect 47443 5729 47452 5763
rect 47400 5720 47452 5729
rect 47032 5652 47084 5704
rect 48412 5652 48464 5704
rect 39212 5516 39264 5568
rect 39304 5516 39356 5568
rect 39672 5516 39724 5568
rect 40684 5584 40736 5636
rect 41144 5627 41196 5636
rect 41144 5593 41153 5627
rect 41153 5593 41187 5627
rect 41187 5593 41196 5627
rect 41144 5584 41196 5593
rect 40960 5559 41012 5568
rect 40960 5525 40969 5559
rect 40969 5525 41003 5559
rect 41003 5525 41012 5559
rect 40960 5516 41012 5525
rect 41972 5627 42024 5636
rect 41972 5593 41981 5627
rect 41981 5593 42015 5627
rect 42015 5593 42024 5627
rect 41972 5584 42024 5593
rect 41420 5516 41472 5568
rect 46848 5516 46900 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 25688 5312 25740 5364
rect 26424 5312 26476 5364
rect 27252 5312 27304 5364
rect 28356 5312 28408 5364
rect 28448 5312 28500 5364
rect 29000 5312 29052 5364
rect 29460 5355 29512 5364
rect 29460 5321 29469 5355
rect 29469 5321 29503 5355
rect 29503 5321 29512 5355
rect 29460 5312 29512 5321
rect 29828 5312 29880 5364
rect 30656 5312 30708 5364
rect 31668 5312 31720 5364
rect 31944 5355 31996 5364
rect 31944 5321 31953 5355
rect 31953 5321 31987 5355
rect 31987 5321 31996 5355
rect 31944 5312 31996 5321
rect 32312 5312 32364 5364
rect 33140 5312 33192 5364
rect 39120 5312 39172 5364
rect 40500 5312 40552 5364
rect 40684 5355 40736 5364
rect 40684 5321 40693 5355
rect 40693 5321 40727 5355
rect 40727 5321 40736 5355
rect 40684 5312 40736 5321
rect 41972 5312 42024 5364
rect 45376 5312 45428 5364
rect 46480 5312 46532 5364
rect 46848 5312 46900 5364
rect 26976 5176 27028 5228
rect 27712 5176 27764 5228
rect 28632 5244 28684 5296
rect 28724 5219 28776 5228
rect 28724 5185 28733 5219
rect 28733 5185 28767 5219
rect 28767 5185 28776 5219
rect 28724 5176 28776 5185
rect 28816 5219 28868 5228
rect 28816 5185 28825 5219
rect 28825 5185 28859 5219
rect 28859 5185 28868 5219
rect 28816 5176 28868 5185
rect 30932 5244 30984 5296
rect 31024 5176 31076 5228
rect 31484 5176 31536 5228
rect 27620 5151 27672 5160
rect 27620 5117 27629 5151
rect 27629 5117 27663 5151
rect 27663 5117 27672 5151
rect 27620 5108 27672 5117
rect 28080 5108 28132 5160
rect 30380 5108 30432 5160
rect 31208 5108 31260 5160
rect 32128 5219 32180 5228
rect 32128 5185 32137 5219
rect 32137 5185 32171 5219
rect 32171 5185 32180 5219
rect 32128 5176 32180 5185
rect 35440 5244 35492 5296
rect 36452 5287 36504 5296
rect 36452 5253 36461 5287
rect 36461 5253 36495 5287
rect 36495 5253 36504 5287
rect 36452 5244 36504 5253
rect 35992 5176 36044 5228
rect 36268 5219 36320 5228
rect 36268 5185 36277 5219
rect 36277 5185 36311 5219
rect 36311 5185 36320 5219
rect 36268 5176 36320 5185
rect 39488 5219 39540 5228
rect 39488 5185 39497 5219
rect 39497 5185 39531 5219
rect 39531 5185 39540 5219
rect 39488 5176 39540 5185
rect 39580 5176 39632 5228
rect 44456 5244 44508 5296
rect 46020 5244 46072 5296
rect 33876 5108 33928 5160
rect 36084 5108 36136 5160
rect 36176 5151 36228 5160
rect 36176 5117 36185 5151
rect 36185 5117 36219 5151
rect 36219 5117 36228 5151
rect 36176 5108 36228 5117
rect 36728 5108 36780 5160
rect 40960 5219 41012 5228
rect 40960 5185 40969 5219
rect 40969 5185 41003 5219
rect 41003 5185 41012 5219
rect 40960 5176 41012 5185
rect 41236 5219 41288 5228
rect 41236 5185 41245 5219
rect 41245 5185 41279 5219
rect 41279 5185 41288 5219
rect 41236 5176 41288 5185
rect 41512 5219 41564 5228
rect 41512 5185 41521 5219
rect 41521 5185 41555 5219
rect 41555 5185 41564 5219
rect 41512 5176 41564 5185
rect 41144 5108 41196 5160
rect 42432 5151 42484 5160
rect 42432 5117 42441 5151
rect 42441 5117 42475 5151
rect 42475 5117 42484 5151
rect 42432 5108 42484 5117
rect 36544 5040 36596 5092
rect 27068 5015 27120 5024
rect 27068 4981 27077 5015
rect 27077 4981 27111 5015
rect 27111 4981 27120 5015
rect 27068 4972 27120 4981
rect 29460 4972 29512 5024
rect 30656 4972 30708 5024
rect 32496 4972 32548 5024
rect 33048 4972 33100 5024
rect 33600 4972 33652 5024
rect 36636 5015 36688 5024
rect 36636 4981 36645 5015
rect 36645 4981 36679 5015
rect 36679 4981 36688 5015
rect 36636 4972 36688 4981
rect 37188 4972 37240 5024
rect 39672 5015 39724 5024
rect 39672 4981 39681 5015
rect 39681 4981 39715 5015
rect 39715 4981 39724 5015
rect 39672 4972 39724 4981
rect 40316 4972 40368 5024
rect 40776 5015 40828 5024
rect 40776 4981 40785 5015
rect 40785 4981 40819 5015
rect 40819 4981 40828 5015
rect 40776 4972 40828 4981
rect 43720 5151 43772 5160
rect 43720 5117 43729 5151
rect 43729 5117 43763 5151
rect 43763 5117 43772 5151
rect 43720 5108 43772 5117
rect 46112 5108 46164 5160
rect 45100 4972 45152 5024
rect 45284 5015 45336 5024
rect 45284 4981 45293 5015
rect 45293 4981 45327 5015
rect 45327 4981 45336 5015
rect 45284 4972 45336 4981
rect 45928 4972 45980 5024
rect 46480 5219 46532 5228
rect 46480 5185 46489 5219
rect 46489 5185 46523 5219
rect 46523 5185 46532 5219
rect 46480 5176 46532 5185
rect 46572 5219 46624 5228
rect 46572 5185 46607 5219
rect 46607 5185 46624 5219
rect 46572 5176 46624 5185
rect 46848 5219 46900 5228
rect 46848 5185 46857 5219
rect 46857 5185 46891 5219
rect 46891 5185 46900 5219
rect 46848 5176 46900 5185
rect 46940 5176 46992 5228
rect 47584 5219 47636 5228
rect 47584 5185 47593 5219
rect 47593 5185 47627 5219
rect 47627 5185 47636 5219
rect 47584 5176 47636 5185
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 27068 4768 27120 4820
rect 27620 4768 27672 4820
rect 28540 4768 28592 4820
rect 30472 4768 30524 4820
rect 32496 4768 32548 4820
rect 33600 4811 33652 4820
rect 33600 4777 33609 4811
rect 33609 4777 33643 4811
rect 33643 4777 33652 4811
rect 33600 4768 33652 4777
rect 35440 4768 35492 4820
rect 36084 4811 36136 4820
rect 36084 4777 36093 4811
rect 36093 4777 36127 4811
rect 36127 4777 36136 4811
rect 36084 4768 36136 4777
rect 37464 4768 37516 4820
rect 28908 4700 28960 4752
rect 34060 4700 34112 4752
rect 36268 4700 36320 4752
rect 25596 4632 25648 4684
rect 31852 4675 31904 4684
rect 31852 4641 31861 4675
rect 31861 4641 31895 4675
rect 31895 4641 31904 4675
rect 31852 4632 31904 4641
rect 32772 4632 32824 4684
rect 33876 4632 33928 4684
rect 27436 4564 27488 4616
rect 30656 4564 30708 4616
rect 30932 4607 30984 4616
rect 30932 4573 30941 4607
rect 30941 4573 30975 4607
rect 30975 4573 30984 4607
rect 30932 4564 30984 4573
rect 27068 4496 27120 4548
rect 27988 4539 28040 4548
rect 27988 4505 27997 4539
rect 27997 4505 28031 4539
rect 28031 4505 28040 4539
rect 27988 4496 28040 4505
rect 30564 4496 30616 4548
rect 34612 4564 34664 4616
rect 35992 4607 36044 4616
rect 35992 4573 36001 4607
rect 36001 4573 36035 4607
rect 36035 4573 36044 4607
rect 35992 4564 36044 4573
rect 39488 4811 39540 4820
rect 39488 4777 39497 4811
rect 39497 4777 39531 4811
rect 39531 4777 39540 4811
rect 39488 4768 39540 4777
rect 40776 4768 40828 4820
rect 42432 4768 42484 4820
rect 43720 4768 43772 4820
rect 44456 4811 44508 4820
rect 44456 4777 44465 4811
rect 44465 4777 44499 4811
rect 44499 4777 44508 4811
rect 44456 4768 44508 4777
rect 45284 4768 45336 4820
rect 45928 4768 45980 4820
rect 38384 4700 38436 4752
rect 39396 4700 39448 4752
rect 36544 4607 36596 4616
rect 36544 4573 36579 4607
rect 36579 4573 36596 4607
rect 36544 4564 36596 4573
rect 36728 4607 36780 4616
rect 36728 4573 36737 4607
rect 36737 4573 36771 4607
rect 36771 4573 36780 4607
rect 36728 4564 36780 4573
rect 36820 4607 36872 4616
rect 36820 4573 36829 4607
rect 36829 4573 36863 4607
rect 36863 4573 36872 4607
rect 36820 4564 36872 4573
rect 31392 4496 31444 4548
rect 33140 4496 33192 4548
rect 29000 4428 29052 4480
rect 35992 4471 36044 4480
rect 35992 4437 36001 4471
rect 36001 4437 36035 4471
rect 36035 4437 36044 4471
rect 35992 4428 36044 4437
rect 37556 4539 37608 4548
rect 37556 4505 37565 4539
rect 37565 4505 37599 4539
rect 37599 4505 37608 4539
rect 37556 4496 37608 4505
rect 38200 4607 38252 4616
rect 38200 4573 38209 4607
rect 38209 4573 38243 4607
rect 38243 4573 38252 4607
rect 38200 4564 38252 4573
rect 38660 4564 38712 4616
rect 39580 4632 39632 4684
rect 45100 4632 45152 4684
rect 47032 4632 47084 4684
rect 37464 4471 37516 4480
rect 37464 4437 37473 4471
rect 37473 4437 37507 4471
rect 37507 4437 37516 4471
rect 37464 4428 37516 4437
rect 40040 4539 40092 4548
rect 40040 4505 40049 4539
rect 40049 4505 40083 4539
rect 40083 4505 40092 4539
rect 40040 4496 40092 4505
rect 40132 4539 40184 4548
rect 40132 4505 40141 4539
rect 40141 4505 40175 4539
rect 40175 4505 40184 4539
rect 40132 4496 40184 4505
rect 40500 4564 40552 4616
rect 43904 4564 43956 4616
rect 41328 4496 41380 4548
rect 47584 4607 47636 4616
rect 47584 4573 47593 4607
rect 47593 4573 47627 4607
rect 47627 4573 47636 4607
rect 47584 4564 47636 4573
rect 38200 4428 38252 4480
rect 39028 4428 39080 4480
rect 40224 4428 40276 4480
rect 40408 4471 40460 4480
rect 40408 4437 40417 4471
rect 40417 4437 40451 4471
rect 40451 4437 40460 4471
rect 40408 4428 40460 4437
rect 48320 4564 48372 4616
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 27068 4267 27120 4276
rect 27068 4233 27077 4267
rect 27077 4233 27111 4267
rect 27111 4233 27120 4267
rect 27068 4224 27120 4233
rect 28632 4224 28684 4276
rect 28356 4156 28408 4208
rect 26976 4131 27028 4140
rect 26976 4097 26985 4131
rect 26985 4097 27019 4131
rect 27019 4097 27028 4131
rect 26976 4088 27028 4097
rect 28356 4020 28408 4072
rect 28724 4156 28776 4208
rect 31668 4224 31720 4276
rect 35992 4224 36044 4276
rect 29092 4088 29144 4140
rect 29552 4088 29604 4140
rect 30104 4131 30156 4140
rect 30104 4097 30113 4131
rect 30113 4097 30147 4131
rect 30147 4097 30156 4131
rect 30104 4088 30156 4097
rect 31576 4156 31628 4208
rect 34796 4156 34848 4208
rect 32128 4088 32180 4140
rect 33324 4088 33376 4140
rect 33876 4131 33928 4140
rect 33876 4097 33885 4131
rect 33885 4097 33919 4131
rect 33919 4097 33928 4131
rect 33876 4088 33928 4097
rect 36636 4224 36688 4276
rect 36728 4224 36780 4276
rect 38200 4224 38252 4276
rect 38384 4224 38436 4276
rect 38476 4267 38528 4276
rect 38476 4233 38485 4267
rect 38485 4233 38519 4267
rect 38519 4233 38528 4267
rect 38476 4224 38528 4233
rect 38614 4224 38666 4276
rect 39028 4224 39080 4276
rect 39396 4224 39448 4276
rect 40224 4224 40276 4276
rect 36452 4156 36504 4208
rect 36268 4131 36320 4140
rect 36268 4097 36277 4131
rect 36277 4097 36311 4131
rect 36311 4097 36320 4131
rect 36268 4088 36320 4097
rect 37464 4088 37516 4140
rect 37740 4131 37792 4140
rect 37740 4097 37749 4131
rect 37749 4097 37783 4131
rect 37783 4097 37792 4131
rect 37740 4088 37792 4097
rect 28908 3952 28960 4004
rect 28724 3927 28776 3936
rect 28724 3893 28733 3927
rect 28733 3893 28767 3927
rect 28767 3893 28776 3927
rect 28724 3884 28776 3893
rect 29828 3927 29880 3936
rect 29828 3893 29837 3927
rect 29837 3893 29871 3927
rect 29871 3893 29880 3927
rect 29828 3884 29880 3893
rect 30656 4020 30708 4072
rect 33140 4020 33192 4072
rect 37188 4020 37240 4072
rect 36820 3952 36872 4004
rect 38384 4131 38436 4140
rect 38384 4097 38393 4131
rect 38393 4097 38427 4131
rect 38427 4097 38436 4131
rect 38384 4088 38436 4097
rect 40132 4156 40184 4208
rect 40316 4156 40368 4208
rect 39396 4131 39448 4140
rect 39396 4097 39405 4131
rect 39405 4097 39439 4131
rect 39439 4097 39448 4131
rect 39396 4088 39448 4097
rect 40500 4199 40552 4208
rect 40500 4165 40509 4199
rect 40509 4165 40543 4199
rect 40543 4165 40552 4199
rect 40500 4156 40552 4165
rect 30472 3884 30524 3936
rect 36544 3884 36596 3936
rect 38108 3952 38160 4004
rect 38292 3952 38344 4004
rect 39212 4020 39264 4072
rect 39948 4063 40000 4072
rect 39948 4029 39957 4063
rect 39957 4029 39991 4063
rect 39991 4029 40000 4063
rect 39948 4020 40000 4029
rect 40592 4020 40644 4072
rect 37556 3927 37608 3936
rect 37556 3893 37565 3927
rect 37565 3893 37599 3927
rect 37599 3893 37608 3927
rect 37556 3884 37608 3893
rect 38568 3884 38620 3936
rect 40040 3884 40092 3936
rect 41420 3884 41472 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 28724 3680 28776 3732
rect 28908 3680 28960 3732
rect 30104 3723 30156 3732
rect 30104 3689 30113 3723
rect 30113 3689 30147 3723
rect 30147 3689 30156 3723
rect 30104 3680 30156 3689
rect 30748 3723 30800 3732
rect 30748 3689 30757 3723
rect 30757 3689 30791 3723
rect 30791 3689 30800 3723
rect 30748 3680 30800 3689
rect 28632 3544 28684 3596
rect 34796 3723 34848 3732
rect 34796 3689 34805 3723
rect 34805 3689 34839 3723
rect 34839 3689 34848 3723
rect 34796 3680 34848 3689
rect 37740 3680 37792 3732
rect 39396 3680 39448 3732
rect 39948 3680 40000 3732
rect 38384 3612 38436 3664
rect 41420 3612 41472 3664
rect 31852 3544 31904 3596
rect 37372 3544 37424 3596
rect 38292 3544 38344 3596
rect 40040 3587 40092 3596
rect 40040 3553 40049 3587
rect 40049 3553 40083 3587
rect 40083 3553 40092 3587
rect 40040 3544 40092 3553
rect 41328 3544 41380 3596
rect 27804 3340 27856 3392
rect 30472 3519 30524 3528
rect 30472 3485 30481 3519
rect 30481 3485 30515 3519
rect 30515 3485 30524 3519
rect 30472 3476 30524 3485
rect 34612 3476 34664 3528
rect 36268 3519 36320 3528
rect 36268 3485 36277 3519
rect 36277 3485 36311 3519
rect 36311 3485 36320 3519
rect 36268 3476 36320 3485
rect 36820 3476 36872 3528
rect 29092 3408 29144 3460
rect 30656 3408 30708 3460
rect 31392 3408 31444 3460
rect 32312 3408 32364 3460
rect 33048 3451 33100 3460
rect 33048 3417 33057 3451
rect 33057 3417 33091 3451
rect 33091 3417 33100 3451
rect 33048 3408 33100 3417
rect 36544 3408 36596 3460
rect 29000 3340 29052 3392
rect 35900 3383 35952 3392
rect 35900 3349 35909 3383
rect 35909 3349 35943 3383
rect 35943 3349 35952 3383
rect 35900 3340 35952 3349
rect 38200 3408 38252 3460
rect 39304 3476 39356 3528
rect 68468 3519 68520 3528
rect 68468 3485 68477 3519
rect 68477 3485 68511 3519
rect 68511 3485 68520 3519
rect 68468 3476 68520 3485
rect 40408 3408 40460 3460
rect 39396 3340 39448 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 27436 3136 27488 3188
rect 27804 3068 27856 3120
rect 28448 3068 28500 3120
rect 29828 3136 29880 3188
rect 30472 3136 30524 3188
rect 31576 3179 31628 3188
rect 31576 3145 31585 3179
rect 31585 3145 31619 3179
rect 31619 3145 31628 3179
rect 31576 3136 31628 3145
rect 31668 3179 31720 3188
rect 31668 3145 31677 3179
rect 31677 3145 31711 3179
rect 31711 3145 31720 3179
rect 31668 3136 31720 3145
rect 32312 3136 32364 3188
rect 32864 3136 32916 3188
rect 34704 3136 34756 3188
rect 30380 3068 30432 3120
rect 32128 3043 32180 3052
rect 32128 3009 32137 3043
rect 32137 3009 32171 3043
rect 32171 3009 32180 3043
rect 32128 3000 32180 3009
rect 36360 3068 36412 3120
rect 37372 3136 37424 3188
rect 38292 3136 38344 3188
rect 37648 3068 37700 3120
rect 38660 3000 38712 3052
rect 39028 3000 39080 3052
rect 30656 2932 30708 2984
rect 31392 2932 31444 2984
rect 33048 2932 33100 2984
rect 33876 2932 33928 2984
rect 29092 2864 29144 2916
rect 31852 2864 31904 2916
rect 22560 2796 22612 2848
rect 31116 2796 31168 2848
rect 35348 2975 35400 2984
rect 35348 2941 35357 2975
rect 35357 2941 35391 2975
rect 35391 2941 35400 2975
rect 35348 2932 35400 2941
rect 37556 2975 37608 2984
rect 37556 2941 37565 2975
rect 37565 2941 37599 2975
rect 37599 2941 37608 2975
rect 37556 2932 37608 2941
rect 37648 2932 37700 2984
rect 39304 3043 39356 3052
rect 39304 3009 39313 3043
rect 39313 3009 39347 3043
rect 39347 3009 39356 3043
rect 39304 3000 39356 3009
rect 40040 3068 40092 3120
rect 40684 3068 40736 3120
rect 39120 2839 39172 2848
rect 39120 2805 39129 2839
rect 39129 2805 39163 2839
rect 39163 2805 39172 2839
rect 39120 2796 39172 2805
rect 39948 2975 40000 2984
rect 39948 2941 39957 2975
rect 39957 2941 39991 2975
rect 39991 2941 40000 2975
rect 39948 2932 40000 2941
rect 48320 2796 48372 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 28448 2592 28500 2644
rect 30380 2635 30432 2644
rect 30380 2601 30389 2635
rect 30389 2601 30423 2635
rect 30423 2601 30432 2635
rect 30380 2592 30432 2601
rect 32128 2592 32180 2644
rect 34612 2592 34664 2644
rect 35348 2592 35400 2644
rect 36360 2592 36412 2644
rect 38660 2592 38712 2644
rect 39948 2592 40000 2644
rect 40684 2635 40736 2644
rect 40684 2601 40693 2635
rect 40693 2601 40727 2635
rect 40727 2601 40736 2635
rect 40684 2592 40736 2601
rect 20 2524 72 2576
rect 35808 2524 35860 2576
rect 940 2388 992 2440
rect 1952 2388 2004 2440
rect 4528 2388 4580 2440
rect 7104 2388 7156 2440
rect 9680 2388 9732 2440
rect 17408 2388 17460 2440
rect 25136 2388 25188 2440
rect 28356 2388 28408 2440
rect 30472 2388 30524 2440
rect 33140 2431 33192 2440
rect 33140 2397 33149 2431
rect 33149 2397 33183 2431
rect 33183 2397 33192 2431
rect 33140 2388 33192 2397
rect 35900 2388 35952 2440
rect 40592 2524 40644 2576
rect 38292 2388 38344 2440
rect 39672 2456 39724 2508
rect 39396 2431 39448 2440
rect 39396 2397 39405 2431
rect 39405 2397 39439 2431
rect 39439 2397 39448 2431
rect 39396 2388 39448 2397
rect 40132 2388 40184 2440
rect 43168 2388 43220 2440
rect 45744 2388 45796 2440
rect 48320 2388 48372 2440
rect 50896 2388 50948 2440
rect 53472 2388 53524 2440
rect 56048 2388 56100 2440
rect 58624 2388 58676 2440
rect 66352 2388 66404 2440
rect 68468 2431 68520 2440
rect 68468 2397 68477 2431
rect 68477 2397 68511 2431
rect 68511 2397 68520 2431
rect 68468 2388 68520 2397
rect 68652 2388 68704 2440
rect 31760 2320 31812 2372
rect 39212 2320 39264 2372
rect 12348 2252 12400 2304
rect 48320 2252 48372 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 18 69200 74 70000
rect 1950 69306 2006 70000
rect 4526 69306 4582 70000
rect 7102 69306 7158 70000
rect 9678 69306 9734 70000
rect 12254 69306 12310 70000
rect 14830 69306 14886 70000
rect 17406 69306 17462 70000
rect 19982 69306 20038 70000
rect 22558 69306 22614 70000
rect 25134 69306 25190 70000
rect 27710 69306 27766 70000
rect 1950 69278 2268 69306
rect 1950 69200 2006 69278
rect 938 67416 994 67425
rect 938 67351 994 67360
rect 952 67250 980 67351
rect 2240 67250 2268 69278
rect 4526 69278 4844 69306
rect 4526 69200 4582 69278
rect 4816 67250 4844 69278
rect 7102 69278 7420 69306
rect 7102 69200 7158 69278
rect 7392 67250 7420 69278
rect 9678 69278 9996 69306
rect 9678 69200 9734 69278
rect 9968 67250 9996 69278
rect 12254 69278 12388 69306
rect 12254 69200 12310 69278
rect 12360 67266 12388 69278
rect 14830 69278 15148 69306
rect 14830 69200 14886 69278
rect 12360 67250 12480 67266
rect 15120 67250 15148 69278
rect 17406 69278 17724 69306
rect 17406 69200 17462 69278
rect 17696 67250 17724 69278
rect 19982 69278 20300 69306
rect 19982 69200 20038 69278
rect 19574 67484 19882 67493
rect 19574 67482 19580 67484
rect 19636 67482 19660 67484
rect 19716 67482 19740 67484
rect 19796 67482 19820 67484
rect 19876 67482 19882 67484
rect 19636 67430 19638 67482
rect 19818 67430 19820 67482
rect 19574 67428 19580 67430
rect 19636 67428 19660 67430
rect 19716 67428 19740 67430
rect 19796 67428 19820 67430
rect 19876 67428 19882 67430
rect 19574 67419 19882 67428
rect 20272 67250 20300 69278
rect 22558 69278 22876 69306
rect 22558 69200 22614 69278
rect 22848 67250 22876 69278
rect 25134 69278 25452 69306
rect 25134 69200 25190 69278
rect 25424 67250 25452 69278
rect 27710 69278 28028 69306
rect 27710 69200 27766 69278
rect 28000 67250 28028 69278
rect 30286 69200 30342 70000
rect 32862 69306 32918 70000
rect 32862 69278 33088 69306
rect 32862 69200 32918 69278
rect 30300 67266 30328 69200
rect 33060 67538 33088 69278
rect 35438 69200 35494 70000
rect 38014 69306 38070 70000
rect 40590 69306 40646 70000
rect 38014 69278 38332 69306
rect 38014 69200 38070 69278
rect 33060 67510 33180 67538
rect 30300 67250 30420 67266
rect 33152 67250 33180 67510
rect 38304 67250 38332 69278
rect 40590 69278 40908 69306
rect 40590 69200 40646 69278
rect 40880 67250 40908 69278
rect 43166 69200 43222 70000
rect 45742 69306 45798 70000
rect 45742 69278 46060 69306
rect 45742 69200 45798 69278
rect 46032 67250 46060 69278
rect 48318 69200 48374 70000
rect 50894 69200 50950 70000
rect 53470 69306 53526 70000
rect 56046 69306 56102 70000
rect 58622 69306 58678 70000
rect 61198 69306 61254 70000
rect 63774 69306 63830 70000
rect 53470 69278 53788 69306
rect 53470 69200 53526 69278
rect 50294 67484 50602 67493
rect 50294 67482 50300 67484
rect 50356 67482 50380 67484
rect 50436 67482 50460 67484
rect 50516 67482 50540 67484
rect 50596 67482 50602 67484
rect 50356 67430 50358 67482
rect 50538 67430 50540 67482
rect 50294 67428 50300 67430
rect 50356 67428 50380 67430
rect 50436 67428 50460 67430
rect 50516 67428 50540 67430
rect 50596 67428 50602 67430
rect 50294 67419 50602 67428
rect 53760 67250 53788 69278
rect 56046 69278 56180 69306
rect 56046 69200 56102 69278
rect 56152 67386 56180 69278
rect 58622 69278 58940 69306
rect 58622 69200 58678 69278
rect 56140 67380 56192 67386
rect 56140 67322 56192 67328
rect 58912 67250 58940 69278
rect 61198 69278 61516 69306
rect 61198 69200 61254 69278
rect 61488 67250 61516 69278
rect 63774 69278 64092 69306
rect 63774 69200 63830 69278
rect 64064 67250 64092 69278
rect 66350 69200 66406 70000
rect 68926 69200 68982 70000
rect 68940 67250 68968 69200
rect 940 67244 992 67250
rect 940 67186 992 67192
rect 2228 67244 2280 67250
rect 2228 67186 2280 67192
rect 4804 67244 4856 67250
rect 4804 67186 4856 67192
rect 7380 67244 7432 67250
rect 7380 67186 7432 67192
rect 9956 67244 10008 67250
rect 12360 67244 12492 67250
rect 12360 67238 12440 67244
rect 9956 67186 10008 67192
rect 12440 67186 12492 67192
rect 15108 67244 15160 67250
rect 15108 67186 15160 67192
rect 17684 67244 17736 67250
rect 17684 67186 17736 67192
rect 20260 67244 20312 67250
rect 20260 67186 20312 67192
rect 22836 67244 22888 67250
rect 22836 67186 22888 67192
rect 25412 67244 25464 67250
rect 25412 67186 25464 67192
rect 27988 67244 28040 67250
rect 30300 67244 30432 67250
rect 30300 67238 30380 67244
rect 27988 67186 28040 67192
rect 30380 67186 30432 67192
rect 33140 67244 33192 67250
rect 33140 67186 33192 67192
rect 38292 67244 38344 67250
rect 38292 67186 38344 67192
rect 40868 67244 40920 67250
rect 40868 67186 40920 67192
rect 46020 67244 46072 67250
rect 46020 67186 46072 67192
rect 53748 67244 53800 67250
rect 53748 67186 53800 67192
rect 58900 67244 58952 67250
rect 58900 67186 58952 67192
rect 61476 67244 61528 67250
rect 61476 67186 61528 67192
rect 64052 67244 64104 67250
rect 64052 67186 64104 67192
rect 68928 67244 68980 67250
rect 68928 67186 68980 67192
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 19574 66396 19882 66405
rect 19574 66394 19580 66396
rect 19636 66394 19660 66396
rect 19716 66394 19740 66396
rect 19796 66394 19820 66396
rect 19876 66394 19882 66396
rect 19636 66342 19638 66394
rect 19818 66342 19820 66394
rect 19574 66340 19580 66342
rect 19636 66340 19660 66342
rect 19716 66340 19740 66342
rect 19796 66340 19820 66342
rect 19876 66340 19882 66342
rect 19574 66331 19882 66340
rect 50294 66396 50602 66405
rect 50294 66394 50300 66396
rect 50356 66394 50380 66396
rect 50436 66394 50460 66396
rect 50516 66394 50540 66396
rect 50596 66394 50602 66396
rect 50356 66342 50358 66394
rect 50538 66342 50540 66394
rect 50294 66340 50300 66342
rect 50356 66340 50380 66342
rect 50436 66340 50460 66342
rect 50516 66340 50540 66342
rect 50596 66340 50602 66342
rect 50294 66331 50602 66340
rect 68466 66056 68522 66065
rect 68466 65991 68468 66000
rect 68520 65991 68522 66000
rect 68468 65962 68520 65968
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 19574 65308 19882 65317
rect 19574 65306 19580 65308
rect 19636 65306 19660 65308
rect 19716 65306 19740 65308
rect 19796 65306 19820 65308
rect 19876 65306 19882 65308
rect 19636 65254 19638 65306
rect 19818 65254 19820 65306
rect 19574 65252 19580 65254
rect 19636 65252 19660 65254
rect 19716 65252 19740 65254
rect 19796 65252 19820 65254
rect 19876 65252 19882 65254
rect 19574 65243 19882 65252
rect 50294 65308 50602 65317
rect 50294 65306 50300 65308
rect 50356 65306 50380 65308
rect 50436 65306 50460 65308
rect 50516 65306 50540 65308
rect 50596 65306 50602 65308
rect 50356 65254 50358 65306
rect 50538 65254 50540 65306
rect 50294 65252 50300 65254
rect 50356 65252 50380 65254
rect 50436 65252 50460 65254
rect 50516 65252 50540 65254
rect 50596 65252 50602 65254
rect 50294 65243 50602 65252
rect 1584 64932 1636 64938
rect 1584 64874 1636 64880
rect 1596 64841 1624 64874
rect 1582 64832 1638 64841
rect 1582 64767 1638 64776
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 34934 64764 35242 64773
rect 34934 64762 34940 64764
rect 34996 64762 35020 64764
rect 35076 64762 35100 64764
rect 35156 64762 35180 64764
rect 35236 64762 35242 64764
rect 34996 64710 34998 64762
rect 35178 64710 35180 64762
rect 34934 64708 34940 64710
rect 34996 64708 35020 64710
rect 35076 64708 35100 64710
rect 35156 64708 35180 64710
rect 35236 64708 35242 64710
rect 34934 64699 35242 64708
rect 65654 64764 65962 64773
rect 65654 64762 65660 64764
rect 65716 64762 65740 64764
rect 65796 64762 65820 64764
rect 65876 64762 65900 64764
rect 65956 64762 65962 64764
rect 65716 64710 65718 64762
rect 65898 64710 65900 64762
rect 65654 64708 65660 64710
rect 65716 64708 65740 64710
rect 65796 64708 65820 64710
rect 65876 64708 65900 64710
rect 65956 64708 65962 64710
rect 65654 64699 65962 64708
rect 19574 64220 19882 64229
rect 19574 64218 19580 64220
rect 19636 64218 19660 64220
rect 19716 64218 19740 64220
rect 19796 64218 19820 64220
rect 19876 64218 19882 64220
rect 19636 64166 19638 64218
rect 19818 64166 19820 64218
rect 19574 64164 19580 64166
rect 19636 64164 19660 64166
rect 19716 64164 19740 64166
rect 19796 64164 19820 64166
rect 19876 64164 19882 64166
rect 19574 64155 19882 64164
rect 50294 64220 50602 64229
rect 50294 64218 50300 64220
rect 50356 64218 50380 64220
rect 50436 64218 50460 64220
rect 50516 64218 50540 64220
rect 50596 64218 50602 64220
rect 50356 64166 50358 64218
rect 50538 64166 50540 64218
rect 50294 64164 50300 64166
rect 50356 64164 50380 64166
rect 50436 64164 50460 64166
rect 50516 64164 50540 64166
rect 50596 64164 50602 64166
rect 50294 64155 50602 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 34934 63676 35242 63685
rect 34934 63674 34940 63676
rect 34996 63674 35020 63676
rect 35076 63674 35100 63676
rect 35156 63674 35180 63676
rect 35236 63674 35242 63676
rect 34996 63622 34998 63674
rect 35178 63622 35180 63674
rect 34934 63620 34940 63622
rect 34996 63620 35020 63622
rect 35076 63620 35100 63622
rect 35156 63620 35180 63622
rect 35236 63620 35242 63622
rect 34934 63611 35242 63620
rect 65654 63676 65962 63685
rect 65654 63674 65660 63676
rect 65716 63674 65740 63676
rect 65796 63674 65820 63676
rect 65876 63674 65900 63676
rect 65956 63674 65962 63676
rect 65716 63622 65718 63674
rect 65898 63622 65900 63674
rect 65654 63620 65660 63622
rect 65716 63620 65740 63622
rect 65796 63620 65820 63622
rect 65876 63620 65900 63622
rect 65956 63620 65962 63622
rect 65654 63611 65962 63620
rect 68468 63368 68520 63374
rect 68466 63336 68468 63345
rect 68520 63336 68522 63345
rect 68466 63271 68522 63280
rect 19574 63132 19882 63141
rect 19574 63130 19580 63132
rect 19636 63130 19660 63132
rect 19716 63130 19740 63132
rect 19796 63130 19820 63132
rect 19876 63130 19882 63132
rect 19636 63078 19638 63130
rect 19818 63078 19820 63130
rect 19574 63076 19580 63078
rect 19636 63076 19660 63078
rect 19716 63076 19740 63078
rect 19796 63076 19820 63078
rect 19876 63076 19882 63078
rect 19574 63067 19882 63076
rect 50294 63132 50602 63141
rect 50294 63130 50300 63132
rect 50356 63130 50380 63132
rect 50436 63130 50460 63132
rect 50516 63130 50540 63132
rect 50596 63130 50602 63132
rect 50356 63078 50358 63130
rect 50538 63078 50540 63130
rect 50294 63076 50300 63078
rect 50356 63076 50380 63078
rect 50436 63076 50460 63078
rect 50516 63076 50540 63078
rect 50596 63076 50602 63078
rect 50294 63067 50602 63076
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 34934 62588 35242 62597
rect 34934 62586 34940 62588
rect 34996 62586 35020 62588
rect 35076 62586 35100 62588
rect 35156 62586 35180 62588
rect 35236 62586 35242 62588
rect 34996 62534 34998 62586
rect 35178 62534 35180 62586
rect 34934 62532 34940 62534
rect 34996 62532 35020 62534
rect 35076 62532 35100 62534
rect 35156 62532 35180 62534
rect 35236 62532 35242 62534
rect 34934 62523 35242 62532
rect 65654 62588 65962 62597
rect 65654 62586 65660 62588
rect 65716 62586 65740 62588
rect 65796 62586 65820 62588
rect 65876 62586 65900 62588
rect 65956 62586 65962 62588
rect 65716 62534 65718 62586
rect 65898 62534 65900 62586
rect 65654 62532 65660 62534
rect 65716 62532 65740 62534
rect 65796 62532 65820 62534
rect 65876 62532 65900 62534
rect 65956 62532 65962 62534
rect 65654 62523 65962 62532
rect 19574 62044 19882 62053
rect 19574 62042 19580 62044
rect 19636 62042 19660 62044
rect 19716 62042 19740 62044
rect 19796 62042 19820 62044
rect 19876 62042 19882 62044
rect 19636 61990 19638 62042
rect 19818 61990 19820 62042
rect 19574 61988 19580 61990
rect 19636 61988 19660 61990
rect 19716 61988 19740 61990
rect 19796 61988 19820 61990
rect 19876 61988 19882 61990
rect 19574 61979 19882 61988
rect 50294 62044 50602 62053
rect 50294 62042 50300 62044
rect 50356 62042 50380 62044
rect 50436 62042 50460 62044
rect 50516 62042 50540 62044
rect 50596 62042 50602 62044
rect 50356 61990 50358 62042
rect 50538 61990 50540 62042
rect 50294 61988 50300 61990
rect 50356 61988 50380 61990
rect 50436 61988 50460 61990
rect 50516 61988 50540 61990
rect 50596 61988 50602 61990
rect 50294 61979 50602 61988
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 65654 61500 65962 61509
rect 65654 61498 65660 61500
rect 65716 61498 65740 61500
rect 65796 61498 65820 61500
rect 65876 61498 65900 61500
rect 65956 61498 65962 61500
rect 65716 61446 65718 61498
rect 65898 61446 65900 61498
rect 65654 61444 65660 61446
rect 65716 61444 65740 61446
rect 65796 61444 65820 61446
rect 65876 61444 65900 61446
rect 65956 61444 65962 61446
rect 65654 61435 65962 61444
rect 19574 60956 19882 60965
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60891 19882 60900
rect 50294 60956 50602 60965
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60891 50602 60900
rect 68192 60716 68244 60722
rect 68192 60658 68244 60664
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 65654 60412 65962 60421
rect 65654 60410 65660 60412
rect 65716 60410 65740 60412
rect 65796 60410 65820 60412
rect 65876 60410 65900 60412
rect 65956 60410 65962 60412
rect 65716 60358 65718 60410
rect 65898 60358 65900 60410
rect 65654 60356 65660 60358
rect 65716 60356 65740 60358
rect 65796 60356 65820 60358
rect 65876 60356 65900 60358
rect 65956 60356 65962 60358
rect 65654 60347 65962 60356
rect 19574 59868 19882 59877
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59803 19882 59812
rect 50294 59868 50602 59877
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59803 50602 59812
rect 1584 59424 1636 59430
rect 1584 59366 1636 59372
rect 1596 59265 1624 59366
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 1582 59256 1638 59265
rect 4214 59259 4522 59268
rect 34934 59324 35242 59333
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59259 35242 59268
rect 65654 59324 65962 59333
rect 65654 59322 65660 59324
rect 65716 59322 65740 59324
rect 65796 59322 65820 59324
rect 65876 59322 65900 59324
rect 65956 59322 65962 59324
rect 65716 59270 65718 59322
rect 65898 59270 65900 59322
rect 65654 59268 65660 59270
rect 65716 59268 65740 59270
rect 65796 59268 65820 59270
rect 65876 59268 65900 59270
rect 65956 59268 65962 59270
rect 65654 59259 65962 59268
rect 1582 59191 1638 59200
rect 19574 58780 19882 58789
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58715 19882 58724
rect 50294 58780 50602 58789
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58715 50602 58724
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 34934 58236 35242 58245
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58171 35242 58180
rect 65654 58236 65962 58245
rect 65654 58234 65660 58236
rect 65716 58234 65740 58236
rect 65796 58234 65820 58236
rect 65876 58234 65900 58236
rect 65956 58234 65962 58236
rect 65716 58182 65718 58234
rect 65898 58182 65900 58234
rect 65654 58180 65660 58182
rect 65716 58180 65740 58182
rect 65796 58180 65820 58182
rect 65876 58180 65900 58182
rect 65956 58180 65962 58182
rect 65654 58171 65962 58180
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 1584 56840 1636 56846
rect 1584 56782 1636 56788
rect 1596 56545 1624 56782
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 1582 56536 1638 56545
rect 19574 56539 19882 56548
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 1582 56471 1638 56480
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 65654 56060 65962 56069
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 940 51400 992 51406
rect 940 51342 992 51348
rect 952 51105 980 51342
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 938 51096 994 51105
rect 19574 51099 19882 51108
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 938 51031 994 51040
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 940 48544 992 48550
rect 940 48486 992 48492
rect 952 48385 980 48486
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 938 48376 994 48385
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 938 48311 994 48320
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 65654 46268 65962 46277
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 940 45960 992 45966
rect 940 45902 992 45908
rect 952 45665 980 45902
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 938 45656 994 45665
rect 19574 45659 19882 45668
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 938 45591 994 45600
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 65654 44092 65962 44101
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 940 43104 992 43110
rect 940 43046 992 43052
rect 952 42945 980 43046
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 938 42936 994 42945
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 938 42871 994 42880
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 65654 40828 65962 40837
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 940 37664 992 37670
rect 940 37606 992 37612
rect 952 37505 980 37606
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 938 37496 994 37505
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 938 37431 994 37440
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 940 35080 992 35086
rect 940 35022 992 35028
rect 952 34785 980 35022
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 938 34776 994 34785
rect 19574 34779 19882 34788
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 938 34711 994 34720
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 940 32224 992 32230
rect 940 32166 992 32172
rect 952 32065 980 32166
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 938 32056 994 32065
rect 4214 32059 4522 32068
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 938 31991 994 32000
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 940 29640 992 29646
rect 940 29582 992 29588
rect 952 29345 980 29582
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 938 29336 994 29345
rect 19574 29339 19882 29348
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 938 29271 994 29280
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 940 26784 992 26790
rect 940 26726 992 26732
rect 952 26625 980 26726
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 938 26616 994 26625
rect 4214 26619 4522 26628
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 938 26551 994 26560
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 31208 25288 31260 25294
rect 31208 25230 31260 25236
rect 28816 25152 28868 25158
rect 28816 25094 28868 25100
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 28828 24886 28856 25094
rect 28816 24880 28868 24886
rect 28816 24822 28868 24828
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 28920 24410 28948 25230
rect 29552 25220 29604 25226
rect 29552 25162 29604 25168
rect 29460 24608 29512 24614
rect 29460 24550 29512 24556
rect 28908 24404 28960 24410
rect 28908 24346 28960 24352
rect 29472 24290 29500 24550
rect 29564 24410 29592 25162
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 30288 24812 30340 24818
rect 30288 24754 30340 24760
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 29552 24404 29604 24410
rect 29552 24346 29604 24352
rect 29472 24262 29592 24290
rect 29564 24206 29592 24262
rect 940 24200 992 24206
rect 940 24142 992 24148
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 952 23905 980 24142
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 938 23896 994 23905
rect 19574 23899 19882 23908
rect 938 23831 994 23840
rect 29092 23792 29144 23798
rect 29092 23734 29144 23740
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 28448 23724 28500 23730
rect 28448 23666 28500 23672
rect 26976 23520 27028 23526
rect 26976 23462 27028 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 26608 23112 26660 23118
rect 26608 23054 26660 23060
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 26620 21622 26648 23054
rect 26988 23050 27016 23462
rect 26976 23044 27028 23050
rect 26976 22986 27028 22992
rect 27172 22778 27200 23666
rect 28080 23520 28132 23526
rect 28080 23462 28132 23468
rect 28092 22778 28120 23462
rect 28460 23322 28488 23666
rect 28908 23656 28960 23662
rect 28908 23598 28960 23604
rect 28448 23316 28500 23322
rect 28448 23258 28500 23264
rect 28920 23118 28948 23598
rect 29104 23118 29132 23734
rect 29472 23730 29500 24142
rect 29564 23798 29592 24142
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 29552 23792 29604 23798
rect 29552 23734 29604 23740
rect 29184 23724 29236 23730
rect 29184 23666 29236 23672
rect 29460 23724 29512 23730
rect 29460 23666 29512 23672
rect 29196 23186 29224 23666
rect 29472 23186 29500 23666
rect 29932 23186 29960 24006
rect 29184 23180 29236 23186
rect 29184 23122 29236 23128
rect 29460 23180 29512 23186
rect 29460 23122 29512 23128
rect 29920 23180 29972 23186
rect 29920 23122 29972 23128
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 29092 23112 29144 23118
rect 29092 23054 29144 23060
rect 28540 22976 28592 22982
rect 28540 22918 28592 22924
rect 29104 22930 29132 23054
rect 29276 22976 29328 22982
rect 29104 22924 29276 22930
rect 29104 22918 29328 22924
rect 27160 22772 27212 22778
rect 27160 22714 27212 22720
rect 28080 22772 28132 22778
rect 28080 22714 28132 22720
rect 26700 22568 26752 22574
rect 26700 22510 26752 22516
rect 26608 21616 26660 21622
rect 26608 21558 26660 21564
rect 940 21548 992 21554
rect 940 21490 992 21496
rect 952 21185 980 21490
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 952 18465 980 18702
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1780 17882 1808 21286
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 24964 20466 24992 21422
rect 26516 20868 26568 20874
rect 26516 20810 26568 20816
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 25792 20534 25820 20742
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 26528 20058 26556 20810
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26620 19786 26648 20402
rect 26712 19922 26740 22510
rect 28080 22024 28132 22030
rect 28080 21966 28132 21972
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27632 21554 27660 21830
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27620 21548 27672 21554
rect 27620 21490 27672 21496
rect 26884 21344 26936 21350
rect 26884 21286 26936 21292
rect 26896 20942 26924 21286
rect 27172 21146 27200 21490
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 27448 21010 27476 21490
rect 28092 21350 28120 21966
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 27436 21004 27488 21010
rect 27436 20946 27488 20952
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 27160 20936 27212 20942
rect 27160 20878 27212 20884
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 26804 20602 26832 20878
rect 26792 20596 26844 20602
rect 26792 20538 26844 20544
rect 27172 20398 27200 20878
rect 27160 20392 27212 20398
rect 27160 20334 27212 20340
rect 27620 20392 27672 20398
rect 27672 20340 27752 20346
rect 27620 20334 27752 20340
rect 27632 20318 27752 20334
rect 27620 20256 27672 20262
rect 27620 20198 27672 20204
rect 27632 20058 27660 20198
rect 27620 20052 27672 20058
rect 27620 19994 27672 20000
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 26252 18766 26280 19110
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 25240 17678 25268 18702
rect 26712 18426 26740 19858
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26988 19514 27016 19654
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 27172 18766 27200 19790
rect 27264 19360 27292 19790
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 27344 19372 27396 19378
rect 27264 19332 27344 19360
rect 27264 18970 27292 19332
rect 27344 19314 27396 19320
rect 27448 19174 27476 19654
rect 27436 19168 27488 19174
rect 27436 19110 27488 19116
rect 27540 19122 27568 19790
rect 27632 19242 27660 19790
rect 27724 19514 27752 20318
rect 27816 20058 27844 20878
rect 28092 20602 28120 21286
rect 28552 21078 28580 22918
rect 29104 22902 29316 22918
rect 29104 22234 29132 22902
rect 29092 22228 29144 22234
rect 29092 22170 29144 22176
rect 29092 22092 29144 22098
rect 29092 22034 29144 22040
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 28736 21146 28764 21490
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 28540 21072 28592 21078
rect 28540 21014 28592 21020
rect 28080 20596 28132 20602
rect 28080 20538 28132 20544
rect 28552 20466 28580 21014
rect 28828 20942 28856 21830
rect 29104 21690 29132 22034
rect 30024 22030 30052 24686
rect 30300 23866 30328 24754
rect 30564 24336 30616 24342
rect 30564 24278 30616 24284
rect 30576 24206 30604 24278
rect 30564 24200 30616 24206
rect 30564 24142 30616 24148
rect 30288 23860 30340 23866
rect 30288 23802 30340 23808
rect 30944 23662 30972 25094
rect 31220 24954 31248 25230
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 31208 24948 31260 24954
rect 31208 24890 31260 24896
rect 31668 24948 31720 24954
rect 31668 24890 31720 24896
rect 31220 24562 31248 24890
rect 31128 24534 31248 24562
rect 31024 24268 31076 24274
rect 31024 24210 31076 24216
rect 30932 23656 30984 23662
rect 30932 23598 30984 23604
rect 30196 23520 30248 23526
rect 30196 23462 30248 23468
rect 30208 23322 30236 23462
rect 31036 23322 31064 24210
rect 30196 23316 30248 23322
rect 30196 23258 30248 23264
rect 31024 23316 31076 23322
rect 31024 23258 31076 23264
rect 30208 22982 30236 23258
rect 31036 22982 31064 23258
rect 31128 23186 31156 24534
rect 31208 24404 31260 24410
rect 31208 24346 31260 24352
rect 31576 24404 31628 24410
rect 31576 24346 31628 24352
rect 31116 23180 31168 23186
rect 31116 23122 31168 23128
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 30380 22976 30432 22982
rect 30380 22918 30432 22924
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 30288 22772 30340 22778
rect 30288 22714 30340 22720
rect 30300 22094 30328 22714
rect 30116 22066 30328 22094
rect 30012 22024 30064 22030
rect 30012 21966 30064 21972
rect 29092 21684 29144 21690
rect 29092 21626 29144 21632
rect 28908 21616 28960 21622
rect 28908 21558 28960 21564
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28920 20466 28948 21558
rect 29104 21554 29132 21626
rect 30024 21622 30052 21966
rect 30116 21962 30144 22066
rect 30104 21956 30156 21962
rect 30104 21898 30156 21904
rect 30012 21616 30064 21622
rect 30012 21558 30064 21564
rect 29092 21548 29144 21554
rect 29092 21490 29144 21496
rect 29368 20868 29420 20874
rect 29368 20810 29420 20816
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 28080 20256 28132 20262
rect 28080 20198 28132 20204
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 27816 19718 27844 19994
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27804 19372 27856 19378
rect 27724 19332 27804 19360
rect 27620 19236 27672 19242
rect 27620 19178 27672 19184
rect 27724 19122 27752 19332
rect 27804 19314 27856 19320
rect 27540 19094 27752 19122
rect 27252 18964 27304 18970
rect 27252 18906 27304 18912
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 26700 18420 26752 18426
rect 26700 18362 26752 18368
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 25240 16590 25268 17614
rect 26608 17196 26660 17202
rect 26608 17138 26660 17144
rect 25780 16992 25832 16998
rect 25780 16934 25832 16940
rect 25792 16590 25820 16934
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 25240 15978 25268 16526
rect 26620 16250 26648 17138
rect 26712 16250 26740 18362
rect 27264 18290 27292 18906
rect 27540 18630 27568 19094
rect 28092 18970 28120 20198
rect 28632 19916 28684 19922
rect 28632 19858 28684 19864
rect 28644 19786 28672 19858
rect 28736 19854 28764 20402
rect 28920 19922 28948 20402
rect 28908 19916 28960 19922
rect 28908 19858 28960 19864
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 28448 19780 28500 19786
rect 28448 19722 28500 19728
rect 28632 19780 28684 19786
rect 28632 19722 28684 19728
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28080 18964 28132 18970
rect 28080 18906 28132 18912
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27264 17882 27292 18226
rect 28368 18154 28396 19110
rect 28460 18698 28488 19722
rect 28644 19378 28672 19722
rect 28736 19378 28764 19790
rect 29104 19514 29132 20402
rect 29092 19508 29144 19514
rect 29092 19450 29144 19456
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 28644 19242 28672 19314
rect 28908 19304 28960 19310
rect 28908 19246 28960 19252
rect 28632 19236 28684 19242
rect 28632 19178 28684 19184
rect 28448 18692 28500 18698
rect 28448 18634 28500 18640
rect 27804 18148 27856 18154
rect 27804 18090 27856 18096
rect 28356 18148 28408 18154
rect 28356 18090 28408 18096
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 27816 17746 27844 18090
rect 27988 18080 28040 18086
rect 27988 18022 28040 18028
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 28000 17678 28028 18022
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 26884 16448 26936 16454
rect 26884 16390 26936 16396
rect 26976 16448 27028 16454
rect 26976 16390 27028 16396
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26700 16244 26752 16250
rect 26700 16186 26752 16192
rect 26148 16176 26200 16182
rect 26200 16124 26372 16130
rect 26148 16118 26372 16124
rect 26056 16108 26108 16114
rect 26160 16102 26372 16118
rect 26056 16050 26108 16056
rect 25228 15972 25280 15978
rect 25228 15914 25280 15920
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 24860 15904 24912 15910
rect 24860 15846 24912 15852
rect 952 15745 980 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 938 15736 994 15745
rect 4214 15739 4522 15748
rect 938 15671 994 15680
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 24872 15026 24900 15846
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 25148 14822 25176 15438
rect 25240 14958 25268 15914
rect 26068 15706 26096 16050
rect 26148 16040 26200 16046
rect 26200 16000 26280 16028
rect 26148 15982 26200 15988
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 26252 15570 26280 16000
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26068 15162 26096 15438
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 22388 13326 22416 13806
rect 23216 13530 23244 13806
rect 23952 13530 23980 13942
rect 24872 13870 24900 14418
rect 25148 14414 25176 14758
rect 26068 14482 26096 15098
rect 26056 14476 26108 14482
rect 26056 14418 26108 14424
rect 26252 14414 26280 15302
rect 26344 14618 26372 16102
rect 26896 15586 26924 16390
rect 26988 16250 27016 16390
rect 27356 16250 27384 16390
rect 26976 16244 27028 16250
rect 26976 16186 27028 16192
rect 27344 16244 27396 16250
rect 27344 16186 27396 16192
rect 27540 16046 27568 17070
rect 27988 16584 28040 16590
rect 27988 16526 28040 16532
rect 28000 16250 28028 16526
rect 27988 16244 28040 16250
rect 27988 16186 28040 16192
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 26896 15558 27016 15586
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 26608 15360 26660 15366
rect 26608 15302 26660 15308
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 26620 14414 26648 15302
rect 26896 14618 26924 15438
rect 26988 15434 27016 15558
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 26976 15428 27028 15434
rect 26976 15370 27028 15376
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 26988 14414 27016 15370
rect 27068 15360 27120 15366
rect 27068 15302 27120 15308
rect 27080 15026 27108 15302
rect 27264 15026 27292 15506
rect 27356 15026 27384 15642
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 27632 15162 27660 15438
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 28092 15026 28120 15438
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 28080 15020 28132 15026
rect 28080 14962 28132 14968
rect 27356 14414 27384 14962
rect 27896 14816 27948 14822
rect 27896 14758 27948 14764
rect 25136 14408 25188 14414
rect 25136 14350 25188 14356
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 27344 14408 27396 14414
rect 27344 14350 27396 14356
rect 25964 14272 26016 14278
rect 25964 14214 26016 14220
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 952 13025 980 13262
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 938 13016 994 13025
rect 19574 13019 19882 13028
rect 938 12951 994 12960
rect 22388 12782 22416 13262
rect 23584 12986 23612 13262
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 22388 11218 22416 12718
rect 23676 12442 23704 12854
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23860 12238 23888 13262
rect 24872 13258 24900 13806
rect 24952 13456 25004 13462
rect 24952 13398 25004 13404
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24504 12442 24532 12718
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 24872 12170 24900 12786
rect 24964 12306 24992 13398
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 25320 13252 25372 13258
rect 25320 13194 25372 13200
rect 25780 13252 25832 13258
rect 25780 13194 25832 13200
rect 25056 12986 25084 13194
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25332 12782 25360 13194
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25320 12776 25372 12782
rect 25320 12718 25372 12724
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 25240 12238 25268 12718
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 24860 12164 24912 12170
rect 24860 12106 24912 12112
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 23584 10690 23612 12038
rect 24872 11642 24900 12106
rect 24780 11614 24900 11642
rect 24400 11212 24452 11218
rect 24400 11154 24452 11160
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 23676 10810 23704 11018
rect 24412 10810 24440 11154
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 23584 10674 23704 10690
rect 24780 10674 24808 11614
rect 25240 11558 25268 12174
rect 24860 11552 24912 11558
rect 24860 11494 24912 11500
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 24872 10810 24900 11494
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 23584 10668 23716 10674
rect 23584 10662 23664 10668
rect 23664 10610 23716 10616
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 952 10305 980 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 938 10296 994 10305
rect 4214 10299 4522 10308
rect 938 10231 994 10240
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 23492 9518 23520 9862
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 23216 8634 23244 9318
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23492 8566 23520 9318
rect 23584 9178 23612 9590
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23676 8906 23704 10610
rect 24780 9722 24808 10610
rect 25056 10606 25084 10950
rect 25148 10606 25176 11086
rect 25240 10742 25268 11494
rect 25332 11150 25360 12718
rect 25516 12714 25544 13126
rect 25504 12708 25556 12714
rect 25504 12650 25556 12656
rect 25516 11218 25544 12650
rect 25792 11898 25820 13194
rect 25976 12434 26004 14214
rect 27080 13394 27108 14350
rect 27908 14074 27936 14758
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 28368 13870 28396 17614
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 28356 13864 28408 13870
rect 28356 13806 28408 13812
rect 27804 13728 27856 13734
rect 27804 13670 27856 13676
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 26516 13252 26568 13258
rect 26516 13194 26568 13200
rect 26240 12640 26292 12646
rect 26240 12582 26292 12588
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 25976 12406 26096 12434
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25504 11212 25556 11218
rect 25504 11154 25556 11160
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25332 10810 25360 11086
rect 25516 11082 25544 11154
rect 25504 11076 25556 11082
rect 25504 11018 25556 11024
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24872 9586 24900 9930
rect 25240 9586 25268 10678
rect 25424 10538 25452 10950
rect 25516 10810 25544 11018
rect 25700 10810 25728 11698
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25792 11014 25820 11086
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25688 10804 25740 10810
rect 25688 10746 25740 10752
rect 25412 10532 25464 10538
rect 25412 10474 25464 10480
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25516 9994 25544 10406
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25608 9602 25636 9998
rect 25700 9926 25728 10746
rect 25884 10674 25912 11086
rect 25976 10742 26004 11154
rect 26068 11150 26096 12406
rect 26252 12306 26280 12582
rect 26344 12374 26372 12582
rect 26528 12442 26556 13194
rect 26700 13184 26752 13190
rect 26700 13126 26752 13132
rect 26712 12986 26740 13126
rect 26700 12980 26752 12986
rect 26700 12922 26752 12928
rect 26712 12646 26740 12922
rect 27080 12850 27108 13330
rect 27816 12850 27844 13670
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 26884 12708 26936 12714
rect 26884 12650 26936 12656
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26516 12436 26568 12442
rect 26516 12378 26568 12384
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26712 11830 26740 12582
rect 26896 11830 26924 12650
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27448 12238 27476 12582
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27436 12096 27488 12102
rect 27436 12038 27488 12044
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 26700 11824 26752 11830
rect 26528 11784 26700 11812
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26436 11558 26464 11698
rect 26424 11552 26476 11558
rect 26424 11494 26476 11500
rect 26436 11234 26464 11494
rect 26528 11354 26556 11784
rect 26884 11824 26936 11830
rect 26752 11784 26832 11812
rect 26700 11766 26752 11772
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26620 11354 26648 11494
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 26240 11212 26292 11218
rect 26436 11206 26556 11234
rect 26240 11154 26292 11160
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 26252 11014 26280 11154
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26240 11008 26292 11014
rect 26240 10950 26292 10956
rect 26436 10810 26464 11086
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 25964 10736 26016 10742
rect 25964 10678 26016 10684
rect 26056 10736 26108 10742
rect 26056 10678 26108 10684
rect 26332 10736 26384 10742
rect 26332 10678 26384 10684
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 25792 10554 25820 10610
rect 26068 10554 26096 10678
rect 25792 10526 26096 10554
rect 25792 10130 25820 10526
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 25688 9920 25740 9926
rect 25688 9862 25740 9868
rect 25700 9738 25728 9862
rect 25700 9710 25820 9738
rect 25792 9654 25820 9710
rect 26068 9654 26096 9998
rect 26148 9920 26200 9926
rect 26148 9862 26200 9868
rect 26160 9722 26188 9862
rect 26344 9722 26372 10678
rect 26436 10266 26464 10746
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26528 9926 26556 11206
rect 26804 11082 26832 11784
rect 26884 11766 26936 11772
rect 27172 11354 27200 11834
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27448 11150 27476 12038
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 28092 11354 28120 11698
rect 28080 11348 28132 11354
rect 28080 11290 28132 11296
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 28080 11144 28132 11150
rect 28080 11086 28132 11092
rect 26792 11076 26844 11082
rect 26792 11018 26844 11024
rect 27356 10810 27384 11086
rect 26792 10804 26844 10810
rect 26792 10746 26844 10752
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 26804 10198 26832 10746
rect 27528 10736 27580 10742
rect 27528 10678 27580 10684
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 27356 10266 27384 10542
rect 27344 10260 27396 10266
rect 27344 10202 27396 10208
rect 26792 10192 26844 10198
rect 26792 10134 26844 10140
rect 27540 10062 27568 10678
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 26516 9920 26568 9926
rect 26516 9862 26568 9868
rect 26148 9716 26200 9722
rect 26148 9658 26200 9664
rect 26332 9716 26384 9722
rect 26332 9658 26384 9664
rect 25688 9648 25740 9654
rect 25608 9596 25688 9602
rect 25608 9590 25740 9596
rect 25780 9648 25832 9654
rect 25780 9590 25832 9596
rect 26056 9648 26108 9654
rect 26056 9590 26108 9596
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25608 9574 25728 9590
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24688 8906 24716 9454
rect 24780 9178 24808 9522
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 25608 9042 25636 9574
rect 25792 9518 25820 9590
rect 25780 9512 25832 9518
rect 25780 9454 25832 9460
rect 26056 9444 26108 9450
rect 26056 9386 26108 9392
rect 26068 9178 26096 9386
rect 26344 9382 26372 9658
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24676 8900 24728 8906
rect 24676 8842 24728 8848
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 24412 7886 24440 8842
rect 24492 8560 24544 8566
rect 24492 8502 24544 8508
rect 24504 8090 24532 8502
rect 24964 8362 24992 8978
rect 26160 8634 26188 9114
rect 26528 8974 26556 9862
rect 26608 9648 26660 9654
rect 26608 9590 26660 9596
rect 26620 9178 26648 9590
rect 26792 9512 26844 9518
rect 26792 9454 26844 9460
rect 26804 9178 26832 9454
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 26792 9172 26844 9178
rect 26792 9114 26844 9120
rect 26516 8968 26568 8974
rect 26896 8922 26924 9998
rect 27436 9920 27488 9926
rect 27436 9862 27488 9868
rect 27448 9586 27476 9862
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 26516 8910 26568 8916
rect 26620 8894 26924 8922
rect 26620 8838 26648 8894
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24492 8084 24544 8090
rect 24492 8026 24544 8032
rect 25608 7954 25636 8570
rect 26712 8498 26740 8774
rect 26988 8498 27016 9522
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 27252 9376 27304 9382
rect 27252 9318 27304 9324
rect 27264 9178 27292 9318
rect 27252 9172 27304 9178
rect 27252 9114 27304 9120
rect 27632 8974 27660 9454
rect 27712 9376 27764 9382
rect 27712 9318 27764 9324
rect 27724 9178 27752 9318
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 26700 8492 26752 8498
rect 26700 8434 26752 8440
rect 26976 8492 27028 8498
rect 26976 8434 27028 8440
rect 26240 8288 26292 8294
rect 26240 8230 26292 8236
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 940 7880 992 7886
rect 940 7822 992 7828
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 952 7585 980 7822
rect 24768 7812 24820 7818
rect 24768 7754 24820 7760
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 938 7576 994 7585
rect 19574 7579 19882 7588
rect 938 7511 994 7520
rect 24780 7478 24808 7754
rect 24768 7472 24820 7478
rect 24768 7414 24820 7420
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 25608 6798 25636 7890
rect 26252 7750 26280 8230
rect 26988 8090 27016 8434
rect 26976 8084 27028 8090
rect 26976 8026 27028 8032
rect 27632 7954 27660 8910
rect 28092 8566 28120 11086
rect 28184 11014 28212 13806
rect 28356 11348 28408 11354
rect 28356 11290 28408 11296
rect 28368 11150 28396 11290
rect 28356 11144 28408 11150
rect 28356 11086 28408 11092
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 28184 10742 28212 10950
rect 28172 10736 28224 10742
rect 28172 10678 28224 10684
rect 28368 10470 28396 11086
rect 28460 10810 28488 18634
rect 28920 18630 28948 19246
rect 29184 18692 29236 18698
rect 29184 18634 29236 18640
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 29196 17270 29224 18634
rect 29276 17604 29328 17610
rect 29276 17546 29328 17552
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 28908 17128 28960 17134
rect 28736 17076 28908 17082
rect 28736 17070 28960 17076
rect 28736 17054 28948 17070
rect 28736 16794 28764 17054
rect 28816 16992 28868 16998
rect 28816 16934 28868 16940
rect 28828 16794 28856 16934
rect 28724 16788 28776 16794
rect 28724 16730 28776 16736
rect 28816 16788 28868 16794
rect 28816 16730 28868 16736
rect 29196 16658 29224 17206
rect 29184 16652 29236 16658
rect 29184 16594 29236 16600
rect 28724 16584 28776 16590
rect 28724 16526 28776 16532
rect 28632 16448 28684 16454
rect 28632 16390 28684 16396
rect 28540 15972 28592 15978
rect 28540 15914 28592 15920
rect 28552 15706 28580 15914
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28644 15570 28672 16390
rect 28736 15910 28764 16526
rect 28908 16516 28960 16522
rect 28908 16458 28960 16464
rect 28920 16402 28948 16458
rect 28920 16374 29040 16402
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28724 15904 28776 15910
rect 28724 15846 28776 15852
rect 28736 15570 28764 15846
rect 28828 15706 28856 16050
rect 28816 15700 28868 15706
rect 28816 15642 28868 15648
rect 28632 15564 28684 15570
rect 28632 15506 28684 15512
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 28724 15360 28776 15366
rect 28724 15302 28776 15308
rect 28736 15026 28764 15302
rect 28920 15162 28948 16186
rect 29012 16046 29040 16374
rect 29288 16114 29316 17546
rect 29380 17542 29408 20810
rect 30024 20398 30052 21558
rect 30392 21350 30420 22918
rect 31220 22778 31248 24346
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31300 24132 31352 24138
rect 31300 24074 31352 24080
rect 31312 23798 31340 24074
rect 31300 23792 31352 23798
rect 31300 23734 31352 23740
rect 31300 23044 31352 23050
rect 31300 22986 31352 22992
rect 31208 22772 31260 22778
rect 31208 22714 31260 22720
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30472 22432 30524 22438
rect 30472 22374 30524 22380
rect 30748 22432 30800 22438
rect 30748 22374 30800 22380
rect 30484 22030 30512 22374
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 30760 21690 30788 22374
rect 30852 22094 30880 22578
rect 31312 22574 31340 22986
rect 31300 22568 31352 22574
rect 31300 22510 31352 22516
rect 31404 22094 31432 24142
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 31496 23202 31524 24006
rect 31588 23798 31616 24346
rect 31576 23792 31628 23798
rect 31576 23734 31628 23740
rect 31680 23610 31708 24890
rect 34060 24880 34112 24886
rect 34060 24822 34112 24828
rect 31852 24812 31904 24818
rect 31852 24754 31904 24760
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 31864 24274 31892 24754
rect 31852 24268 31904 24274
rect 31852 24210 31904 24216
rect 31760 24064 31812 24070
rect 31760 24006 31812 24012
rect 31772 23730 31800 24006
rect 32220 23860 32272 23866
rect 32220 23802 32272 23808
rect 32232 23730 32260 23802
rect 31760 23724 31812 23730
rect 31760 23666 31812 23672
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32404 23724 32456 23730
rect 32404 23666 32456 23672
rect 31944 23656 31996 23662
rect 31680 23604 31944 23610
rect 31680 23598 31996 23604
rect 31680 23582 31984 23598
rect 31496 23186 31892 23202
rect 31496 23180 31904 23186
rect 31496 23174 31852 23180
rect 31852 23122 31904 23128
rect 31668 23112 31720 23118
rect 31668 23054 31720 23060
rect 32312 23112 32364 23118
rect 32416 23100 32444 23666
rect 32508 23118 32536 24754
rect 32956 23656 33008 23662
rect 32956 23598 33008 23604
rect 32680 23316 32732 23322
rect 32680 23258 32732 23264
rect 32968 23304 32996 23598
rect 33048 23316 33100 23322
rect 32968 23276 33048 23304
rect 32364 23072 32444 23100
rect 32312 23054 32364 23060
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 31496 22710 31524 22918
rect 31484 22704 31536 22710
rect 31484 22646 31536 22652
rect 31680 22574 31708 23054
rect 32036 23044 32088 23050
rect 32036 22986 32088 22992
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 32048 22574 32076 22986
rect 32140 22778 32168 22986
rect 32128 22772 32180 22778
rect 32128 22714 32180 22720
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31668 22568 31720 22574
rect 31668 22510 31720 22516
rect 32036 22568 32088 22574
rect 32036 22510 32088 22516
rect 31588 22234 31616 22510
rect 32416 22438 32444 23072
rect 32496 23112 32548 23118
rect 32496 23054 32548 23060
rect 32692 23050 32720 23258
rect 32680 23044 32732 23050
rect 32680 22986 32732 22992
rect 32496 22976 32548 22982
rect 32496 22918 32548 22924
rect 32508 22710 32536 22918
rect 32496 22704 32548 22710
rect 32496 22646 32548 22652
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 31576 22228 31628 22234
rect 31576 22170 31628 22176
rect 30852 22066 31064 22094
rect 31404 22066 31524 22094
rect 31036 21690 31064 22066
rect 30748 21684 30800 21690
rect 30748 21626 30800 21632
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 30656 21616 30708 21622
rect 30656 21558 30708 21564
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30116 21146 30144 21286
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30564 20460 30616 20466
rect 30564 20402 30616 20408
rect 30012 20392 30064 20398
rect 30012 20334 30064 20340
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 30012 20256 30064 20262
rect 30012 20198 30064 20204
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29564 18290 29592 18566
rect 29656 18358 29684 19790
rect 29748 19718 29776 20198
rect 30024 20058 30052 20198
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 29932 19378 29960 19654
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 30024 18358 30052 19994
rect 30208 19854 30236 20198
rect 30576 20058 30604 20402
rect 30668 20262 30696 21558
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30196 19848 30248 19854
rect 30196 19790 30248 19796
rect 31496 19378 31524 22066
rect 31760 21548 31812 21554
rect 31760 21490 31812 21496
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 31772 20942 31800 21490
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31668 20256 31720 20262
rect 31668 20198 31720 20204
rect 31680 19990 31708 20198
rect 31668 19984 31720 19990
rect 31668 19926 31720 19932
rect 31772 19378 31800 20878
rect 32220 20800 32272 20806
rect 32220 20742 32272 20748
rect 32036 20528 32088 20534
rect 32036 20470 32088 20476
rect 32048 20058 32076 20470
rect 32232 20466 32260 20742
rect 32220 20460 32272 20466
rect 32220 20402 32272 20408
rect 32600 20058 32628 21490
rect 32968 21010 32996 23276
rect 33048 23258 33100 23264
rect 34072 22642 34100 24822
rect 34244 24812 34296 24818
rect 34244 24754 34296 24760
rect 36084 24812 36136 24818
rect 36084 24754 36136 24760
rect 34256 23594 34284 24754
rect 35348 24608 35400 24614
rect 35348 24550 35400 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24410 35388 24550
rect 35348 24404 35400 24410
rect 35348 24346 35400 24352
rect 35532 24336 35584 24342
rect 35532 24278 35584 24284
rect 35348 23860 35400 23866
rect 35348 23802 35400 23808
rect 34704 23792 34756 23798
rect 34704 23734 34756 23740
rect 34244 23588 34296 23594
rect 34244 23530 34296 23536
rect 34716 23322 34744 23734
rect 35360 23594 35388 23802
rect 35544 23730 35572 24278
rect 35900 24268 35952 24274
rect 35900 24210 35952 24216
rect 35912 24154 35940 24210
rect 35820 24126 35940 24154
rect 35532 23724 35584 23730
rect 35532 23666 35584 23672
rect 35820 23662 35848 24126
rect 35900 24064 35952 24070
rect 35900 24006 35952 24012
rect 35912 23662 35940 24006
rect 36096 23866 36124 24754
rect 36820 24608 36872 24614
rect 36820 24550 36872 24556
rect 37004 24608 37056 24614
rect 37004 24550 37056 24556
rect 36268 24268 36320 24274
rect 36268 24210 36320 24216
rect 36084 23860 36136 23866
rect 36084 23802 36136 23808
rect 35624 23656 35676 23662
rect 35624 23598 35676 23604
rect 35808 23656 35860 23662
rect 35808 23598 35860 23604
rect 35900 23656 35952 23662
rect 35900 23598 35952 23604
rect 35348 23588 35400 23594
rect 35348 23530 35400 23536
rect 35440 23520 35492 23526
rect 35440 23462 35492 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34520 23316 34572 23322
rect 34520 23258 34572 23264
rect 34704 23316 34756 23322
rect 34704 23258 34756 23264
rect 35348 23316 35400 23322
rect 35348 23258 35400 23264
rect 34532 23118 34560 23258
rect 34520 23112 34572 23118
rect 34520 23054 34572 23060
rect 35360 22982 35388 23258
rect 35452 23118 35480 23462
rect 35636 23254 35664 23598
rect 35624 23248 35676 23254
rect 35624 23190 35676 23196
rect 35440 23112 35492 23118
rect 35440 23054 35492 23060
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 34808 22778 34836 22918
rect 34796 22772 34848 22778
rect 34796 22714 34848 22720
rect 34060 22636 34112 22642
rect 34060 22578 34112 22584
rect 33324 22568 33376 22574
rect 33244 22528 33324 22556
rect 33244 22166 33272 22528
rect 33324 22510 33376 22516
rect 34072 22166 34100 22578
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 33232 22160 33284 22166
rect 33232 22102 33284 22108
rect 34060 22160 34112 22166
rect 34060 22102 34112 22108
rect 34704 22160 34756 22166
rect 34704 22102 34756 22108
rect 33244 21026 33272 22102
rect 34072 21690 34100 22102
rect 34060 21684 34112 21690
rect 34060 21626 34112 21632
rect 33508 21548 33560 21554
rect 33508 21490 33560 21496
rect 33416 21344 33468 21350
rect 33416 21286 33468 21292
rect 33428 21146 33456 21286
rect 33416 21140 33468 21146
rect 33416 21082 33468 21088
rect 32956 21004 33008 21010
rect 32956 20946 33008 20952
rect 33152 20998 33272 21026
rect 32036 20052 32088 20058
rect 32036 19994 32088 20000
rect 32588 20052 32640 20058
rect 32588 19994 32640 20000
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32232 19446 32260 19790
rect 32968 19514 32996 20946
rect 33152 19938 33180 20998
rect 33232 20936 33284 20942
rect 33232 20878 33284 20884
rect 33244 20602 33272 20878
rect 33324 20800 33376 20806
rect 33324 20742 33376 20748
rect 33232 20596 33284 20602
rect 33232 20538 33284 20544
rect 33336 20466 33364 20742
rect 33324 20460 33376 20466
rect 33324 20402 33376 20408
rect 33324 20256 33376 20262
rect 33324 20198 33376 20204
rect 33336 19990 33364 20198
rect 33520 19990 33548 21490
rect 33692 21412 33744 21418
rect 33692 21354 33744 21360
rect 33704 21146 33732 21354
rect 33692 21140 33744 21146
rect 33692 21082 33744 21088
rect 34716 21010 34744 22102
rect 35256 22024 35308 22030
rect 35256 21966 35308 21972
rect 35268 21690 35296 21966
rect 35360 21690 35388 22918
rect 35452 22778 35480 23054
rect 36280 22778 36308 24210
rect 36544 24200 36596 24206
rect 36544 24142 36596 24148
rect 36728 24200 36780 24206
rect 36728 24142 36780 24148
rect 36452 24132 36504 24138
rect 36452 24074 36504 24080
rect 36360 24064 36412 24070
rect 36360 24006 36412 24012
rect 36372 23866 36400 24006
rect 36464 23866 36492 24074
rect 36360 23860 36412 23866
rect 36360 23802 36412 23808
rect 36452 23860 36504 23866
rect 36452 23802 36504 23808
rect 36464 23186 36492 23802
rect 36556 23798 36584 24142
rect 36544 23792 36596 23798
rect 36544 23734 36596 23740
rect 36556 23322 36584 23734
rect 36740 23322 36768 24142
rect 36832 23730 36860 24550
rect 37016 24410 37044 24550
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 37004 24404 37056 24410
rect 37004 24346 37056 24352
rect 37740 24132 37792 24138
rect 37740 24074 37792 24080
rect 37556 24064 37608 24070
rect 37556 24006 37608 24012
rect 36820 23724 36872 23730
rect 36820 23666 36872 23672
rect 37188 23724 37240 23730
rect 37188 23666 37240 23672
rect 36832 23594 36860 23666
rect 36820 23588 36872 23594
rect 36820 23530 36872 23536
rect 36544 23316 36596 23322
rect 36544 23258 36596 23264
rect 36728 23316 36780 23322
rect 36728 23258 36780 23264
rect 36832 23304 36860 23530
rect 37096 23316 37148 23322
rect 36832 23276 37096 23304
rect 36452 23180 36504 23186
rect 36452 23122 36504 23128
rect 36556 23118 36584 23258
rect 36544 23112 36596 23118
rect 36544 23054 36596 23060
rect 36832 22982 36860 23276
rect 37096 23258 37148 23264
rect 37200 23186 37228 23666
rect 37372 23520 37424 23526
rect 37372 23462 37424 23468
rect 37464 23520 37516 23526
rect 37464 23462 37516 23468
rect 37384 23186 37412 23462
rect 37188 23180 37240 23186
rect 37188 23122 37240 23128
rect 37372 23180 37424 23186
rect 37372 23122 37424 23128
rect 37476 23118 37504 23462
rect 37568 23254 37596 24006
rect 37752 23322 37780 24074
rect 37832 24064 37884 24070
rect 37832 24006 37884 24012
rect 38292 24064 38344 24070
rect 38292 24006 38344 24012
rect 37844 23662 37872 24006
rect 37832 23656 37884 23662
rect 37832 23598 37884 23604
rect 37740 23316 37792 23322
rect 37740 23258 37792 23264
rect 37556 23248 37608 23254
rect 37556 23190 37608 23196
rect 37464 23112 37516 23118
rect 37464 23054 37516 23060
rect 36820 22976 36872 22982
rect 36820 22918 36872 22924
rect 37740 22976 37792 22982
rect 37740 22918 37792 22924
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 35624 22772 35676 22778
rect 35624 22714 35676 22720
rect 36268 22772 36320 22778
rect 36268 22714 36320 22720
rect 35636 22098 35664 22714
rect 37372 22704 37424 22710
rect 37372 22646 37424 22652
rect 35624 22092 35676 22098
rect 35624 22034 35676 22040
rect 36544 21888 36596 21894
rect 36544 21830 36596 21836
rect 37280 21888 37332 21894
rect 37280 21830 37332 21836
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 36556 21554 36584 21830
rect 36544 21548 36596 21554
rect 36544 21490 36596 21496
rect 36636 21548 36688 21554
rect 36636 21490 36688 21496
rect 34796 21344 34848 21350
rect 34796 21286 34848 21292
rect 36084 21344 36136 21350
rect 36084 21286 36136 21292
rect 34704 21004 34756 21010
rect 34704 20946 34756 20952
rect 33600 20936 33652 20942
rect 33600 20878 33652 20884
rect 33612 20482 33640 20878
rect 33784 20800 33836 20806
rect 33784 20742 33836 20748
rect 34060 20800 34112 20806
rect 34060 20742 34112 20748
rect 33612 20454 33732 20482
rect 33600 20324 33652 20330
rect 33600 20266 33652 20272
rect 33324 19984 33376 19990
rect 33152 19910 33272 19938
rect 33324 19926 33376 19932
rect 33508 19984 33560 19990
rect 33508 19926 33560 19932
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 32956 19508 33008 19514
rect 32956 19450 33008 19456
rect 31852 19440 31904 19446
rect 31852 19382 31904 19388
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 31484 19372 31536 19378
rect 31404 19320 31484 19334
rect 31404 19314 31536 19320
rect 31576 19372 31628 19378
rect 31576 19314 31628 19320
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31404 19306 31524 19314
rect 31404 18737 31432 19306
rect 31390 18728 31446 18737
rect 30196 18692 30248 18698
rect 31390 18663 31392 18672
rect 30196 18634 30248 18640
rect 31444 18663 31446 18672
rect 31392 18634 31444 18640
rect 30208 18358 30236 18634
rect 29644 18352 29696 18358
rect 29644 18294 29696 18300
rect 30012 18352 30064 18358
rect 30012 18294 30064 18300
rect 30196 18352 30248 18358
rect 30196 18294 30248 18300
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 31300 18080 31352 18086
rect 31300 18022 31352 18028
rect 29736 17876 29788 17882
rect 29736 17818 29788 17824
rect 29748 17610 29776 17818
rect 31312 17678 31340 18022
rect 31404 17882 31432 18634
rect 31588 18290 31616 19314
rect 31864 18970 31892 19382
rect 32864 19168 32916 19174
rect 32864 19110 32916 19116
rect 32876 18970 32904 19110
rect 31852 18964 31904 18970
rect 31852 18906 31904 18912
rect 32864 18964 32916 18970
rect 32864 18906 32916 18912
rect 31852 18420 31904 18426
rect 31852 18362 31904 18368
rect 31760 18352 31812 18358
rect 31760 18294 31812 18300
rect 31576 18284 31628 18290
rect 31576 18226 31628 18232
rect 31576 18080 31628 18086
rect 31576 18022 31628 18028
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 30748 17672 30800 17678
rect 30748 17614 30800 17620
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 29736 17604 29788 17610
rect 29736 17546 29788 17552
rect 30196 17604 30248 17610
rect 30196 17546 30248 17552
rect 29368 17536 29420 17542
rect 29368 17478 29420 17484
rect 30012 17536 30064 17542
rect 30012 17478 30064 17484
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 29368 16448 29420 16454
rect 29368 16390 29420 16396
rect 29380 16250 29408 16390
rect 29368 16244 29420 16250
rect 29368 16186 29420 16192
rect 29276 16108 29328 16114
rect 29276 16050 29328 16056
rect 29380 16046 29408 16186
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 28908 15156 28960 15162
rect 28908 15098 28960 15104
rect 29012 15042 29040 15982
rect 29368 15632 29420 15638
rect 29368 15574 29420 15580
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 29104 15162 29132 15438
rect 29092 15156 29144 15162
rect 29092 15098 29144 15104
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28828 15014 29040 15042
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 28644 14074 28672 14214
rect 28632 14068 28684 14074
rect 28632 14010 28684 14016
rect 28828 12434 28856 15014
rect 29276 14816 29328 14822
rect 29276 14758 29328 14764
rect 29288 14618 29316 14758
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 29012 12850 29040 13806
rect 29000 12844 29052 12850
rect 29000 12786 29052 12792
rect 28828 12406 28948 12434
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 28644 11354 28672 12106
rect 28920 11558 28948 12406
rect 29012 11694 29040 12786
rect 29276 12640 29328 12646
rect 29276 12582 29328 12588
rect 29288 12306 29316 12582
rect 29380 12442 29408 15574
rect 29472 15026 29500 16526
rect 30024 16250 30052 17478
rect 30208 17082 30236 17546
rect 30208 17054 30420 17082
rect 30012 16244 30064 16250
rect 30012 16186 30064 16192
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29644 15564 29696 15570
rect 29644 15506 29696 15512
rect 29552 15360 29604 15366
rect 29552 15302 29604 15308
rect 29564 15094 29592 15302
rect 29552 15088 29604 15094
rect 29552 15030 29604 15036
rect 29460 15020 29512 15026
rect 29460 14962 29512 14968
rect 29656 14414 29684 15506
rect 29932 14550 29960 15982
rect 30208 15638 30236 17054
rect 30392 16998 30420 17054
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 30380 16992 30432 16998
rect 30380 16934 30432 16940
rect 30300 16590 30328 16934
rect 30288 16584 30340 16590
rect 30288 16526 30340 16532
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 30300 16046 30328 16390
rect 30656 16108 30708 16114
rect 30656 16050 30708 16056
rect 30288 16040 30340 16046
rect 30288 15982 30340 15988
rect 30196 15632 30248 15638
rect 30196 15574 30248 15580
rect 30104 15496 30156 15502
rect 30104 15438 30156 15444
rect 29920 14544 29972 14550
rect 29920 14486 29972 14492
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29748 13530 29776 13874
rect 30116 13734 30144 15438
rect 30668 15366 30696 16050
rect 30760 15502 30788 17614
rect 31588 17202 31616 18022
rect 31772 17338 31800 18294
rect 31760 17332 31812 17338
rect 31760 17274 31812 17280
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31864 17134 31892 18362
rect 32968 18358 32996 19450
rect 33152 18766 33180 19790
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 33244 18442 33272 19910
rect 33612 19854 33640 20266
rect 33704 19990 33732 20454
rect 33692 19984 33744 19990
rect 33692 19926 33744 19932
rect 33508 19848 33560 19854
rect 33508 19790 33560 19796
rect 33600 19848 33652 19854
rect 33600 19790 33652 19796
rect 33692 19848 33744 19854
rect 33692 19790 33744 19796
rect 33520 19514 33548 19790
rect 33704 19530 33732 19790
rect 33796 19718 33824 20742
rect 33876 20256 33928 20262
rect 33876 20198 33928 20204
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33508 19508 33560 19514
rect 33508 19450 33560 19456
rect 33612 19502 33732 19530
rect 33324 19236 33376 19242
rect 33324 19178 33376 19184
rect 33336 18834 33364 19178
rect 33324 18828 33376 18834
rect 33324 18770 33376 18776
rect 33060 18414 33272 18442
rect 32956 18352 33008 18358
rect 32956 18294 33008 18300
rect 32036 18216 32088 18222
rect 32036 18158 32088 18164
rect 32128 18216 32180 18222
rect 32128 18158 32180 18164
rect 32048 17814 32076 18158
rect 32140 17882 32168 18158
rect 32220 18148 32272 18154
rect 32220 18090 32272 18096
rect 32232 17882 32260 18090
rect 32404 18080 32456 18086
rect 32404 18022 32456 18028
rect 32864 18080 32916 18086
rect 32864 18022 32916 18028
rect 32128 17876 32180 17882
rect 32128 17818 32180 17824
rect 32220 17876 32272 17882
rect 32220 17818 32272 17824
rect 32036 17808 32088 17814
rect 32036 17750 32088 17756
rect 32048 17202 32076 17750
rect 32416 17678 32444 18022
rect 32876 17746 32904 18022
rect 32864 17740 32916 17746
rect 32864 17682 32916 17688
rect 32404 17672 32456 17678
rect 32404 17614 32456 17620
rect 32036 17196 32088 17202
rect 32036 17138 32088 17144
rect 31760 17128 31812 17134
rect 31760 17070 31812 17076
rect 31852 17128 31904 17134
rect 31852 17070 31904 17076
rect 31772 16250 31800 17070
rect 32128 17060 32180 17066
rect 32128 17002 32180 17008
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 31484 16176 31536 16182
rect 31484 16118 31536 16124
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 31128 15706 31156 16050
rect 31208 16040 31260 16046
rect 31208 15982 31260 15988
rect 31116 15700 31168 15706
rect 31116 15642 31168 15648
rect 30748 15496 30800 15502
rect 30748 15438 30800 15444
rect 30656 15360 30708 15366
rect 30656 15302 30708 15308
rect 30104 13728 30156 13734
rect 30104 13670 30156 13676
rect 29736 13524 29788 13530
rect 29736 13466 29788 13472
rect 30116 13394 30144 13670
rect 30104 13388 30156 13394
rect 30104 13330 30156 13336
rect 30012 13320 30064 13326
rect 30012 13262 30064 13268
rect 30024 12986 30052 13262
rect 30564 13184 30616 13190
rect 30564 13126 30616 13132
rect 30576 12986 30604 13126
rect 30012 12980 30064 12986
rect 30012 12922 30064 12928
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30472 12708 30524 12714
rect 30472 12650 30524 12656
rect 29368 12436 29420 12442
rect 29368 12378 29420 12384
rect 29276 12300 29328 12306
rect 29276 12242 29328 12248
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 29276 12096 29328 12102
rect 29276 12038 29328 12044
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 29288 11898 29316 12038
rect 29276 11892 29328 11898
rect 29276 11834 29328 11840
rect 29000 11688 29052 11694
rect 29000 11630 29052 11636
rect 28908 11552 28960 11558
rect 28908 11494 28960 11500
rect 28632 11348 28684 11354
rect 28632 11290 28684 11296
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28448 10804 28500 10810
rect 28448 10746 28500 10752
rect 28552 10674 28580 11086
rect 28540 10668 28592 10674
rect 28540 10610 28592 10616
rect 28920 10606 28948 11494
rect 29012 10742 29040 11630
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 28908 10600 28960 10606
rect 28908 10542 28960 10548
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 28356 10464 28408 10470
rect 28356 10406 28408 10412
rect 28920 9994 28948 10542
rect 29288 10198 29316 10542
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29276 10192 29328 10198
rect 29276 10134 29328 10140
rect 28264 9988 28316 9994
rect 28264 9930 28316 9936
rect 28908 9988 28960 9994
rect 28908 9930 28960 9936
rect 28276 9518 28304 9930
rect 29564 9654 29592 10406
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 28264 9512 28316 9518
rect 28264 9454 28316 9460
rect 30024 9466 30052 11086
rect 30208 10742 30236 12038
rect 30392 11898 30420 12174
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30196 10736 30248 10742
rect 30196 10678 30248 10684
rect 30024 9438 30144 9466
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 30024 8974 30052 9318
rect 30012 8968 30064 8974
rect 30012 8910 30064 8916
rect 29368 8832 29420 8838
rect 29368 8774 29420 8780
rect 29380 8634 29408 8774
rect 29368 8628 29420 8634
rect 29368 8570 29420 8576
rect 28080 8560 28132 8566
rect 28080 8502 28132 8508
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 26332 7812 26384 7818
rect 26332 7754 26384 7760
rect 27896 7812 27948 7818
rect 27896 7754 27948 7760
rect 29276 7812 29328 7818
rect 29276 7754 29328 7760
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 26344 7546 26372 7754
rect 27908 7546 27936 7754
rect 29288 7546 29316 7754
rect 29552 7744 29604 7750
rect 29552 7686 29604 7692
rect 26332 7540 26384 7546
rect 26332 7482 26384 7488
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 29564 7478 29592 7686
rect 29552 7472 29604 7478
rect 28460 7398 28764 7426
rect 29552 7414 29604 7420
rect 28460 7274 28488 7398
rect 28540 7336 28592 7342
rect 28540 7278 28592 7284
rect 28632 7336 28684 7342
rect 28736 7324 28764 7398
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 28816 7336 28868 7342
rect 28736 7296 28816 7324
rect 28632 7278 28684 7284
rect 28816 7278 28868 7284
rect 28448 7268 28500 7274
rect 28448 7210 28500 7216
rect 28552 6934 28580 7278
rect 28644 7206 28672 7278
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28540 6928 28592 6934
rect 28540 6870 28592 6876
rect 28736 6866 28948 6882
rect 27896 6860 27948 6866
rect 27896 6802 27948 6808
rect 28736 6860 28960 6866
rect 28736 6854 28908 6860
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 25608 5642 25636 6734
rect 26608 6724 26660 6730
rect 26608 6666 26660 6672
rect 27436 6724 27488 6730
rect 27436 6666 27488 6672
rect 26620 6458 26648 6666
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26976 6316 27028 6322
rect 26976 6258 27028 6264
rect 25596 5636 25648 5642
rect 25596 5578 25648 5584
rect 25688 5636 25740 5642
rect 25688 5578 25740 5584
rect 26424 5636 26476 5642
rect 26424 5578 26476 5584
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 25608 4690 25636 5578
rect 25700 5370 25728 5578
rect 26436 5370 26464 5578
rect 25688 5364 25740 5370
rect 25688 5306 25740 5312
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 26988 5234 27016 6258
rect 27448 5914 27476 6666
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27540 6458 27568 6598
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 27908 6322 27936 6802
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 28356 6316 28408 6322
rect 28356 6258 28408 6264
rect 27988 6180 28040 6186
rect 27988 6122 28040 6128
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 28000 5778 28028 6122
rect 27988 5772 28040 5778
rect 27988 5714 28040 5720
rect 27252 5568 27304 5574
rect 27252 5510 27304 5516
rect 27712 5568 27764 5574
rect 27712 5510 27764 5516
rect 27264 5370 27292 5510
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27724 5234 27752 5510
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 26988 4146 27016 5170
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27068 5024 27120 5030
rect 27068 4966 27120 4972
rect 27080 4826 27108 4966
rect 27632 4826 27660 5102
rect 27068 4820 27120 4826
rect 27068 4762 27120 4768
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27068 4548 27120 4554
rect 27068 4490 27120 4496
rect 27080 4282 27108 4490
rect 27068 4276 27120 4282
rect 27068 4218 27120 4224
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 27448 3194 27476 4558
rect 28000 4554 28028 5714
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 28092 5166 28120 5646
rect 28368 5370 28396 6258
rect 28460 6254 28488 6734
rect 28632 6452 28684 6458
rect 28632 6394 28684 6400
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 28644 5710 28672 6394
rect 28736 6186 28764 6854
rect 28908 6802 28960 6808
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 28828 6458 28856 6734
rect 28908 6724 28960 6730
rect 28908 6666 28960 6672
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 28814 6352 28870 6361
rect 28814 6287 28816 6296
rect 28868 6287 28870 6296
rect 28816 6258 28868 6264
rect 28920 6254 28948 6666
rect 29012 6458 29040 7346
rect 29552 6996 29604 7002
rect 29552 6938 29604 6944
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 29564 6322 29592 6938
rect 29736 6656 29788 6662
rect 29736 6598 29788 6604
rect 29552 6316 29604 6322
rect 29552 6258 29604 6264
rect 28908 6248 28960 6254
rect 28908 6190 28960 6196
rect 28724 6180 28776 6186
rect 28724 6122 28776 6128
rect 28540 5704 28592 5710
rect 28540 5646 28592 5652
rect 28632 5704 28684 5710
rect 28632 5646 28684 5652
rect 28448 5568 28500 5574
rect 28448 5510 28500 5516
rect 28460 5370 28488 5510
rect 28356 5364 28408 5370
rect 28356 5306 28408 5312
rect 28448 5364 28500 5370
rect 28448 5306 28500 5312
rect 28080 5160 28132 5166
rect 28080 5102 28132 5108
rect 27988 4548 28040 4554
rect 27988 4490 28040 4496
rect 28368 4214 28396 5306
rect 28552 4826 28580 5646
rect 28644 5302 28672 5646
rect 28816 5568 28868 5574
rect 28816 5510 28868 5516
rect 28632 5296 28684 5302
rect 28632 5238 28684 5244
rect 28828 5234 28856 5510
rect 28724 5228 28776 5234
rect 28724 5170 28776 5176
rect 28816 5228 28868 5234
rect 28816 5170 28868 5176
rect 28540 4820 28592 4826
rect 28540 4762 28592 4768
rect 28632 4276 28684 4282
rect 28632 4218 28684 4224
rect 28356 4208 28408 4214
rect 28356 4150 28408 4156
rect 28356 4072 28408 4078
rect 28356 4014 28408 4020
rect 27804 3392 27856 3398
rect 27710 3360 27766 3369
rect 27804 3334 27856 3340
rect 27710 3295 27766 3304
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 9680 2440 9732 2446
rect 17408 2440 17460 2446
rect 9680 2382 9732 2388
rect 952 2145 980 2382
rect 938 2136 994 2145
rect 938 2071 994 2080
rect 1964 800 1992 2382
rect 4540 800 4568 2382
rect 7116 800 7144 2382
rect 9692 800 9720 2382
rect 12268 2366 12388 2394
rect 17408 2382 17460 2388
rect 12268 800 12296 2366
rect 12360 2310 12388 2366
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 17420 800 17448 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 22572 800 22600 2790
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25148 800 25176 2382
rect 27724 800 27752 3295
rect 27816 3126 27844 3334
rect 27804 3120 27856 3126
rect 27804 3062 27856 3068
rect 28368 2446 28396 4014
rect 28644 3602 28672 4218
rect 28736 4214 28764 5170
rect 28920 4758 28948 6190
rect 29564 5914 29592 6258
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29458 5400 29514 5409
rect 29000 5364 29052 5370
rect 29458 5335 29460 5344
rect 29000 5306 29052 5312
rect 29512 5335 29514 5344
rect 29460 5306 29512 5312
rect 28908 4752 28960 4758
rect 28908 4694 28960 4700
rect 29012 4486 29040 5306
rect 29472 5030 29500 5306
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 28724 4208 28776 4214
rect 28724 4150 28776 4156
rect 28908 4004 28960 4010
rect 28908 3946 28960 3952
rect 28724 3936 28776 3942
rect 28724 3878 28776 3884
rect 28736 3738 28764 3878
rect 28920 3738 28948 3946
rect 28724 3732 28776 3738
rect 28724 3674 28776 3680
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 28632 3596 28684 3602
rect 28632 3538 28684 3544
rect 29012 3398 29040 4422
rect 29564 4146 29592 5850
rect 29748 5794 29776 6598
rect 29840 6458 29868 7822
rect 29932 7206 29960 7890
rect 30012 7744 30064 7750
rect 30012 7686 30064 7692
rect 29920 7200 29972 7206
rect 29920 7142 29972 7148
rect 29828 6452 29880 6458
rect 29828 6394 29880 6400
rect 29932 6322 29960 7142
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 30024 6254 30052 7686
rect 30116 7410 30144 9438
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 30392 7954 30420 8910
rect 30380 7948 30432 7954
rect 30380 7890 30432 7896
rect 30484 7834 30512 12650
rect 30564 11552 30616 11558
rect 30564 11494 30616 11500
rect 30576 11286 30604 11494
rect 30564 11280 30616 11286
rect 30564 11222 30616 11228
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30576 10606 30604 11086
rect 30668 11082 30696 15302
rect 30760 15026 30788 15438
rect 30748 15020 30800 15026
rect 30748 14962 30800 14968
rect 31024 14952 31076 14958
rect 31024 14894 31076 14900
rect 31036 14618 31064 14894
rect 31024 14612 31076 14618
rect 31024 14554 31076 14560
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 30760 11082 30788 14418
rect 31128 14414 31156 15642
rect 31220 15162 31248 15982
rect 31208 15156 31260 15162
rect 31208 15098 31260 15104
rect 31496 14414 31524 16118
rect 32140 16046 32168 17002
rect 32128 16040 32180 16046
rect 32128 15982 32180 15988
rect 31852 15904 31904 15910
rect 31852 15846 31904 15852
rect 31668 15428 31720 15434
rect 31668 15370 31720 15376
rect 31680 15162 31708 15370
rect 31864 15162 31892 15846
rect 32968 15706 32996 18294
rect 33060 16794 33088 18414
rect 33336 18290 33364 18770
rect 33520 18630 33548 19450
rect 33612 19446 33640 19502
rect 33600 19440 33652 19446
rect 33600 19382 33652 19388
rect 33692 19372 33744 19378
rect 33692 19314 33744 19320
rect 33888 19334 33916 20198
rect 33968 19848 34020 19854
rect 33968 19790 34020 19796
rect 33980 19446 34008 19790
rect 34072 19514 34100 20742
rect 34716 20534 34744 20946
rect 34808 20942 34836 21286
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 20936 34848 20942
rect 34796 20878 34848 20884
rect 36096 20806 36124 21286
rect 36556 20874 36584 21490
rect 36268 20868 36320 20874
rect 36268 20810 36320 20816
rect 36544 20868 36596 20874
rect 36544 20810 36596 20816
rect 36084 20800 36136 20806
rect 36084 20742 36136 20748
rect 34704 20528 34756 20534
rect 34704 20470 34756 20476
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34336 19848 34388 19854
rect 34336 19790 34388 19796
rect 34060 19508 34112 19514
rect 34060 19450 34112 19456
rect 33968 19440 34020 19446
rect 33968 19382 34020 19388
rect 34060 19372 34112 19378
rect 33704 18630 33732 19314
rect 33888 19306 34008 19334
rect 34060 19314 34112 19320
rect 33980 18698 34008 19306
rect 34072 18970 34100 19314
rect 34152 19168 34204 19174
rect 34152 19110 34204 19116
rect 34060 18964 34112 18970
rect 34060 18906 34112 18912
rect 33968 18692 34020 18698
rect 33968 18634 34020 18640
rect 33508 18624 33560 18630
rect 33508 18566 33560 18572
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 33704 18426 33732 18566
rect 34164 18426 34192 19110
rect 33692 18420 33744 18426
rect 34152 18420 34204 18426
rect 33692 18362 33744 18368
rect 34072 18380 34152 18408
rect 33600 18352 33652 18358
rect 33600 18294 33652 18300
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 33612 17678 33640 18294
rect 34072 17882 34100 18380
rect 34152 18362 34204 18368
rect 34152 18148 34204 18154
rect 34152 18090 34204 18096
rect 34164 17882 34192 18090
rect 34060 17876 34112 17882
rect 34060 17818 34112 17824
rect 34152 17876 34204 17882
rect 34152 17818 34204 17824
rect 33600 17672 33652 17678
rect 33600 17614 33652 17620
rect 33968 17672 34020 17678
rect 34348 17660 34376 19790
rect 34532 19786 34560 20402
rect 34716 19922 34744 20470
rect 36096 20466 36124 20742
rect 36280 20466 36308 20810
rect 36648 20482 36676 21490
rect 37292 21350 37320 21830
rect 36912 21344 36964 21350
rect 36912 21286 36964 21292
rect 37280 21344 37332 21350
rect 37280 21286 37332 21292
rect 36924 21146 36952 21286
rect 36912 21140 36964 21146
rect 36912 21082 36964 21088
rect 37384 20482 37412 22646
rect 37464 22568 37516 22574
rect 37464 22510 37516 22516
rect 37476 22234 37504 22510
rect 37464 22228 37516 22234
rect 37464 22170 37516 22176
rect 37752 22030 37780 22918
rect 37844 22098 37872 23598
rect 38304 23594 38332 24006
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 38568 23792 38620 23798
rect 38568 23734 38620 23740
rect 38292 23588 38344 23594
rect 38292 23530 38344 23536
rect 38580 23526 38608 23734
rect 39304 23724 39356 23730
rect 39304 23666 39356 23672
rect 45560 23724 45612 23730
rect 45560 23666 45612 23672
rect 46848 23724 46900 23730
rect 46848 23666 46900 23672
rect 38384 23520 38436 23526
rect 38384 23462 38436 23468
rect 38568 23520 38620 23526
rect 38568 23462 38620 23468
rect 38396 23254 38424 23462
rect 38384 23248 38436 23254
rect 38384 23190 38436 23196
rect 38580 23186 38608 23462
rect 39316 23322 39344 23666
rect 45572 23474 45600 23666
rect 45480 23446 45600 23474
rect 46112 23520 46164 23526
rect 46112 23462 46164 23468
rect 39304 23316 39356 23322
rect 39304 23258 39356 23264
rect 38568 23180 38620 23186
rect 38568 23122 38620 23128
rect 45480 23118 45508 23446
rect 45468 23112 45520 23118
rect 45468 23054 45520 23060
rect 46124 23050 46152 23462
rect 46860 23254 46888 23666
rect 47032 23656 47084 23662
rect 47032 23598 47084 23604
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 46848 23248 46900 23254
rect 46848 23190 46900 23196
rect 46952 23118 46980 23462
rect 46940 23112 46992 23118
rect 46940 23054 46992 23060
rect 38016 23044 38068 23050
rect 38016 22986 38068 22992
rect 38292 23044 38344 23050
rect 38292 22986 38344 22992
rect 46112 23044 46164 23050
rect 46112 22986 46164 22992
rect 38028 22710 38056 22986
rect 38304 22778 38332 22986
rect 44456 22976 44508 22982
rect 44456 22918 44508 22924
rect 45100 22976 45152 22982
rect 45100 22918 45152 22924
rect 38292 22772 38344 22778
rect 38292 22714 38344 22720
rect 38016 22704 38068 22710
rect 38016 22646 38068 22652
rect 44088 22704 44140 22710
rect 44088 22646 44140 22652
rect 43628 22568 43680 22574
rect 43628 22510 43680 22516
rect 39028 22500 39080 22506
rect 39028 22442 39080 22448
rect 38752 22432 38804 22438
rect 38752 22374 38804 22380
rect 37832 22092 37884 22098
rect 38764 22094 38792 22374
rect 37832 22034 37884 22040
rect 38672 22066 38792 22094
rect 37740 22024 37792 22030
rect 37740 21966 37792 21972
rect 37464 21956 37516 21962
rect 37464 21898 37516 21904
rect 37476 21690 37504 21898
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37752 21486 37780 21966
rect 37740 21480 37792 21486
rect 37740 21422 37792 21428
rect 36084 20460 36136 20466
rect 36084 20402 36136 20408
rect 36268 20460 36320 20466
rect 36648 20454 36768 20482
rect 36268 20402 36320 20408
rect 36268 20256 36320 20262
rect 36268 20198 36320 20204
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34704 19916 34756 19922
rect 34704 19858 34756 19864
rect 34612 19848 34664 19854
rect 34612 19790 34664 19796
rect 34520 19780 34572 19786
rect 34520 19722 34572 19728
rect 34532 18766 34560 19722
rect 34624 18970 34652 19790
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 34808 19514 34836 19654
rect 34796 19508 34848 19514
rect 34796 19450 34848 19456
rect 36084 19304 36136 19310
rect 36084 19246 36136 19252
rect 35348 19168 35400 19174
rect 35348 19110 35400 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34612 18964 34664 18970
rect 34612 18906 34664 18912
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 35360 18698 35388 19110
rect 36096 18970 36124 19246
rect 36176 19168 36228 19174
rect 36176 19110 36228 19116
rect 36084 18964 36136 18970
rect 36084 18906 36136 18912
rect 36188 18766 36216 19110
rect 36280 18766 36308 20198
rect 36636 19780 36688 19786
rect 36636 19722 36688 19728
rect 36648 19514 36676 19722
rect 36740 19718 36768 20454
rect 37292 20454 37412 20482
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 36728 19712 36780 19718
rect 36728 19654 36780 19660
rect 37004 19712 37056 19718
rect 37004 19654 37056 19660
rect 36636 19508 36688 19514
rect 36636 19450 36688 19456
rect 36912 19304 36964 19310
rect 37016 19292 37044 19654
rect 37200 19334 37228 19790
rect 37292 19786 37320 20454
rect 37372 20324 37424 20330
rect 37372 20266 37424 20272
rect 37384 20058 37412 20266
rect 37844 20058 37872 22034
rect 38672 22030 38700 22066
rect 38660 22024 38712 22030
rect 38660 21966 38712 21972
rect 38292 21616 38344 21622
rect 38292 21558 38344 21564
rect 38304 20942 38332 21558
rect 39040 21350 39068 22442
rect 39212 21888 39264 21894
rect 39212 21830 39264 21836
rect 39224 21690 39252 21830
rect 39212 21684 39264 21690
rect 39212 21626 39264 21632
rect 42706 21584 42762 21593
rect 42432 21548 42484 21554
rect 43640 21554 43668 22510
rect 42706 21519 42708 21528
rect 42432 21490 42484 21496
rect 42760 21519 42762 21528
rect 42800 21548 42852 21554
rect 42708 21490 42760 21496
rect 42800 21490 42852 21496
rect 43628 21548 43680 21554
rect 43628 21490 43680 21496
rect 39028 21344 39080 21350
rect 39028 21286 39080 21292
rect 38660 21072 38712 21078
rect 38660 21014 38712 21020
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38016 20868 38068 20874
rect 38016 20810 38068 20816
rect 37924 20800 37976 20806
rect 37924 20742 37976 20748
rect 37936 20262 37964 20742
rect 38028 20398 38056 20810
rect 38292 20800 38344 20806
rect 38292 20742 38344 20748
rect 38016 20392 38068 20398
rect 38016 20334 38068 20340
rect 37924 20256 37976 20262
rect 37924 20198 37976 20204
rect 37372 20052 37424 20058
rect 37372 19994 37424 20000
rect 37832 20052 37884 20058
rect 37832 19994 37884 20000
rect 37280 19780 37332 19786
rect 37280 19722 37332 19728
rect 36964 19264 37044 19292
rect 37108 19306 37228 19334
rect 36912 19246 36964 19252
rect 36360 19236 36412 19242
rect 36360 19178 36412 19184
rect 36372 18766 36400 19178
rect 36740 19094 37044 19122
rect 36740 18834 36768 19094
rect 36820 18964 36872 18970
rect 36872 18924 36952 18952
rect 36820 18906 36872 18912
rect 36728 18828 36780 18834
rect 36728 18770 36780 18776
rect 36176 18760 36228 18766
rect 36176 18702 36228 18708
rect 36268 18760 36320 18766
rect 36268 18702 36320 18708
rect 36360 18760 36412 18766
rect 36360 18702 36412 18708
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 35348 18692 35400 18698
rect 35348 18634 35400 18640
rect 35360 18290 35388 18634
rect 35348 18284 35400 18290
rect 35348 18226 35400 18232
rect 35808 18284 35860 18290
rect 35808 18226 35860 18232
rect 34704 18216 34756 18222
rect 34704 18158 34756 18164
rect 34716 17678 34744 18158
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34428 17672 34480 17678
rect 34348 17632 34428 17660
rect 33968 17614 34020 17620
rect 34428 17614 34480 17620
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 33140 17536 33192 17542
rect 33140 17478 33192 17484
rect 33232 17536 33284 17542
rect 33232 17478 33284 17484
rect 33048 16788 33100 16794
rect 33048 16730 33100 16736
rect 33060 16114 33088 16730
rect 33048 16108 33100 16114
rect 33048 16050 33100 16056
rect 33152 15994 33180 17478
rect 33244 17202 33272 17478
rect 33612 17338 33640 17614
rect 33600 17332 33652 17338
rect 33600 17274 33652 17280
rect 33980 17202 34008 17614
rect 33232 17196 33284 17202
rect 33232 17138 33284 17144
rect 33968 17196 34020 17202
rect 33968 17138 34020 17144
rect 33416 16108 33468 16114
rect 33416 16050 33468 16056
rect 33152 15966 33272 15994
rect 33140 15904 33192 15910
rect 33140 15846 33192 15852
rect 32956 15700 33008 15706
rect 32956 15642 33008 15648
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 31668 15156 31720 15162
rect 31668 15098 31720 15104
rect 31852 15156 31904 15162
rect 31852 15098 31904 15104
rect 31864 14618 31892 15098
rect 32324 14958 32352 15438
rect 32312 14952 32364 14958
rect 32312 14894 32364 14900
rect 31852 14612 31904 14618
rect 31852 14554 31904 14560
rect 32968 14414 32996 15642
rect 33152 15434 33180 15846
rect 33140 15428 33192 15434
rect 33140 15370 33192 15376
rect 33140 15020 33192 15026
rect 33140 14962 33192 14968
rect 33152 14618 33180 14962
rect 33140 14612 33192 14618
rect 33140 14554 33192 14560
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 31484 14408 31536 14414
rect 31484 14350 31536 14356
rect 31944 14408 31996 14414
rect 32956 14408 33008 14414
rect 31944 14350 31996 14356
rect 31956 14074 31984 14350
rect 32600 14346 32720 14362
rect 32956 14350 33008 14356
rect 32600 14340 32732 14346
rect 32600 14334 32680 14340
rect 32496 14272 32548 14278
rect 32496 14214 32548 14220
rect 31944 14068 31996 14074
rect 31944 14010 31996 14016
rect 32220 13932 32272 13938
rect 32220 13874 32272 13880
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31668 13728 31720 13734
rect 31668 13670 31720 13676
rect 30932 12980 30984 12986
rect 30932 12922 30984 12928
rect 30944 12306 30972 12922
rect 31128 12850 31156 13670
rect 31680 13394 31708 13670
rect 31484 13388 31536 13394
rect 31668 13388 31720 13394
rect 31484 13330 31536 13336
rect 31588 13348 31668 13376
rect 31208 12980 31260 12986
rect 31208 12922 31260 12928
rect 31116 12844 31168 12850
rect 31116 12786 31168 12792
rect 30932 12300 30984 12306
rect 30932 12242 30984 12248
rect 30840 12232 30892 12238
rect 30840 12174 30892 12180
rect 30852 11558 30880 12174
rect 30944 11830 30972 12242
rect 30932 11824 30984 11830
rect 30932 11766 30984 11772
rect 31220 11762 31248 12922
rect 31392 12776 31444 12782
rect 31392 12718 31444 12724
rect 31404 11830 31432 12718
rect 31496 12374 31524 13330
rect 31588 12646 31616 13348
rect 31668 13330 31720 13336
rect 31944 13388 31996 13394
rect 31944 13330 31996 13336
rect 31956 12782 31984 13330
rect 32232 13326 32260 13874
rect 32508 13326 32536 14214
rect 32220 13320 32272 13326
rect 32220 13262 32272 13268
rect 32404 13320 32456 13326
rect 32404 13262 32456 13268
rect 32496 13320 32548 13326
rect 32496 13262 32548 13268
rect 32128 13184 32180 13190
rect 32128 13126 32180 13132
rect 32140 13002 32168 13126
rect 32048 12974 32168 13002
rect 32048 12918 32076 12974
rect 32036 12912 32088 12918
rect 32036 12854 32088 12860
rect 31668 12776 31720 12782
rect 31668 12718 31720 12724
rect 31944 12776 31996 12782
rect 31944 12718 31996 12724
rect 31576 12640 31628 12646
rect 31576 12582 31628 12588
rect 31484 12368 31536 12374
rect 31484 12310 31536 12316
rect 31392 11824 31444 11830
rect 31392 11766 31444 11772
rect 31496 11762 31524 12310
rect 31680 12306 31708 12718
rect 31668 12300 31720 12306
rect 31668 12242 31720 12248
rect 31668 12096 31720 12102
rect 31668 12038 31720 12044
rect 31680 11898 31708 12038
rect 31668 11892 31720 11898
rect 31668 11834 31720 11840
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31484 11756 31536 11762
rect 31484 11698 31536 11704
rect 32232 11694 32260 13262
rect 32416 12986 32444 13262
rect 32404 12980 32456 12986
rect 32404 12922 32456 12928
rect 32312 12436 32364 12442
rect 32600 12434 32628 14334
rect 32680 14282 32732 14288
rect 32772 14272 32824 14278
rect 32692 14220 32772 14226
rect 32692 14214 32824 14220
rect 32692 14198 32812 14214
rect 32692 12442 32720 14198
rect 33048 14000 33100 14006
rect 33048 13942 33100 13948
rect 33060 13326 33088 13942
rect 33244 13870 33272 15966
rect 33428 15026 33456 16050
rect 33784 16040 33836 16046
rect 33784 15982 33836 15988
rect 33796 15162 33824 15982
rect 34440 15473 34468 17614
rect 34716 17338 34744 17614
rect 34704 17332 34756 17338
rect 34704 17274 34756 17280
rect 35360 17270 35388 18226
rect 35820 17882 35848 18226
rect 36372 18086 36400 18702
rect 36360 18080 36412 18086
rect 36360 18022 36412 18028
rect 35808 17876 35860 17882
rect 35808 17818 35860 17824
rect 36176 17536 36228 17542
rect 36176 17478 36228 17484
rect 35348 17264 35400 17270
rect 35348 17206 35400 17212
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16454 35388 17206
rect 36188 17202 36216 17478
rect 36372 17338 36400 18022
rect 36464 17882 36492 18702
rect 36820 18692 36872 18698
rect 36820 18634 36872 18640
rect 36728 18624 36780 18630
rect 36832 18601 36860 18634
rect 36728 18566 36780 18572
rect 36818 18592 36874 18601
rect 36740 18204 36768 18566
rect 36818 18527 36874 18536
rect 36924 18340 36952 18924
rect 37016 18902 37044 19094
rect 37004 18896 37056 18902
rect 37004 18838 37056 18844
rect 37108 18766 37136 19306
rect 37096 18760 37148 18766
rect 37096 18702 37148 18708
rect 37188 18760 37240 18766
rect 37188 18702 37240 18708
rect 37004 18352 37056 18358
rect 36924 18312 37004 18340
rect 37004 18294 37056 18300
rect 37096 18216 37148 18222
rect 36740 18176 37096 18204
rect 37096 18158 37148 18164
rect 36912 18080 36964 18086
rect 36912 18022 36964 18028
rect 36452 17876 36504 17882
rect 36452 17818 36504 17824
rect 36464 17592 36492 17818
rect 36924 17678 36952 18022
rect 36912 17672 36964 17678
rect 36912 17614 36964 17620
rect 36636 17604 36688 17610
rect 36464 17564 36636 17592
rect 36360 17332 36412 17338
rect 36360 17274 36412 17280
rect 36464 17202 36492 17564
rect 36636 17546 36688 17552
rect 35900 17196 35952 17202
rect 35900 17138 35952 17144
rect 36176 17196 36228 17202
rect 36176 17138 36228 17144
rect 36452 17196 36504 17202
rect 36452 17138 36504 17144
rect 35624 16992 35676 16998
rect 35624 16934 35676 16940
rect 35636 16590 35664 16934
rect 35624 16584 35676 16590
rect 35624 16526 35676 16532
rect 35348 16448 35400 16454
rect 35348 16390 35400 16396
rect 34520 16108 34572 16114
rect 34520 16050 34572 16056
rect 34426 15464 34482 15473
rect 34348 15422 34426 15450
rect 33968 15360 34020 15366
rect 33968 15302 34020 15308
rect 33784 15156 33836 15162
rect 33784 15098 33836 15104
rect 33416 15020 33468 15026
rect 33416 14962 33468 14968
rect 33600 14816 33652 14822
rect 33600 14758 33652 14764
rect 33692 14816 33744 14822
rect 33692 14758 33744 14764
rect 33612 14618 33640 14758
rect 33600 14612 33652 14618
rect 33600 14554 33652 14560
rect 33324 14408 33376 14414
rect 33324 14350 33376 14356
rect 33232 13864 33284 13870
rect 33232 13806 33284 13812
rect 33336 13530 33364 14350
rect 33324 13524 33376 13530
rect 33324 13466 33376 13472
rect 33048 13320 33100 13326
rect 33048 13262 33100 13268
rect 32864 13252 32916 13258
rect 32864 13194 32916 13200
rect 32876 12986 32904 13194
rect 32864 12980 32916 12986
rect 32864 12922 32916 12928
rect 32772 12640 32824 12646
rect 32772 12582 32824 12588
rect 32312 12378 32364 12384
rect 32508 12406 32628 12434
rect 32680 12436 32732 12442
rect 32324 11898 32352 12378
rect 32404 12232 32456 12238
rect 32404 12174 32456 12180
rect 32312 11892 32364 11898
rect 32312 11834 32364 11840
rect 32220 11688 32272 11694
rect 32220 11630 32272 11636
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 31300 11552 31352 11558
rect 31300 11494 31352 11500
rect 30656 11076 30708 11082
rect 30656 11018 30708 11024
rect 30748 11076 30800 11082
rect 30748 11018 30800 11024
rect 30564 10600 30616 10606
rect 30564 10542 30616 10548
rect 30576 10062 30604 10542
rect 30748 10124 30800 10130
rect 30748 10066 30800 10072
rect 30564 10056 30616 10062
rect 30564 9998 30616 10004
rect 30760 9722 30788 10066
rect 30748 9716 30800 9722
rect 30748 9658 30800 9664
rect 30748 8288 30800 8294
rect 30748 8230 30800 8236
rect 30392 7818 30512 7834
rect 30760 7818 30788 8230
rect 30380 7812 30512 7818
rect 30432 7806 30512 7812
rect 30748 7812 30800 7818
rect 30380 7754 30432 7760
rect 30748 7754 30800 7760
rect 30852 7698 30880 11494
rect 30932 10124 30984 10130
rect 30932 10066 30984 10072
rect 30944 9722 30972 10066
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 31116 9920 31168 9926
rect 31116 9862 31168 9868
rect 31036 9722 31064 9862
rect 30932 9716 30984 9722
rect 30932 9658 30984 9664
rect 31024 9716 31076 9722
rect 31024 9658 31076 9664
rect 31128 9602 31156 9862
rect 30944 9586 31156 9602
rect 30932 9580 31156 9586
rect 30984 9574 31156 9580
rect 30932 9522 30984 9528
rect 31312 8974 31340 11494
rect 31392 11144 31444 11150
rect 31392 11086 31444 11092
rect 31404 10062 31432 11086
rect 31392 10056 31444 10062
rect 31392 9998 31444 10004
rect 31404 9722 31432 9998
rect 32220 9988 32272 9994
rect 32220 9930 32272 9936
rect 31392 9716 31444 9722
rect 31392 9658 31444 9664
rect 32232 9586 32260 9930
rect 32220 9580 32272 9586
rect 32220 9522 32272 9528
rect 31576 9512 31628 9518
rect 31576 9454 31628 9460
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 30760 7670 30880 7698
rect 30104 7404 30156 7410
rect 30104 7346 30156 7352
rect 30380 7268 30432 7274
rect 30380 7210 30432 7216
rect 30104 6656 30156 6662
rect 30104 6598 30156 6604
rect 30116 6458 30144 6598
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 30012 6248 30064 6254
rect 30012 6190 30064 6196
rect 29748 5778 29960 5794
rect 29748 5772 29972 5778
rect 29748 5766 29920 5772
rect 29920 5714 29972 5720
rect 30024 5710 30052 6190
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 30288 6112 30340 6118
rect 30288 6054 30340 6060
rect 30116 5710 30144 6054
rect 30300 5914 30328 6054
rect 30392 5914 30420 7210
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30656 6316 30708 6322
rect 30656 6258 30708 6264
rect 30288 5908 30340 5914
rect 30288 5850 30340 5856
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 29828 5704 29880 5710
rect 29828 5646 29880 5652
rect 30012 5704 30064 5710
rect 30012 5646 30064 5652
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 29840 5370 29868 5646
rect 29828 5364 29880 5370
rect 29828 5306 29880 5312
rect 30392 5166 30420 5646
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30484 4826 30512 6258
rect 30576 5778 30604 6258
rect 30564 5772 30616 5778
rect 30564 5714 30616 5720
rect 30472 4820 30524 4826
rect 30472 4762 30524 4768
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 30104 4140 30156 4146
rect 30104 4082 30156 4088
rect 29104 3466 29132 4082
rect 29828 3936 29880 3942
rect 29828 3878 29880 3884
rect 29092 3460 29144 3466
rect 29092 3402 29144 3408
rect 29000 3392 29052 3398
rect 29000 3334 29052 3340
rect 28448 3120 28500 3126
rect 28448 3062 28500 3068
rect 28460 2650 28488 3062
rect 29104 2922 29132 3402
rect 29840 3194 29868 3878
rect 30116 3738 30144 4082
rect 30484 3942 30512 4762
rect 30576 4554 30604 5714
rect 30668 5370 30696 6258
rect 30760 5778 30788 7670
rect 31116 7472 31168 7478
rect 31116 7414 31168 7420
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 30852 6361 30880 6598
rect 30838 6352 30894 6361
rect 30838 6287 30894 6296
rect 31024 6112 31076 6118
rect 31024 6054 31076 6060
rect 30748 5772 30800 5778
rect 30748 5714 30800 5720
rect 30840 5704 30892 5710
rect 30840 5646 30892 5652
rect 30852 5409 30880 5646
rect 30838 5400 30894 5409
rect 30656 5364 30708 5370
rect 30838 5335 30894 5344
rect 30656 5306 30708 5312
rect 30932 5296 30984 5302
rect 30932 5238 30984 5244
rect 30656 5024 30708 5030
rect 30656 4966 30708 4972
rect 30668 4622 30696 4966
rect 30944 4622 30972 5238
rect 31036 5234 31064 6054
rect 31024 5228 31076 5234
rect 31024 5170 31076 5176
rect 30656 4616 30708 4622
rect 30932 4616 30984 4622
rect 30656 4558 30708 4564
rect 30760 4564 30932 4570
rect 30760 4558 30984 4564
rect 30564 4548 30616 4554
rect 30564 4490 30616 4496
rect 30668 4078 30696 4558
rect 30760 4542 30972 4558
rect 30656 4072 30708 4078
rect 30656 4014 30708 4020
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30472 3528 30524 3534
rect 30472 3470 30524 3476
rect 30484 3194 30512 3470
rect 30668 3466 30696 4014
rect 30760 3738 30788 4542
rect 30748 3732 30800 3738
rect 30748 3674 30800 3680
rect 30656 3460 30708 3466
rect 30656 3402 30708 3408
rect 29828 3188 29880 3194
rect 29828 3130 29880 3136
rect 30472 3188 30524 3194
rect 30472 3130 30524 3136
rect 30380 3120 30432 3126
rect 30380 3062 30432 3068
rect 29092 2916 29144 2922
rect 29092 2858 29144 2864
rect 30392 2650 30420 3062
rect 30668 2990 30696 3402
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 31128 2854 31156 7414
rect 31588 7410 31616 9454
rect 32416 8634 32444 12174
rect 32508 9586 32536 12406
rect 32680 12378 32732 12384
rect 32680 12096 32732 12102
rect 32680 12038 32732 12044
rect 32692 11762 32720 12038
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32600 11150 32628 11630
rect 32784 11626 32812 12582
rect 32876 12238 32904 12922
rect 32956 12436 33008 12442
rect 32956 12378 33008 12384
rect 32968 12238 32996 12378
rect 32864 12232 32916 12238
rect 32864 12174 32916 12180
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32864 12096 32916 12102
rect 32864 12038 32916 12044
rect 32772 11620 32824 11626
rect 32772 11562 32824 11568
rect 32680 11552 32732 11558
rect 32680 11494 32732 11500
rect 32692 11286 32720 11494
rect 32680 11280 32732 11286
rect 32680 11222 32732 11228
rect 32588 11144 32640 11150
rect 32588 11086 32640 11092
rect 32876 11014 32904 12038
rect 33060 11694 33088 13262
rect 33232 12640 33284 12646
rect 33232 12582 33284 12588
rect 33244 12434 33272 12582
rect 33704 12434 33732 14758
rect 33980 14482 34008 15302
rect 34244 14952 34296 14958
rect 34244 14894 34296 14900
rect 33968 14476 34020 14482
rect 33968 14418 34020 14424
rect 34256 13938 34284 14894
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 33968 13932 34020 13938
rect 33968 13874 34020 13880
rect 34244 13932 34296 13938
rect 34244 13874 34296 13880
rect 33796 12714 33824 13874
rect 33876 13728 33928 13734
rect 33876 13670 33928 13676
rect 33888 12850 33916 13670
rect 33980 12986 34008 13874
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 34060 13252 34112 13258
rect 34060 13194 34112 13200
rect 34072 12986 34100 13194
rect 34164 12986 34192 13806
rect 33968 12980 34020 12986
rect 33968 12922 34020 12928
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 34152 12980 34204 12986
rect 34152 12922 34204 12928
rect 33980 12850 34008 12922
rect 33876 12844 33928 12850
rect 33876 12786 33928 12792
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 33784 12708 33836 12714
rect 33784 12650 33836 12656
rect 33152 12406 33272 12434
rect 33612 12406 33732 12434
rect 33152 12306 33180 12406
rect 33140 12300 33192 12306
rect 33140 12242 33192 12248
rect 33612 12238 33640 12406
rect 33600 12232 33652 12238
rect 33600 12174 33652 12180
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 33704 11898 33732 12038
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 33048 11688 33100 11694
rect 33048 11630 33100 11636
rect 33968 11552 34020 11558
rect 33968 11494 34020 11500
rect 32772 11008 32824 11014
rect 32772 10950 32824 10956
rect 32864 11008 32916 11014
rect 32864 10950 32916 10956
rect 32784 10538 32812 10950
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 33048 10668 33100 10674
rect 33048 10610 33100 10616
rect 32772 10532 32824 10538
rect 32772 10474 32824 10480
rect 33060 10266 33088 10610
rect 33232 10464 33284 10470
rect 33232 10406 33284 10412
rect 33508 10464 33560 10470
rect 33508 10406 33560 10412
rect 33244 10266 33272 10406
rect 33048 10260 33100 10266
rect 33048 10202 33100 10208
rect 33232 10260 33284 10266
rect 33232 10202 33284 10208
rect 33520 10062 33548 10406
rect 33612 10062 33640 10746
rect 33692 10464 33744 10470
rect 33692 10406 33744 10412
rect 32772 10056 32824 10062
rect 32772 9998 32824 10004
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33600 10056 33652 10062
rect 33600 9998 33652 10004
rect 32680 9648 32732 9654
rect 32784 9636 32812 9998
rect 33048 9920 33100 9926
rect 33048 9862 33100 9868
rect 33060 9654 33088 9862
rect 32732 9608 32812 9636
rect 33048 9648 33100 9654
rect 32680 9590 32732 9596
rect 33048 9590 33100 9596
rect 32496 9580 32548 9586
rect 32496 9522 32548 9528
rect 33506 9480 33562 9489
rect 33506 9415 33562 9424
rect 33520 9382 33548 9415
rect 33508 9376 33560 9382
rect 33508 9318 33560 9324
rect 32772 8832 32824 8838
rect 32772 8774 32824 8780
rect 32784 8634 32812 8774
rect 32404 8628 32456 8634
rect 32404 8570 32456 8576
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32220 8084 32272 8090
rect 32220 8026 32272 8032
rect 31944 7880 31996 7886
rect 31944 7822 31996 7828
rect 31668 7812 31720 7818
rect 31668 7754 31720 7760
rect 31680 7546 31708 7754
rect 31956 7546 31984 7822
rect 31668 7540 31720 7546
rect 31668 7482 31720 7488
rect 31944 7540 31996 7546
rect 31944 7482 31996 7488
rect 31576 7404 31628 7410
rect 31576 7346 31628 7352
rect 31668 7404 31720 7410
rect 31668 7346 31720 7352
rect 31680 6390 31708 7346
rect 32232 7342 32260 8026
rect 32416 7478 32444 8570
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 32784 8090 32812 8366
rect 33232 8356 33284 8362
rect 33232 8298 33284 8304
rect 32772 8084 32824 8090
rect 32772 8026 32824 8032
rect 32772 7948 32824 7954
rect 32772 7890 32824 7896
rect 32404 7472 32456 7478
rect 32404 7414 32456 7420
rect 32784 7342 32812 7890
rect 33244 7426 33272 8298
rect 33324 8288 33376 8294
rect 33324 8230 33376 8236
rect 33336 7818 33364 8230
rect 33324 7812 33376 7818
rect 33324 7754 33376 7760
rect 33416 7744 33468 7750
rect 33416 7686 33468 7692
rect 33428 7546 33456 7686
rect 33416 7540 33468 7546
rect 33416 7482 33468 7488
rect 33244 7398 33364 7426
rect 32220 7336 32272 7342
rect 32220 7278 32272 7284
rect 32772 7336 32824 7342
rect 32772 7278 32824 7284
rect 33232 7336 33284 7342
rect 33232 7278 33284 7284
rect 32232 6866 32260 7278
rect 32220 6860 32272 6866
rect 32220 6802 32272 6808
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 31772 6458 31800 6734
rect 31760 6452 31812 6458
rect 31760 6394 31812 6400
rect 31668 6384 31720 6390
rect 31668 6326 31720 6332
rect 31576 6112 31628 6118
rect 31576 6054 31628 6060
rect 31588 5710 31616 6054
rect 31680 5778 31708 6326
rect 32508 6186 32536 6734
rect 32588 6656 32640 6662
rect 32588 6598 32640 6604
rect 32496 6180 32548 6186
rect 32496 6122 32548 6128
rect 31944 5908 31996 5914
rect 31944 5850 31996 5856
rect 31668 5772 31720 5778
rect 31668 5714 31720 5720
rect 31576 5704 31628 5710
rect 31576 5646 31628 5652
rect 31208 5636 31260 5642
rect 31208 5578 31260 5584
rect 31220 5166 31248 5578
rect 31484 5568 31536 5574
rect 31484 5510 31536 5516
rect 31576 5568 31628 5574
rect 31576 5510 31628 5516
rect 31496 5234 31524 5510
rect 31484 5228 31536 5234
rect 31484 5170 31536 5176
rect 31208 5160 31260 5166
rect 31208 5102 31260 5108
rect 31392 4548 31444 4554
rect 31392 4490 31444 4496
rect 31404 3466 31432 4490
rect 31588 4214 31616 5510
rect 31680 5370 31708 5714
rect 31956 5710 31984 5850
rect 32508 5710 32536 6122
rect 32600 5710 32628 6598
rect 32784 6254 32812 7278
rect 32864 7200 32916 7206
rect 32864 7142 32916 7148
rect 32772 6248 32824 6254
rect 32772 6190 32824 6196
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 32312 5704 32364 5710
rect 32312 5646 32364 5652
rect 32496 5704 32548 5710
rect 32496 5646 32548 5652
rect 32588 5704 32640 5710
rect 32588 5646 32640 5652
rect 31956 5370 31984 5646
rect 32128 5568 32180 5574
rect 32128 5510 32180 5516
rect 31668 5364 31720 5370
rect 31668 5306 31720 5312
rect 31944 5364 31996 5370
rect 31944 5306 31996 5312
rect 32140 5234 32168 5510
rect 32324 5370 32352 5646
rect 32312 5364 32364 5370
rect 32312 5306 32364 5312
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32496 5024 32548 5030
rect 32496 4966 32548 4972
rect 32508 4826 32536 4966
rect 32496 4820 32548 4826
rect 32496 4762 32548 4768
rect 32784 4690 32812 6190
rect 31852 4684 31904 4690
rect 31852 4626 31904 4632
rect 32772 4684 32824 4690
rect 32772 4626 32824 4632
rect 31668 4276 31720 4282
rect 31668 4218 31720 4224
rect 31576 4208 31628 4214
rect 31576 4150 31628 4156
rect 31392 3460 31444 3466
rect 31392 3402 31444 3408
rect 31404 2990 31432 3402
rect 31588 3194 31616 4150
rect 31680 3194 31708 4218
rect 31864 3602 31892 4626
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 31852 3596 31904 3602
rect 31852 3538 31904 3544
rect 31576 3188 31628 3194
rect 31576 3130 31628 3136
rect 31668 3188 31720 3194
rect 31668 3130 31720 3136
rect 32140 3058 32168 4082
rect 32312 3460 32364 3466
rect 32312 3402 32364 3408
rect 32324 3194 32352 3402
rect 32876 3194 32904 7142
rect 33244 6730 33272 7278
rect 33232 6724 33284 6730
rect 33232 6666 33284 6672
rect 33048 6248 33100 6254
rect 33048 6190 33100 6196
rect 33060 5914 33088 6190
rect 33048 5908 33100 5914
rect 33048 5850 33100 5856
rect 33140 5704 33192 5710
rect 33140 5646 33192 5652
rect 33152 5370 33180 5646
rect 33140 5364 33192 5370
rect 33140 5306 33192 5312
rect 33048 5024 33100 5030
rect 33048 4966 33100 4972
rect 33060 3466 33088 4966
rect 33140 4548 33192 4554
rect 33140 4490 33192 4496
rect 33152 4078 33180 4490
rect 33336 4146 33364 7398
rect 33428 6934 33456 7482
rect 33520 6934 33548 9318
rect 33612 8974 33640 9998
rect 33600 8968 33652 8974
rect 33600 8910 33652 8916
rect 33704 7546 33732 10406
rect 33980 8634 34008 11494
rect 34060 10600 34112 10606
rect 34060 10542 34112 10548
rect 34072 10266 34100 10542
rect 34060 10260 34112 10266
rect 34060 10202 34112 10208
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 33692 7540 33744 7546
rect 33692 7482 33744 7488
rect 33980 7206 34008 8570
rect 34256 8430 34284 13874
rect 34348 13802 34376 15422
rect 34426 15399 34482 15408
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 34440 14618 34468 15098
rect 34532 15026 34560 16050
rect 34612 15972 34664 15978
rect 34612 15914 34664 15920
rect 34520 15020 34572 15026
rect 34520 14962 34572 14968
rect 34428 14612 34480 14618
rect 34428 14554 34480 14560
rect 34532 14414 34560 14962
rect 34624 14618 34652 15914
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15502 35388 16390
rect 35348 15496 35400 15502
rect 35348 15438 35400 15444
rect 34796 15428 34848 15434
rect 34796 15370 34848 15376
rect 34704 15360 34756 15366
rect 34704 15302 34756 15308
rect 34716 15094 34744 15302
rect 34704 15088 34756 15094
rect 34704 15030 34756 15036
rect 34612 14612 34664 14618
rect 34612 14554 34664 14560
rect 34520 14408 34572 14414
rect 34520 14350 34572 14356
rect 34624 14226 34652 14554
rect 34716 14414 34744 15030
rect 34808 14618 34836 15370
rect 35360 15026 35388 15438
rect 35348 15020 35400 15026
rect 35348 14962 35400 14968
rect 35256 14816 35308 14822
rect 35308 14764 35480 14770
rect 35256 14758 35480 14764
rect 35268 14742 35480 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34796 14612 34848 14618
rect 34796 14554 34848 14560
rect 34704 14408 34756 14414
rect 34704 14350 34756 14356
rect 35348 14408 35400 14414
rect 35348 14350 35400 14356
rect 35072 14340 35124 14346
rect 35072 14282 35124 14288
rect 34532 14198 34652 14226
rect 34336 13796 34388 13802
rect 34336 13738 34388 13744
rect 34428 13184 34480 13190
rect 34428 13126 34480 13132
rect 34440 12918 34468 13126
rect 34428 12912 34480 12918
rect 34428 12854 34480 12860
rect 34532 12714 34560 14198
rect 34612 14068 34664 14074
rect 34612 14010 34664 14016
rect 34624 12918 34652 14010
rect 35084 13818 35112 14282
rect 35360 14074 35388 14350
rect 35348 14068 35400 14074
rect 35348 14010 35400 14016
rect 34808 13790 35112 13818
rect 34808 12918 34836 13790
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34612 12912 34664 12918
rect 34612 12854 34664 12860
rect 34796 12912 34848 12918
rect 34796 12854 34848 12860
rect 34808 12764 34836 12854
rect 34624 12736 34836 12764
rect 34520 12708 34572 12714
rect 34520 12650 34572 12656
rect 34624 12442 34652 12736
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34612 12436 34664 12442
rect 34612 12378 34664 12384
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 34612 11756 34664 11762
rect 34612 11698 34664 11704
rect 34520 10668 34572 10674
rect 34520 10610 34572 10616
rect 34532 9994 34560 10610
rect 34520 9988 34572 9994
rect 34520 9930 34572 9936
rect 34532 9722 34560 9930
rect 34520 9716 34572 9722
rect 34520 9658 34572 9664
rect 34428 9648 34480 9654
rect 34428 9590 34480 9596
rect 34440 9178 34468 9590
rect 34428 9172 34480 9178
rect 34428 9114 34480 9120
rect 34428 8900 34480 8906
rect 34428 8842 34480 8848
rect 34440 8430 34468 8842
rect 34624 8786 34652 11698
rect 34808 11150 34836 12174
rect 35072 12164 35124 12170
rect 35072 12106 35124 12112
rect 35084 11898 35112 12106
rect 35164 12096 35216 12102
rect 35164 12038 35216 12044
rect 35072 11892 35124 11898
rect 35072 11834 35124 11840
rect 35176 11762 35204 12038
rect 35164 11756 35216 11762
rect 35164 11698 35216 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 34808 10062 34836 11086
rect 35256 10600 35308 10606
rect 35452 10554 35480 14742
rect 35912 12646 35940 17138
rect 37108 16114 37136 18158
rect 37200 18154 37228 18702
rect 37292 18222 37320 19722
rect 37464 19304 37516 19310
rect 37464 19246 37516 19252
rect 37372 18624 37424 18630
rect 37372 18566 37424 18572
rect 37280 18216 37332 18222
rect 37280 18158 37332 18164
rect 37188 18148 37240 18154
rect 37188 18090 37240 18096
rect 37200 17814 37228 18090
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37188 17808 37240 17814
rect 37188 17750 37240 17756
rect 37292 17678 37320 18022
rect 37384 17882 37412 18566
rect 37372 17876 37424 17882
rect 37372 17818 37424 17824
rect 37188 17672 37240 17678
rect 37188 17614 37240 17620
rect 37280 17672 37332 17678
rect 37280 17614 37332 17620
rect 37096 16108 37148 16114
rect 37096 16050 37148 16056
rect 36084 15360 36136 15366
rect 36084 15302 36136 15308
rect 36096 13938 36124 15302
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 36360 14816 36412 14822
rect 36360 14758 36412 14764
rect 36372 14482 36400 14758
rect 36464 14618 36492 14962
rect 36544 14816 36596 14822
rect 36544 14758 36596 14764
rect 36728 14816 36780 14822
rect 36728 14758 36780 14764
rect 36820 14816 36872 14822
rect 36820 14758 36872 14764
rect 36452 14612 36504 14618
rect 36452 14554 36504 14560
rect 36360 14476 36412 14482
rect 36360 14418 36412 14424
rect 36084 13932 36136 13938
rect 36084 13874 36136 13880
rect 36556 13870 36584 14758
rect 36740 14482 36768 14758
rect 36728 14476 36780 14482
rect 36728 14418 36780 14424
rect 36728 14272 36780 14278
rect 36728 14214 36780 14220
rect 36740 13938 36768 14214
rect 36832 14006 36860 14758
rect 37108 14618 37136 16050
rect 37200 16028 37228 17614
rect 37280 16040 37332 16046
rect 37200 16000 37280 16028
rect 37280 15982 37332 15988
rect 37292 15502 37320 15982
rect 37476 15706 37504 19246
rect 38304 19174 38332 20742
rect 38672 20466 38700 21014
rect 39040 20942 39068 21286
rect 39684 21134 39896 21162
rect 39684 20942 39712 21134
rect 39764 21072 39816 21078
rect 39764 21014 39816 21020
rect 39028 20936 39080 20942
rect 39028 20878 39080 20884
rect 39672 20936 39724 20942
rect 39672 20878 39724 20884
rect 38752 20868 38804 20874
rect 38752 20810 38804 20816
rect 38764 20602 38792 20810
rect 38936 20800 38988 20806
rect 38936 20742 38988 20748
rect 39580 20800 39632 20806
rect 39776 20754 39804 21014
rect 39632 20748 39804 20754
rect 39580 20742 39804 20748
rect 38752 20596 38804 20602
rect 38752 20538 38804 20544
rect 38948 20534 38976 20742
rect 39592 20726 39804 20742
rect 38936 20528 38988 20534
rect 38936 20470 38988 20476
rect 39776 20466 39804 20726
rect 39868 20602 39896 21134
rect 40040 21140 40092 21146
rect 40040 21082 40092 21088
rect 39856 20596 39908 20602
rect 39856 20538 39908 20544
rect 38660 20460 38712 20466
rect 38660 20402 38712 20408
rect 39764 20460 39816 20466
rect 39764 20402 39816 20408
rect 40052 20398 40080 21082
rect 41328 20936 41380 20942
rect 41328 20878 41380 20884
rect 42340 20936 42392 20942
rect 42340 20878 42392 20884
rect 40316 20800 40368 20806
rect 40316 20742 40368 20748
rect 40408 20800 40460 20806
rect 40408 20742 40460 20748
rect 40040 20392 40092 20398
rect 40040 20334 40092 20340
rect 38660 20256 38712 20262
rect 38660 20198 38712 20204
rect 38844 20256 38896 20262
rect 38844 20198 38896 20204
rect 38672 19990 38700 20198
rect 38856 19990 38884 20198
rect 40224 20052 40276 20058
rect 40328 20040 40356 20742
rect 40420 20534 40448 20742
rect 41340 20534 41368 20878
rect 42352 20806 42380 20878
rect 42340 20800 42392 20806
rect 42340 20742 42392 20748
rect 42352 20602 42380 20742
rect 42340 20596 42392 20602
rect 42340 20538 42392 20544
rect 40408 20528 40460 20534
rect 40408 20470 40460 20476
rect 41328 20528 41380 20534
rect 41328 20470 41380 20476
rect 40500 20460 40552 20466
rect 40500 20402 40552 20408
rect 40868 20460 40920 20466
rect 40868 20402 40920 20408
rect 40276 20012 40356 20040
rect 40224 19994 40276 20000
rect 38660 19984 38712 19990
rect 38660 19926 38712 19932
rect 38844 19984 38896 19990
rect 38844 19926 38896 19932
rect 38384 19780 38436 19786
rect 38384 19722 38436 19728
rect 38292 19168 38344 19174
rect 38292 19110 38344 19116
rect 37924 18760 37976 18766
rect 37922 18728 37924 18737
rect 37976 18728 37978 18737
rect 38304 18698 38332 19110
rect 38396 18766 38424 19722
rect 40316 19712 40368 19718
rect 40316 19654 40368 19660
rect 39856 19372 39908 19378
rect 39856 19314 39908 19320
rect 39764 19168 39816 19174
rect 39764 19110 39816 19116
rect 39776 18902 39804 19110
rect 39396 18896 39448 18902
rect 39396 18838 39448 18844
rect 39764 18896 39816 18902
rect 39764 18838 39816 18844
rect 38384 18760 38436 18766
rect 38384 18702 38436 18708
rect 37922 18663 37978 18672
rect 38200 18692 38252 18698
rect 37832 18284 37884 18290
rect 37832 18226 37884 18232
rect 37844 17882 37872 18226
rect 37832 17876 37884 17882
rect 37832 17818 37884 17824
rect 37936 17678 37964 18663
rect 38200 18634 38252 18640
rect 38292 18692 38344 18698
rect 38292 18634 38344 18640
rect 38212 18426 38240 18634
rect 38304 18426 38332 18634
rect 38200 18420 38252 18426
rect 38200 18362 38252 18368
rect 38292 18420 38344 18426
rect 38292 18362 38344 18368
rect 38212 18154 38240 18362
rect 38396 18290 38424 18702
rect 38476 18692 38528 18698
rect 38476 18634 38528 18640
rect 38660 18692 38712 18698
rect 38660 18634 38712 18640
rect 38488 18601 38516 18634
rect 38474 18592 38530 18601
rect 38474 18527 38530 18536
rect 38384 18284 38436 18290
rect 38384 18226 38436 18232
rect 38200 18148 38252 18154
rect 38200 18090 38252 18096
rect 38568 18080 38620 18086
rect 38568 18022 38620 18028
rect 37924 17672 37976 17678
rect 37924 17614 37976 17620
rect 37832 17264 37884 17270
rect 37832 17206 37884 17212
rect 37844 16794 37872 17206
rect 37832 16788 37884 16794
rect 37832 16730 37884 16736
rect 37844 16182 37872 16730
rect 38198 16552 38254 16561
rect 38198 16487 38200 16496
rect 38252 16487 38254 16496
rect 38200 16458 38252 16464
rect 38016 16448 38068 16454
rect 38016 16390 38068 16396
rect 37832 16176 37884 16182
rect 37832 16118 37884 16124
rect 37464 15700 37516 15706
rect 37464 15642 37516 15648
rect 38028 15502 38056 16390
rect 38108 16176 38160 16182
rect 38108 16118 38160 16124
rect 38120 15706 38148 16118
rect 38108 15700 38160 15706
rect 38108 15642 38160 15648
rect 37280 15496 37332 15502
rect 37280 15438 37332 15444
rect 38016 15496 38068 15502
rect 38016 15438 38068 15444
rect 37096 14612 37148 14618
rect 37096 14554 37148 14560
rect 37004 14408 37056 14414
rect 37004 14350 37056 14356
rect 36820 14000 36872 14006
rect 36820 13942 36872 13948
rect 36912 14000 36964 14006
rect 36912 13942 36964 13948
rect 36728 13932 36780 13938
rect 36728 13874 36780 13880
rect 36544 13864 36596 13870
rect 36544 13806 36596 13812
rect 36268 13252 36320 13258
rect 36268 13194 36320 13200
rect 36280 12986 36308 13194
rect 36452 13184 36504 13190
rect 36452 13126 36504 13132
rect 36268 12980 36320 12986
rect 36268 12922 36320 12928
rect 36464 12918 36492 13126
rect 36832 12918 36860 13942
rect 36924 13802 36952 13942
rect 36912 13796 36964 13802
rect 36912 13738 36964 13744
rect 36452 12912 36504 12918
rect 36452 12854 36504 12860
rect 36820 12912 36872 12918
rect 36820 12854 36872 12860
rect 35900 12640 35952 12646
rect 35900 12582 35952 12588
rect 35912 12102 35940 12582
rect 36360 12164 36412 12170
rect 36360 12106 36412 12112
rect 35900 12096 35952 12102
rect 35900 12038 35952 12044
rect 36372 11898 36400 12106
rect 36360 11892 36412 11898
rect 36360 11834 36412 11840
rect 35808 11756 35860 11762
rect 36084 11756 36136 11762
rect 35860 11716 36084 11744
rect 35808 11698 35860 11704
rect 36084 11698 36136 11704
rect 36464 11694 36492 12854
rect 37016 12850 37044 14350
rect 37292 13938 37320 15438
rect 37556 15428 37608 15434
rect 37556 15370 37608 15376
rect 37464 14340 37516 14346
rect 37464 14282 37516 14288
rect 37280 13932 37332 13938
rect 37280 13874 37332 13880
rect 37476 13841 37504 14282
rect 37462 13832 37518 13841
rect 37462 13767 37518 13776
rect 36728 12844 36780 12850
rect 36728 12786 36780 12792
rect 37004 12844 37056 12850
rect 37004 12786 37056 12792
rect 37280 12844 37332 12850
rect 37280 12786 37332 12792
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 36740 12714 36768 12786
rect 37292 12730 37320 12786
rect 36728 12708 36780 12714
rect 37292 12702 37412 12730
rect 36728 12650 36780 12656
rect 36740 12434 36768 12650
rect 37280 12640 37332 12646
rect 37280 12582 37332 12588
rect 36740 12406 37136 12434
rect 37016 12374 37044 12406
rect 37004 12368 37056 12374
rect 37004 12310 37056 12316
rect 36912 12096 36964 12102
rect 36912 12038 36964 12044
rect 36924 11898 36952 12038
rect 36912 11892 36964 11898
rect 36912 11834 36964 11840
rect 36452 11688 36504 11694
rect 36452 11630 36504 11636
rect 36464 11558 36492 11630
rect 35808 11552 35860 11558
rect 35808 11494 35860 11500
rect 36452 11552 36504 11558
rect 36452 11494 36504 11500
rect 37004 11552 37056 11558
rect 37004 11494 37056 11500
rect 35820 11354 35848 11494
rect 35808 11348 35860 11354
rect 35808 11290 35860 11296
rect 35900 11348 35952 11354
rect 35900 11290 35952 11296
rect 35912 11234 35940 11290
rect 35820 11206 35940 11234
rect 35820 10606 35848 11206
rect 35308 10548 35480 10554
rect 35256 10542 35480 10548
rect 35808 10600 35860 10606
rect 35808 10542 35860 10548
rect 35268 10526 35480 10542
rect 35348 10464 35400 10470
rect 35348 10406 35400 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 10056 34848 10062
rect 34796 9998 34848 10004
rect 34796 9444 34848 9450
rect 34796 9386 34848 9392
rect 34808 9178 34836 9386
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 9172 34848 9178
rect 34796 9114 34848 9120
rect 35360 8906 35388 10406
rect 35452 10130 35480 10526
rect 35624 10192 35676 10198
rect 35624 10134 35676 10140
rect 35440 10124 35492 10130
rect 35440 10066 35492 10072
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 35348 8900 35400 8906
rect 35348 8842 35400 8848
rect 34532 8758 34652 8786
rect 34244 8424 34296 8430
rect 34244 8366 34296 8372
rect 34428 8424 34480 8430
rect 34428 8366 34480 8372
rect 34256 7342 34284 8366
rect 34440 7886 34468 8366
rect 34532 8090 34560 8758
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34716 8090 34744 8434
rect 34796 8288 34848 8294
rect 34796 8230 34848 8236
rect 34520 8084 34572 8090
rect 34520 8026 34572 8032
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 34532 7886 34560 8026
rect 34808 7886 34836 8230
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 34520 7880 34572 7886
rect 34520 7822 34572 7828
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 35256 7880 35308 7886
rect 35360 7868 35388 8842
rect 35544 8634 35572 9318
rect 35532 8628 35584 8634
rect 35532 8570 35584 8576
rect 35308 7840 35388 7868
rect 35256 7822 35308 7828
rect 34440 7410 34468 7822
rect 34428 7404 34480 7410
rect 34428 7346 34480 7352
rect 34244 7336 34296 7342
rect 34244 7278 34296 7284
rect 33968 7200 34020 7206
rect 33968 7142 34020 7148
rect 33416 6928 33468 6934
rect 33416 6870 33468 6876
rect 33508 6928 33560 6934
rect 33508 6870 33560 6876
rect 33428 5710 33456 6870
rect 34256 6866 34284 7278
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34244 6860 34296 6866
rect 34244 6802 34296 6808
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 33784 6656 33836 6662
rect 33784 6598 33836 6604
rect 33704 5914 33732 6598
rect 33796 6390 33824 6598
rect 33784 6384 33836 6390
rect 33784 6326 33836 6332
rect 33692 5908 33744 5914
rect 33692 5850 33744 5856
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 33876 5160 33928 5166
rect 33876 5102 33928 5108
rect 33600 5024 33652 5030
rect 33600 4966 33652 4972
rect 33612 4826 33640 4966
rect 33600 4820 33652 4826
rect 33600 4762 33652 4768
rect 33888 4690 33916 5102
rect 34072 4758 34100 6734
rect 35636 6662 35664 10134
rect 35820 9722 35848 10542
rect 35808 9716 35860 9722
rect 35808 9658 35860 9664
rect 35716 9580 35768 9586
rect 35716 9522 35768 9528
rect 35728 8838 35756 9522
rect 35820 9110 35848 9658
rect 35900 9580 35952 9586
rect 35900 9522 35952 9528
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35716 8832 35768 8838
rect 35716 8774 35768 8780
rect 35820 8362 35848 8910
rect 35912 8906 35940 9522
rect 36084 9512 36136 9518
rect 36084 9454 36136 9460
rect 36096 9178 36124 9454
rect 36084 9172 36136 9178
rect 36084 9114 36136 9120
rect 36464 9110 36492 11494
rect 37016 10742 37044 11494
rect 37108 11014 37136 12406
rect 37292 12306 37320 12582
rect 37384 12442 37412 12702
rect 37372 12436 37424 12442
rect 37372 12378 37424 12384
rect 37476 12306 37504 12786
rect 37280 12300 37332 12306
rect 37280 12242 37332 12248
rect 37464 12300 37516 12306
rect 37464 12242 37516 12248
rect 37476 11150 37504 12242
rect 37464 11144 37516 11150
rect 37464 11086 37516 11092
rect 37372 11076 37424 11082
rect 37372 11018 37424 11024
rect 37096 11008 37148 11014
rect 37096 10950 37148 10956
rect 37004 10736 37056 10742
rect 37004 10678 37056 10684
rect 36636 10464 36688 10470
rect 36636 10406 36688 10412
rect 36452 9104 36504 9110
rect 36452 9046 36504 9052
rect 35900 8900 35952 8906
rect 35900 8842 35952 8848
rect 36648 8498 36676 10406
rect 36728 9988 36780 9994
rect 36728 9930 36780 9936
rect 36740 9722 36768 9930
rect 36728 9716 36780 9722
rect 36728 9658 36780 9664
rect 37108 8974 37136 10950
rect 37384 10674 37412 11018
rect 37372 10668 37424 10674
rect 37372 10610 37424 10616
rect 37188 9920 37240 9926
rect 37188 9862 37240 9868
rect 37372 9920 37424 9926
rect 37372 9862 37424 9868
rect 37096 8968 37148 8974
rect 37096 8910 37148 8916
rect 37200 8838 37228 9862
rect 37384 8974 37412 9862
rect 37372 8968 37424 8974
rect 37372 8910 37424 8916
rect 37464 8968 37516 8974
rect 37464 8910 37516 8916
rect 37188 8832 37240 8838
rect 37188 8774 37240 8780
rect 37372 8832 37424 8838
rect 37372 8774 37424 8780
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 36636 8492 36688 8498
rect 36636 8434 36688 8440
rect 35808 8356 35860 8362
rect 35808 8298 35860 8304
rect 34520 6656 34572 6662
rect 34520 6598 34572 6604
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 35624 6656 35676 6662
rect 35624 6598 35676 6604
rect 34532 6118 34560 6598
rect 34520 6112 34572 6118
rect 34520 6054 34572 6060
rect 34532 5710 34560 6054
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34060 4752 34112 4758
rect 34060 4694 34112 4700
rect 33876 4684 33928 4690
rect 33876 4626 33928 4632
rect 33888 4146 33916 4626
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 33324 4140 33376 4146
rect 33324 4082 33376 4088
rect 33876 4140 33928 4146
rect 33876 4082 33928 4088
rect 33140 4072 33192 4078
rect 33140 4014 33192 4020
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 32312 3188 32364 3194
rect 32312 3130 32364 3136
rect 32864 3188 32916 3194
rect 32864 3130 32916 3136
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 31392 2984 31444 2990
rect 31392 2926 31444 2932
rect 31852 2916 31904 2922
rect 31852 2858 31904 2864
rect 31116 2848 31168 2854
rect 31116 2790 31168 2796
rect 31864 2774 31892 2858
rect 31772 2746 31892 2774
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 28356 2440 28408 2446
rect 30472 2440 30524 2446
rect 28356 2382 28408 2388
rect 30300 2400 30472 2428
rect 30300 800 30328 2400
rect 30472 2382 30524 2388
rect 31772 2378 31800 2746
rect 32140 2650 32168 2994
rect 33060 2990 33088 3402
rect 33888 2990 33916 4082
rect 34624 3534 34652 4558
rect 34612 3528 34664 3534
rect 34612 3470 34664 3476
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 33876 2984 33928 2990
rect 33876 2926 33928 2932
rect 34624 2650 34652 3470
rect 34716 3194 34744 6598
rect 35820 6322 35848 8298
rect 36280 8022 36308 8434
rect 36636 8288 36688 8294
rect 36636 8230 36688 8236
rect 36268 8016 36320 8022
rect 36268 7958 36320 7964
rect 36648 7886 36676 8230
rect 36636 7880 36688 7886
rect 36636 7822 36688 7828
rect 35900 7744 35952 7750
rect 35900 7686 35952 7692
rect 35992 7744 36044 7750
rect 35992 7686 36044 7692
rect 35912 7002 35940 7686
rect 36004 7546 36032 7686
rect 35992 7540 36044 7546
rect 35992 7482 36044 7488
rect 36268 7200 36320 7206
rect 36268 7142 36320 7148
rect 37004 7200 37056 7206
rect 37004 7142 37056 7148
rect 35900 6996 35952 7002
rect 35900 6938 35952 6944
rect 36084 6792 36136 6798
rect 36084 6734 36136 6740
rect 35808 6316 35860 6322
rect 35808 6258 35860 6264
rect 36096 6254 36124 6734
rect 36280 6390 36308 7142
rect 37016 6798 37044 7142
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 37188 6792 37240 6798
rect 37188 6734 37240 6740
rect 36268 6384 36320 6390
rect 36268 6326 36320 6332
rect 36360 6316 36412 6322
rect 36360 6258 36412 6264
rect 37096 6316 37148 6322
rect 37096 6258 37148 6264
rect 36084 6248 36136 6254
rect 36084 6190 36136 6196
rect 36176 6248 36228 6254
rect 36176 6190 36228 6196
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 36188 5914 36216 6190
rect 36176 5908 36228 5914
rect 36176 5850 36228 5856
rect 36176 5568 36228 5574
rect 36372 5556 36400 6258
rect 37004 6112 37056 6118
rect 37004 6054 37056 6060
rect 37016 5914 37044 6054
rect 37004 5908 37056 5914
rect 37004 5850 37056 5856
rect 37108 5846 37136 6258
rect 37096 5840 37148 5846
rect 37096 5782 37148 5788
rect 37200 5574 37228 6734
rect 37280 6656 37332 6662
rect 37280 6598 37332 6604
rect 37292 5914 37320 6598
rect 37384 6322 37412 8774
rect 37476 7410 37504 8910
rect 37568 8566 37596 15370
rect 38580 14278 38608 18022
rect 38672 17882 38700 18634
rect 38752 18624 38804 18630
rect 38752 18566 38804 18572
rect 38936 18624 38988 18630
rect 38936 18566 38988 18572
rect 38660 17876 38712 17882
rect 38660 17818 38712 17824
rect 38764 17338 38792 18566
rect 38948 18426 38976 18566
rect 38936 18420 38988 18426
rect 38936 18362 38988 18368
rect 38936 18284 38988 18290
rect 38936 18226 38988 18232
rect 38844 18148 38896 18154
rect 38844 18090 38896 18096
rect 38856 17338 38884 18090
rect 38752 17332 38804 17338
rect 38752 17274 38804 17280
rect 38844 17332 38896 17338
rect 38844 17274 38896 17280
rect 38948 17134 38976 18226
rect 38936 17128 38988 17134
rect 38936 17070 38988 17076
rect 39408 16794 39436 18838
rect 39488 18624 39540 18630
rect 39488 18566 39540 18572
rect 39500 17338 39528 18566
rect 39580 17536 39632 17542
rect 39580 17478 39632 17484
rect 39488 17332 39540 17338
rect 39488 17274 39540 17280
rect 39592 17202 39620 17478
rect 39580 17196 39632 17202
rect 39580 17138 39632 17144
rect 39396 16788 39448 16794
rect 39396 16730 39448 16736
rect 39028 16448 39080 16454
rect 39028 16390 39080 16396
rect 38660 15904 38712 15910
rect 38660 15846 38712 15852
rect 38672 15706 38700 15846
rect 38660 15700 38712 15706
rect 38660 15642 38712 15648
rect 38672 15162 38700 15642
rect 39040 15502 39068 16390
rect 39408 16266 39436 16730
rect 39488 16448 39540 16454
rect 39488 16390 39540 16396
rect 39316 16238 39436 16266
rect 39316 15570 39344 16238
rect 39396 16108 39448 16114
rect 39396 16050 39448 16056
rect 39408 15706 39436 16050
rect 39500 15910 39528 16390
rect 39488 15904 39540 15910
rect 39488 15846 39540 15852
rect 39396 15700 39448 15706
rect 39396 15642 39448 15648
rect 39304 15564 39356 15570
rect 39304 15506 39356 15512
rect 38844 15496 38896 15502
rect 38844 15438 38896 15444
rect 39028 15496 39080 15502
rect 39028 15438 39080 15444
rect 39210 15464 39266 15473
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38856 15094 38884 15438
rect 39210 15399 39212 15408
rect 39264 15399 39266 15408
rect 39212 15370 39264 15376
rect 38844 15088 38896 15094
rect 38844 15030 38896 15036
rect 39488 15020 39540 15026
rect 39488 14962 39540 14968
rect 39212 14952 39264 14958
rect 39212 14894 39264 14900
rect 38936 14816 38988 14822
rect 38936 14758 38988 14764
rect 38568 14272 38620 14278
rect 38568 14214 38620 14220
rect 37648 13252 37700 13258
rect 37648 13194 37700 13200
rect 37660 12986 37688 13194
rect 37648 12980 37700 12986
rect 37648 12922 37700 12928
rect 37832 12844 37884 12850
rect 37832 12786 37884 12792
rect 37924 12844 37976 12850
rect 37924 12786 37976 12792
rect 37844 12434 37872 12786
rect 37752 12406 37872 12434
rect 37752 11898 37780 12406
rect 37832 12232 37884 12238
rect 37832 12174 37884 12180
rect 37844 11898 37872 12174
rect 37740 11892 37792 11898
rect 37740 11834 37792 11840
rect 37832 11892 37884 11898
rect 37832 11834 37884 11840
rect 37936 11150 37964 12786
rect 38292 12640 38344 12646
rect 38292 12582 38344 12588
rect 38016 12164 38068 12170
rect 38016 12106 38068 12112
rect 37924 11144 37976 11150
rect 37924 11086 37976 11092
rect 37648 11008 37700 11014
rect 37648 10950 37700 10956
rect 37660 10538 37688 10950
rect 37740 10668 37792 10674
rect 37740 10610 37792 10616
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37752 10538 37780 10610
rect 37648 10532 37700 10538
rect 37648 10474 37700 10480
rect 37740 10532 37792 10538
rect 37740 10474 37792 10480
rect 37660 10062 37688 10474
rect 37648 10056 37700 10062
rect 37648 9998 37700 10004
rect 37844 9058 37872 10610
rect 37936 9654 37964 11086
rect 37924 9648 37976 9654
rect 37924 9590 37976 9596
rect 37752 9030 37872 9058
rect 37556 8560 37608 8566
rect 37556 8502 37608 8508
rect 37464 7404 37516 7410
rect 37464 7346 37516 7352
rect 37464 6792 37516 6798
rect 37464 6734 37516 6740
rect 37372 6316 37424 6322
rect 37372 6258 37424 6264
rect 37476 5914 37504 6734
rect 37280 5908 37332 5914
rect 37280 5850 37332 5856
rect 37464 5908 37516 5914
rect 37464 5850 37516 5856
rect 36452 5568 36504 5574
rect 36372 5528 36452 5556
rect 36176 5510 36228 5516
rect 36452 5510 36504 5516
rect 36820 5568 36872 5574
rect 36820 5510 36872 5516
rect 37188 5568 37240 5574
rect 37188 5510 37240 5516
rect 35440 5296 35492 5302
rect 35440 5238 35492 5244
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35452 4826 35480 5238
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 35440 4820 35492 4826
rect 35440 4762 35492 4768
rect 36004 4622 36032 5170
rect 36188 5166 36216 5510
rect 36464 5302 36492 5510
rect 36452 5296 36504 5302
rect 36452 5238 36504 5244
rect 36268 5228 36320 5234
rect 36268 5170 36320 5176
rect 36084 5160 36136 5166
rect 36084 5102 36136 5108
rect 36176 5160 36228 5166
rect 36176 5102 36228 5108
rect 36096 4826 36124 5102
rect 36084 4820 36136 4826
rect 36084 4762 36136 4768
rect 36280 4758 36308 5170
rect 36728 5160 36780 5166
rect 36728 5102 36780 5108
rect 36544 5092 36596 5098
rect 36544 5034 36596 5040
rect 36268 4752 36320 4758
rect 36268 4694 36320 4700
rect 36556 4622 36584 5034
rect 36636 5024 36688 5030
rect 36636 4966 36688 4972
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 35992 4480 36044 4486
rect 35992 4422 36044 4428
rect 36004 4282 36032 4422
rect 35992 4276 36044 4282
rect 35992 4218 36044 4224
rect 34796 4208 34848 4214
rect 34796 4150 34848 4156
rect 36452 4208 36504 4214
rect 36556 4162 36584 4558
rect 36648 4282 36676 4966
rect 36740 4622 36768 5102
rect 36832 4622 36860 5510
rect 37188 5024 37240 5030
rect 37188 4966 37240 4972
rect 36728 4616 36780 4622
rect 36728 4558 36780 4564
rect 36820 4616 36872 4622
rect 36820 4558 36872 4564
rect 36740 4282 36768 4558
rect 36636 4276 36688 4282
rect 36636 4218 36688 4224
rect 36728 4276 36780 4282
rect 36728 4218 36780 4224
rect 36504 4156 36584 4162
rect 36452 4150 36584 4156
rect 34808 3738 34836 4150
rect 36268 4140 36320 4146
rect 36464 4134 36584 4150
rect 36268 4082 36320 4088
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3732 34848 3738
rect 34796 3674 34848 3680
rect 36280 3534 36308 4082
rect 36556 3942 36584 4134
rect 36832 4010 36860 4558
rect 37200 4078 37228 4966
rect 37476 4826 37504 5850
rect 37752 5778 37780 9030
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37844 8634 37872 8910
rect 37832 8628 37884 8634
rect 37832 8570 37884 8576
rect 37936 8498 37964 9590
rect 38028 9586 38056 12106
rect 38304 11558 38332 12582
rect 38292 11552 38344 11558
rect 38292 11494 38344 11500
rect 38304 11150 38332 11494
rect 38108 11144 38160 11150
rect 38108 11086 38160 11092
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38120 10742 38148 11086
rect 38580 10810 38608 14214
rect 38660 13932 38712 13938
rect 38660 13874 38712 13880
rect 38672 12986 38700 13874
rect 38844 13864 38896 13870
rect 38844 13806 38896 13812
rect 38752 13728 38804 13734
rect 38752 13670 38804 13676
rect 38660 12980 38712 12986
rect 38660 12922 38712 12928
rect 38764 12918 38792 13670
rect 38856 13394 38884 13806
rect 38844 13388 38896 13394
rect 38844 13330 38896 13336
rect 38752 12912 38804 12918
rect 38752 12854 38804 12860
rect 38660 12708 38712 12714
rect 38660 12650 38712 12656
rect 38672 12442 38700 12650
rect 38764 12594 38792 12854
rect 38948 12714 38976 14758
rect 39028 14068 39080 14074
rect 39028 14010 39080 14016
rect 38936 12708 38988 12714
rect 38936 12650 38988 12656
rect 38764 12566 38884 12594
rect 38660 12436 38712 12442
rect 38660 12378 38712 12384
rect 38856 12238 38884 12566
rect 38948 12374 38976 12650
rect 38936 12368 38988 12374
rect 38936 12310 38988 12316
rect 38844 12232 38896 12238
rect 38844 12174 38896 12180
rect 38936 12232 38988 12238
rect 38936 12174 38988 12180
rect 38752 12096 38804 12102
rect 38752 12038 38804 12044
rect 38764 11762 38792 12038
rect 38752 11756 38804 11762
rect 38752 11698 38804 11704
rect 38844 11756 38896 11762
rect 38844 11698 38896 11704
rect 38856 11218 38884 11698
rect 38948 11354 38976 12174
rect 38936 11348 38988 11354
rect 38936 11290 38988 11296
rect 38844 11212 38896 11218
rect 38844 11154 38896 11160
rect 38568 10804 38620 10810
rect 38568 10746 38620 10752
rect 38108 10736 38160 10742
rect 38108 10678 38160 10684
rect 38292 10532 38344 10538
rect 38292 10474 38344 10480
rect 38304 10130 38332 10474
rect 38844 10464 38896 10470
rect 38844 10406 38896 10412
rect 38292 10124 38344 10130
rect 38292 10066 38344 10072
rect 38016 9580 38068 9586
rect 38016 9522 38068 9528
rect 38200 9512 38252 9518
rect 38198 9480 38200 9489
rect 38252 9480 38254 9489
rect 38198 9415 38254 9424
rect 38212 8498 38240 9415
rect 37924 8492 37976 8498
rect 37924 8434 37976 8440
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 37936 7954 37964 8434
rect 37924 7948 37976 7954
rect 37924 7890 37976 7896
rect 37936 7002 37964 7890
rect 37924 6996 37976 7002
rect 37924 6938 37976 6944
rect 38200 6792 38252 6798
rect 38200 6734 38252 6740
rect 37832 6112 37884 6118
rect 37832 6054 37884 6060
rect 37844 5778 37872 6054
rect 37740 5772 37792 5778
rect 37740 5714 37792 5720
rect 37832 5772 37884 5778
rect 37832 5714 37884 5720
rect 38212 5710 38240 6734
rect 38304 6390 38332 10066
rect 38384 8900 38436 8906
rect 38384 8842 38436 8848
rect 38396 8634 38424 8842
rect 38384 8628 38436 8634
rect 38384 8570 38436 8576
rect 38660 8424 38712 8430
rect 38660 8366 38712 8372
rect 38672 7970 38700 8366
rect 38580 7954 38700 7970
rect 38568 7948 38700 7954
rect 38620 7942 38700 7948
rect 38568 7890 38620 7896
rect 38660 6656 38712 6662
rect 38660 6598 38712 6604
rect 38292 6384 38344 6390
rect 38292 6326 38344 6332
rect 38292 6248 38344 6254
rect 38292 6190 38344 6196
rect 38200 5704 38252 5710
rect 38200 5646 38252 5652
rect 37464 4820 37516 4826
rect 37464 4762 37516 4768
rect 37476 4570 37504 4762
rect 38212 4622 38240 5646
rect 38200 4616 38252 4622
rect 37384 4554 37596 4570
rect 38200 4558 38252 4564
rect 37384 4548 37608 4554
rect 37384 4542 37556 4548
rect 37188 4072 37240 4078
rect 37188 4014 37240 4020
rect 36820 4004 36872 4010
rect 36820 3946 36872 3952
rect 36544 3936 36596 3942
rect 36544 3878 36596 3884
rect 36268 3528 36320 3534
rect 36268 3470 36320 3476
rect 36556 3466 36584 3878
rect 36832 3534 36860 3946
rect 37384 3602 37412 4542
rect 37556 4490 37608 4496
rect 38212 4486 38240 4558
rect 37464 4480 37516 4486
rect 37464 4422 37516 4428
rect 38200 4480 38252 4486
rect 38200 4422 38252 4428
rect 37476 4146 37504 4422
rect 38212 4282 38240 4422
rect 38200 4276 38252 4282
rect 38200 4218 38252 4224
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37740 4140 37792 4146
rect 37740 4082 37792 4088
rect 37556 3936 37608 3942
rect 37556 3878 37608 3884
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 36544 3460 36596 3466
rect 36544 3402 36596 3408
rect 35900 3392 35952 3398
rect 35900 3334 35952 3340
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 35348 2984 35400 2990
rect 35348 2926 35400 2932
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 2650 35388 2926
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 34612 2644 34664 2650
rect 34612 2586 34664 2592
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 35808 2576 35860 2582
rect 35808 2518 35860 2524
rect 33140 2440 33192 2446
rect 32876 2400 33140 2428
rect 31760 2372 31812 2378
rect 31760 2314 31812 2320
rect 32876 800 32904 2400
rect 33140 2382 33192 2388
rect 35452 870 35572 898
rect 35452 800 35480 870
rect 18 0 74 800
rect 1950 0 2006 800
rect 4526 0 4582 800
rect 7102 0 7158 800
rect 9678 0 9734 800
rect 12254 0 12310 800
rect 14830 0 14886 800
rect 17406 0 17462 800
rect 19982 0 20038 800
rect 22558 0 22614 800
rect 25134 0 25190 800
rect 27710 0 27766 800
rect 30286 0 30342 800
rect 32862 0 32918 800
rect 35438 0 35494 800
rect 35544 762 35572 870
rect 35820 762 35848 2518
rect 35912 2446 35940 3334
rect 37384 3194 37412 3538
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 36360 3120 36412 3126
rect 36360 3062 36412 3068
rect 36372 2650 36400 3062
rect 37568 2990 37596 3878
rect 37752 3738 37780 4082
rect 38106 4040 38162 4049
rect 38106 3975 38108 3984
rect 38160 3975 38162 3984
rect 38108 3946 38160 3952
rect 37740 3732 37792 3738
rect 37740 3674 37792 3680
rect 38212 3466 38240 4218
rect 38304 4010 38332 6190
rect 38568 6112 38620 6118
rect 38568 6054 38620 6060
rect 38580 5914 38608 6054
rect 38568 5908 38620 5914
rect 38568 5850 38620 5856
rect 38384 4752 38436 4758
rect 38384 4694 38436 4700
rect 38396 4282 38424 4694
rect 38672 4622 38700 6598
rect 38856 6458 38884 10406
rect 39040 10130 39068 14010
rect 39224 13530 39252 14894
rect 39500 14550 39528 14962
rect 39580 14816 39632 14822
rect 39580 14758 39632 14764
rect 39488 14544 39540 14550
rect 39488 14486 39540 14492
rect 39592 13530 39620 14758
rect 39764 14612 39816 14618
rect 39764 14554 39816 14560
rect 39672 14408 39724 14414
rect 39672 14350 39724 14356
rect 39684 13530 39712 14350
rect 39776 14074 39804 14554
rect 39764 14068 39816 14074
rect 39764 14010 39816 14016
rect 39868 13954 39896 19314
rect 40132 18760 40184 18766
rect 40132 18702 40184 18708
rect 39948 18352 40000 18358
rect 39948 18294 40000 18300
rect 39960 17270 39988 18294
rect 39948 17264 40000 17270
rect 39948 17206 40000 17212
rect 39960 16522 39988 17206
rect 39948 16516 40000 16522
rect 39948 16458 40000 16464
rect 39960 16250 39988 16458
rect 39948 16244 40000 16250
rect 39948 16186 40000 16192
rect 39960 15570 39988 16186
rect 40144 15638 40172 18702
rect 40224 16448 40276 16454
rect 40224 16390 40276 16396
rect 40236 16114 40264 16390
rect 40224 16108 40276 16114
rect 40224 16050 40276 16056
rect 40132 15632 40184 15638
rect 40132 15574 40184 15580
rect 39948 15564 40000 15570
rect 39948 15506 40000 15512
rect 40236 15502 40264 16050
rect 40224 15496 40276 15502
rect 40224 15438 40276 15444
rect 40132 14816 40184 14822
rect 40132 14758 40184 14764
rect 39776 13926 39896 13954
rect 39212 13524 39264 13530
rect 39212 13466 39264 13472
rect 39580 13524 39632 13530
rect 39580 13466 39632 13472
rect 39672 13524 39724 13530
rect 39672 13466 39724 13472
rect 39224 12850 39252 13466
rect 39212 12844 39264 12850
rect 39212 12786 39264 12792
rect 39776 12646 39804 13926
rect 39856 13864 39908 13870
rect 39856 13806 39908 13812
rect 39868 13326 39896 13806
rect 39856 13320 39908 13326
rect 39856 13262 39908 13268
rect 39764 12640 39816 12646
rect 39764 12582 39816 12588
rect 39396 12300 39448 12306
rect 39396 12242 39448 12248
rect 39120 11756 39172 11762
rect 39120 11698 39172 11704
rect 39132 11354 39160 11698
rect 39212 11552 39264 11558
rect 39212 11494 39264 11500
rect 39120 11348 39172 11354
rect 39120 11290 39172 11296
rect 39224 11150 39252 11494
rect 39408 11150 39436 12242
rect 39764 11348 39816 11354
rect 39764 11290 39816 11296
rect 39212 11144 39264 11150
rect 39212 11086 39264 11092
rect 39396 11144 39448 11150
rect 39396 11086 39448 11092
rect 39776 10606 39804 11290
rect 39868 11218 39896 13262
rect 39948 13184 40000 13190
rect 39948 13126 40000 13132
rect 39960 12918 39988 13126
rect 39948 12912 40000 12918
rect 39948 12854 40000 12860
rect 40144 12850 40172 14758
rect 40224 14476 40276 14482
rect 40224 14418 40276 14424
rect 40236 14074 40264 14418
rect 40328 14346 40356 19654
rect 40512 19514 40540 20402
rect 40684 20256 40736 20262
rect 40684 20198 40736 20204
rect 40696 19854 40724 20198
rect 40880 19990 40908 20402
rect 40868 19984 40920 19990
rect 40868 19926 40920 19932
rect 40684 19848 40736 19854
rect 40684 19790 40736 19796
rect 40500 19508 40552 19514
rect 40500 19450 40552 19456
rect 40880 19378 40908 19926
rect 41340 19530 41368 20470
rect 42444 20466 42472 21490
rect 42524 21344 42576 21350
rect 42524 21286 42576 21292
rect 42536 21146 42564 21286
rect 42524 21140 42576 21146
rect 42524 21082 42576 21088
rect 42812 20754 42840 21490
rect 44100 20942 44128 22646
rect 44364 22568 44416 22574
rect 44364 22510 44416 22516
rect 44376 22234 44404 22510
rect 44364 22228 44416 22234
rect 44364 22170 44416 22176
rect 44468 20942 44496 22918
rect 45008 22772 45060 22778
rect 45008 22714 45060 22720
rect 45020 22094 45048 22714
rect 45112 22710 45140 22918
rect 45100 22704 45152 22710
rect 45100 22646 45152 22652
rect 46572 22636 46624 22642
rect 46572 22578 46624 22584
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 44836 22066 45048 22094
rect 44836 22030 44864 22066
rect 44824 22024 44876 22030
rect 44824 21966 44876 21972
rect 45744 22024 45796 22030
rect 45744 21966 45796 21972
rect 45756 21622 45784 21966
rect 46204 21888 46256 21894
rect 46204 21830 46256 21836
rect 46216 21622 46244 21830
rect 46308 21678 46520 21706
rect 44548 21616 44600 21622
rect 44548 21558 44600 21564
rect 45744 21616 45796 21622
rect 45744 21558 45796 21564
rect 46204 21616 46256 21622
rect 46204 21558 46256 21564
rect 44560 21146 44588 21558
rect 45282 21448 45338 21457
rect 45282 21383 45338 21392
rect 44548 21140 44600 21146
rect 44548 21082 44600 21088
rect 45296 20942 45324 21383
rect 45756 21146 45784 21558
rect 46216 21146 46244 21558
rect 46308 21554 46336 21678
rect 46492 21622 46520 21678
rect 46584 21622 46612 22578
rect 46664 22432 46716 22438
rect 46664 22374 46716 22380
rect 46676 22030 46704 22374
rect 46756 22160 46808 22166
rect 46756 22102 46808 22108
rect 46664 22024 46716 22030
rect 46664 21966 46716 21972
rect 46768 21690 46796 22102
rect 46756 21684 46808 21690
rect 46756 21626 46808 21632
rect 46480 21616 46532 21622
rect 46480 21558 46532 21564
rect 46572 21616 46624 21622
rect 46572 21558 46624 21564
rect 46296 21548 46348 21554
rect 46296 21490 46348 21496
rect 46388 21548 46440 21554
rect 46388 21490 46440 21496
rect 46400 21434 46428 21490
rect 46480 21480 46532 21486
rect 46308 21428 46480 21434
rect 46308 21422 46532 21428
rect 46308 21406 46520 21422
rect 45744 21140 45796 21146
rect 45744 21082 45796 21088
rect 46204 21140 46256 21146
rect 46204 21082 46256 21088
rect 46308 21010 46336 21406
rect 46388 21344 46440 21350
rect 46388 21286 46440 21292
rect 46296 21004 46348 21010
rect 46296 20946 46348 20952
rect 44088 20936 44140 20942
rect 44088 20878 44140 20884
rect 44456 20936 44508 20942
rect 44456 20878 44508 20884
rect 45284 20936 45336 20942
rect 46400 20890 46428 21286
rect 46584 21146 46612 21558
rect 46860 21536 46888 22578
rect 46940 22024 46992 22030
rect 46940 21966 46992 21972
rect 46952 21690 46980 21966
rect 47044 21894 47072 23598
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 48044 23180 48096 23186
rect 48044 23122 48096 23128
rect 47952 23044 48004 23050
rect 47952 22986 48004 22992
rect 47584 22976 47636 22982
rect 47584 22918 47636 22924
rect 47124 22772 47176 22778
rect 47124 22714 47176 22720
rect 47032 21888 47084 21894
rect 47032 21830 47084 21836
rect 46940 21684 46992 21690
rect 46940 21626 46992 21632
rect 47032 21684 47084 21690
rect 47136 21672 47164 22714
rect 47308 22704 47360 22710
rect 47308 22646 47360 22652
rect 47320 22234 47348 22646
rect 47596 22574 47624 22918
rect 47584 22568 47636 22574
rect 47584 22510 47636 22516
rect 47400 22432 47452 22438
rect 47400 22374 47452 22380
rect 47308 22228 47360 22234
rect 47308 22170 47360 22176
rect 47412 22098 47440 22374
rect 47400 22092 47452 22098
rect 47400 22034 47452 22040
rect 47492 22024 47544 22030
rect 47492 21966 47544 21972
rect 47308 21956 47360 21962
rect 47308 21898 47360 21904
rect 47084 21644 47164 21672
rect 47032 21626 47084 21632
rect 47320 21622 47348 21898
rect 47308 21616 47360 21622
rect 47308 21558 47360 21564
rect 47032 21548 47084 21554
rect 46860 21508 47032 21536
rect 46572 21140 46624 21146
rect 46572 21082 46624 21088
rect 45284 20878 45336 20884
rect 42720 20726 42840 20754
rect 44180 20800 44232 20806
rect 44180 20742 44232 20748
rect 42720 20602 42748 20726
rect 42708 20596 42760 20602
rect 42708 20538 42760 20544
rect 43536 20528 43588 20534
rect 43536 20470 43588 20476
rect 42432 20460 42484 20466
rect 42432 20402 42484 20408
rect 41604 20392 41656 20398
rect 41604 20334 41656 20340
rect 42800 20392 42852 20398
rect 42800 20334 42852 20340
rect 41512 20256 41564 20262
rect 41512 20198 41564 20204
rect 41524 20058 41552 20198
rect 41512 20052 41564 20058
rect 41512 19994 41564 20000
rect 41248 19502 41368 19530
rect 41248 19446 41276 19502
rect 41236 19440 41288 19446
rect 41236 19382 41288 19388
rect 40408 19372 40460 19378
rect 40408 19314 40460 19320
rect 40868 19372 40920 19378
rect 40868 19314 40920 19320
rect 40420 15502 40448 19314
rect 41144 18964 41196 18970
rect 41144 18906 41196 18912
rect 41052 18692 41104 18698
rect 41052 18634 41104 18640
rect 41064 18426 41092 18634
rect 41052 18420 41104 18426
rect 41052 18362 41104 18368
rect 41156 18290 41184 18906
rect 41248 18698 41276 19382
rect 41328 19372 41380 19378
rect 41328 19314 41380 19320
rect 41236 18692 41288 18698
rect 41236 18634 41288 18640
rect 41340 18329 41368 19314
rect 41616 18630 41644 20334
rect 42812 20058 42840 20334
rect 43548 20058 43576 20470
rect 42800 20052 42852 20058
rect 42800 19994 42852 20000
rect 43536 20052 43588 20058
rect 43536 19994 43588 20000
rect 43444 19984 43496 19990
rect 43444 19926 43496 19932
rect 42616 19848 42668 19854
rect 42616 19790 42668 19796
rect 42628 19514 42656 19790
rect 42616 19508 42668 19514
rect 42616 19450 42668 19456
rect 43456 19446 43484 19926
rect 44192 19922 44220 20742
rect 45296 20602 45324 20878
rect 46216 20874 46428 20890
rect 46204 20868 46428 20874
rect 46256 20862 46428 20868
rect 46204 20810 46256 20816
rect 45284 20596 45336 20602
rect 45284 20538 45336 20544
rect 46112 20460 46164 20466
rect 46112 20402 46164 20408
rect 44272 20256 44324 20262
rect 44272 20198 44324 20204
rect 44456 20256 44508 20262
rect 44456 20198 44508 20204
rect 44180 19916 44232 19922
rect 44180 19858 44232 19864
rect 43444 19440 43496 19446
rect 43444 19382 43496 19388
rect 43628 19440 43680 19446
rect 43628 19382 43680 19388
rect 42524 19304 42576 19310
rect 42524 19246 42576 19252
rect 42536 18834 42564 19246
rect 42616 19168 42668 19174
rect 42616 19110 42668 19116
rect 42524 18828 42576 18834
rect 42524 18770 42576 18776
rect 41604 18624 41656 18630
rect 41604 18566 41656 18572
rect 42628 18426 42656 19110
rect 43456 18766 43484 19382
rect 43536 19304 43588 19310
rect 43536 19246 43588 19252
rect 43548 19174 43576 19246
rect 43536 19168 43588 19174
rect 43536 19110 43588 19116
rect 43444 18760 43496 18766
rect 43444 18702 43496 18708
rect 42616 18420 42668 18426
rect 42616 18362 42668 18368
rect 41326 18320 41382 18329
rect 41144 18284 41196 18290
rect 41144 18226 41196 18232
rect 41236 18284 41288 18290
rect 41326 18255 41328 18264
rect 41236 18226 41288 18232
rect 41380 18255 41382 18264
rect 41328 18226 41380 18232
rect 40960 17128 41012 17134
rect 40960 17070 41012 17076
rect 40868 16992 40920 16998
rect 40868 16934 40920 16940
rect 40880 16250 40908 16934
rect 40868 16244 40920 16250
rect 40868 16186 40920 16192
rect 40972 15978 41000 17070
rect 41248 17066 41276 18226
rect 43456 17882 43484 18702
rect 43444 17876 43496 17882
rect 43444 17818 43496 17824
rect 41604 17604 41656 17610
rect 41604 17546 41656 17552
rect 41616 17338 41644 17546
rect 43168 17536 43220 17542
rect 43168 17478 43220 17484
rect 41604 17332 41656 17338
rect 41604 17274 41656 17280
rect 42800 17128 42852 17134
rect 42800 17070 42852 17076
rect 41236 17060 41288 17066
rect 41236 17002 41288 17008
rect 42616 16652 42668 16658
rect 42616 16594 42668 16600
rect 42248 16448 42300 16454
rect 42248 16390 42300 16396
rect 42524 16448 42576 16454
rect 42524 16390 42576 16396
rect 42260 16250 42288 16390
rect 42536 16250 42564 16390
rect 42248 16244 42300 16250
rect 42248 16186 42300 16192
rect 42524 16244 42576 16250
rect 42524 16186 42576 16192
rect 41050 16144 41106 16153
rect 41050 16079 41052 16088
rect 41104 16079 41106 16088
rect 41052 16050 41104 16056
rect 40960 15972 41012 15978
rect 40960 15914 41012 15920
rect 40408 15496 40460 15502
rect 40408 15438 40460 15444
rect 40420 15162 40448 15438
rect 42628 15162 42656 16594
rect 42812 16182 42840 17070
rect 43180 16726 43208 17478
rect 43168 16720 43220 16726
rect 43168 16662 43220 16668
rect 42892 16516 42944 16522
rect 42892 16458 42944 16464
rect 42800 16176 42852 16182
rect 42800 16118 42852 16124
rect 42812 15570 42840 16118
rect 42904 15706 42932 16458
rect 43444 16448 43496 16454
rect 43444 16390 43496 16396
rect 43456 16182 43484 16390
rect 43444 16176 43496 16182
rect 43444 16118 43496 16124
rect 42892 15700 42944 15706
rect 42892 15642 42944 15648
rect 42800 15564 42852 15570
rect 42800 15506 42852 15512
rect 40408 15156 40460 15162
rect 40408 15098 40460 15104
rect 42616 15156 42668 15162
rect 42616 15098 42668 15104
rect 42904 15026 42932 15642
rect 43640 15570 43668 19382
rect 43720 19372 43772 19378
rect 43720 19314 43772 19320
rect 43732 18766 43760 19314
rect 44088 19304 44140 19310
rect 44088 19246 44140 19252
rect 43812 18828 43864 18834
rect 43812 18770 43864 18776
rect 43720 18760 43772 18766
rect 43720 18702 43772 18708
rect 43732 17814 43760 18702
rect 43720 17808 43772 17814
rect 43720 17750 43772 17756
rect 43824 17678 43852 18770
rect 43904 18760 43956 18766
rect 43904 18702 43956 18708
rect 43916 18154 43944 18702
rect 44100 18698 44128 19246
rect 44284 19242 44312 20198
rect 44468 19514 44496 20198
rect 46020 19916 46072 19922
rect 46020 19858 46072 19864
rect 44824 19848 44876 19854
rect 44824 19790 44876 19796
rect 44836 19514 44864 19790
rect 45468 19712 45520 19718
rect 45468 19654 45520 19660
rect 44456 19508 44508 19514
rect 44456 19450 44508 19456
rect 44824 19508 44876 19514
rect 44824 19450 44876 19456
rect 44272 19236 44324 19242
rect 44272 19178 44324 19184
rect 45008 18964 45060 18970
rect 45008 18906 45060 18912
rect 44364 18760 44416 18766
rect 44364 18702 44416 18708
rect 44088 18692 44140 18698
rect 44088 18634 44140 18640
rect 43904 18148 43956 18154
rect 43904 18090 43956 18096
rect 43916 17678 43944 18090
rect 44100 18086 44128 18634
rect 44376 18426 44404 18702
rect 44824 18692 44876 18698
rect 44824 18634 44876 18640
rect 44364 18420 44416 18426
rect 44364 18362 44416 18368
rect 44836 18290 44864 18634
rect 45020 18630 45048 18906
rect 45008 18624 45060 18630
rect 45008 18566 45060 18572
rect 44364 18284 44416 18290
rect 44364 18226 44416 18232
rect 44824 18284 44876 18290
rect 44824 18226 44876 18232
rect 44088 18080 44140 18086
rect 44088 18022 44140 18028
rect 44100 17882 44128 18022
rect 44088 17876 44140 17882
rect 44088 17818 44140 17824
rect 44376 17678 44404 18226
rect 43812 17672 43864 17678
rect 43812 17614 43864 17620
rect 43904 17672 43956 17678
rect 43904 17614 43956 17620
rect 44364 17672 44416 17678
rect 44364 17614 44416 17620
rect 44456 17672 44508 17678
rect 44456 17614 44508 17620
rect 44376 17338 44404 17614
rect 44364 17332 44416 17338
rect 44364 17274 44416 17280
rect 43904 17196 43956 17202
rect 43904 17138 43956 17144
rect 43812 16584 43864 16590
rect 43812 16526 43864 16532
rect 43824 15910 43852 16526
rect 43916 16250 43944 17138
rect 44088 16652 44140 16658
rect 44088 16594 44140 16600
rect 44100 16250 44128 16594
rect 44272 16584 44324 16590
rect 44192 16532 44272 16538
rect 44192 16526 44324 16532
rect 44192 16510 44312 16526
rect 43904 16244 43956 16250
rect 43904 16186 43956 16192
rect 44088 16244 44140 16250
rect 44088 16186 44140 16192
rect 44192 16153 44220 16510
rect 44272 16448 44324 16454
rect 44272 16390 44324 16396
rect 44178 16144 44234 16153
rect 44088 16108 44140 16114
rect 44178 16079 44234 16088
rect 44088 16050 44140 16056
rect 43812 15904 43864 15910
rect 43812 15846 43864 15852
rect 43628 15564 43680 15570
rect 43628 15506 43680 15512
rect 43824 15094 43852 15846
rect 43812 15088 43864 15094
rect 43812 15030 43864 15036
rect 40408 15020 40460 15026
rect 40408 14962 40460 14968
rect 40500 15020 40552 15026
rect 40500 14962 40552 14968
rect 40776 15020 40828 15026
rect 40776 14962 40828 14968
rect 42800 15020 42852 15026
rect 42800 14962 42852 14968
rect 42892 15020 42944 15026
rect 42892 14962 42944 14968
rect 40316 14340 40368 14346
rect 40316 14282 40368 14288
rect 40224 14068 40276 14074
rect 40224 14010 40276 14016
rect 40420 13954 40448 14962
rect 40512 14618 40540 14962
rect 40684 14816 40736 14822
rect 40684 14758 40736 14764
rect 40696 14618 40724 14758
rect 40500 14612 40552 14618
rect 40500 14554 40552 14560
rect 40684 14612 40736 14618
rect 40684 14554 40736 14560
rect 40500 14272 40552 14278
rect 40500 14214 40552 14220
rect 40512 14074 40540 14214
rect 40500 14068 40552 14074
rect 40500 14010 40552 14016
rect 40420 13926 40540 13954
rect 40512 13530 40540 13926
rect 40788 13734 40816 14962
rect 42248 14952 42300 14958
rect 42248 14894 42300 14900
rect 40960 14816 41012 14822
rect 40960 14758 41012 14764
rect 40972 13938 41000 14758
rect 42260 14618 42288 14894
rect 42248 14612 42300 14618
rect 42248 14554 42300 14560
rect 42812 14550 42840 14962
rect 42904 14618 42932 14962
rect 44100 14958 44128 16050
rect 44192 15366 44220 16079
rect 44180 15360 44232 15366
rect 44180 15302 44232 15308
rect 44284 14958 44312 16390
rect 44468 16046 44496 17614
rect 44916 16992 44968 16998
rect 44916 16934 44968 16940
rect 44548 16516 44600 16522
rect 44548 16458 44600 16464
rect 44456 16040 44508 16046
rect 44456 15982 44508 15988
rect 44364 15428 44416 15434
rect 44364 15370 44416 15376
rect 44376 15162 44404 15370
rect 44364 15156 44416 15162
rect 44364 15098 44416 15104
rect 43812 14952 43864 14958
rect 43812 14894 43864 14900
rect 44088 14952 44140 14958
rect 44088 14894 44140 14900
rect 44272 14952 44324 14958
rect 44272 14894 44324 14900
rect 42892 14612 42944 14618
rect 42892 14554 42944 14560
rect 42708 14544 42760 14550
rect 42708 14486 42760 14492
rect 42800 14544 42852 14550
rect 42800 14486 42852 14492
rect 42524 14408 42576 14414
rect 42720 14396 42748 14486
rect 43824 14414 43852 14894
rect 44100 14414 44128 14894
rect 44180 14816 44232 14822
rect 44180 14758 44232 14764
rect 43076 14408 43128 14414
rect 42720 14368 43076 14396
rect 42524 14350 42576 14356
rect 43076 14350 43128 14356
rect 43812 14408 43864 14414
rect 43812 14350 43864 14356
rect 44088 14408 44140 14414
rect 44088 14350 44140 14356
rect 41236 14272 41288 14278
rect 41236 14214 41288 14220
rect 42248 14272 42300 14278
rect 42248 14214 42300 14220
rect 40960 13932 41012 13938
rect 40960 13874 41012 13880
rect 40776 13728 40828 13734
rect 40776 13670 40828 13676
rect 40500 13524 40552 13530
rect 40500 13466 40552 13472
rect 40788 13444 40816 13670
rect 40868 13456 40920 13462
rect 40788 13416 40868 13444
rect 40868 13398 40920 13404
rect 41052 13252 41104 13258
rect 41052 13194 41104 13200
rect 41064 12986 41092 13194
rect 40224 12980 40276 12986
rect 40224 12922 40276 12928
rect 41052 12980 41104 12986
rect 41052 12922 41104 12928
rect 40040 12844 40092 12850
rect 40040 12786 40092 12792
rect 40132 12844 40184 12850
rect 40132 12786 40184 12792
rect 39856 11212 39908 11218
rect 39856 11154 39908 11160
rect 39764 10600 39816 10606
rect 39764 10542 39816 10548
rect 40052 10130 40080 12786
rect 40236 12238 40264 12922
rect 41248 12850 41276 14214
rect 42260 14074 42288 14214
rect 42248 14068 42300 14074
rect 42248 14010 42300 14016
rect 42536 13394 42564 14350
rect 43168 14272 43220 14278
rect 43168 14214 43220 14220
rect 43180 14074 43208 14214
rect 43168 14068 43220 14074
rect 43168 14010 43220 14016
rect 43824 13802 43852 14350
rect 43812 13796 43864 13802
rect 43812 13738 43864 13744
rect 42800 13728 42852 13734
rect 42800 13670 42852 13676
rect 42524 13388 42576 13394
rect 42524 13330 42576 13336
rect 42248 13320 42300 13326
rect 42248 13262 42300 13268
rect 42340 13320 42392 13326
rect 42812 13308 42840 13670
rect 42984 13320 43036 13326
rect 42812 13280 42984 13308
rect 42340 13262 42392 13268
rect 42984 13262 43036 13268
rect 42260 12850 42288 13262
rect 42352 12986 42380 13262
rect 42432 13184 42484 13190
rect 42432 13126 42484 13132
rect 42340 12980 42392 12986
rect 42340 12922 42392 12928
rect 41236 12844 41288 12850
rect 41236 12786 41288 12792
rect 42156 12844 42208 12850
rect 42156 12786 42208 12792
rect 42248 12844 42300 12850
rect 42248 12786 42300 12792
rect 40776 12640 40828 12646
rect 40776 12582 40828 12588
rect 40788 12434 40816 12582
rect 40788 12406 40908 12434
rect 40592 12368 40644 12374
rect 40592 12310 40644 12316
rect 40224 12232 40276 12238
rect 40224 12174 40276 12180
rect 40604 12102 40632 12310
rect 40880 12238 40908 12406
rect 40684 12232 40736 12238
rect 40684 12174 40736 12180
rect 40868 12232 40920 12238
rect 40868 12174 40920 12180
rect 41236 12232 41288 12238
rect 41236 12174 41288 12180
rect 40408 12096 40460 12102
rect 40408 12038 40460 12044
rect 40592 12096 40644 12102
rect 40592 12038 40644 12044
rect 40420 11762 40448 12038
rect 40604 11830 40632 12038
rect 40592 11824 40644 11830
rect 40592 11766 40644 11772
rect 40408 11756 40460 11762
rect 40408 11698 40460 11704
rect 40132 11076 40184 11082
rect 40132 11018 40184 11024
rect 40144 10538 40172 11018
rect 40132 10532 40184 10538
rect 40132 10474 40184 10480
rect 40590 10296 40646 10305
rect 40590 10231 40646 10240
rect 40604 10198 40632 10231
rect 40592 10192 40644 10198
rect 40592 10134 40644 10140
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 40040 10124 40092 10130
rect 40040 10066 40092 10072
rect 40696 10062 40724 12174
rect 40776 12096 40828 12102
rect 40776 12038 40828 12044
rect 40788 11694 40816 12038
rect 40776 11688 40828 11694
rect 40776 11630 40828 11636
rect 41144 11688 41196 11694
rect 41144 11630 41196 11636
rect 41156 10810 41184 11630
rect 41248 11354 41276 12174
rect 41604 12096 41656 12102
rect 41604 12038 41656 12044
rect 41616 11898 41644 12038
rect 42168 11898 42196 12786
rect 42260 12238 42288 12786
rect 42248 12232 42300 12238
rect 42248 12174 42300 12180
rect 41604 11892 41656 11898
rect 41604 11834 41656 11840
rect 42156 11892 42208 11898
rect 42156 11834 42208 11840
rect 42444 11694 42472 13126
rect 42800 12640 42852 12646
rect 42800 12582 42852 12588
rect 42432 11688 42484 11694
rect 42432 11630 42484 11636
rect 41696 11552 41748 11558
rect 41696 11494 41748 11500
rect 41880 11552 41932 11558
rect 41880 11494 41932 11500
rect 41236 11348 41288 11354
rect 41236 11290 41288 11296
rect 41328 11144 41380 11150
rect 41328 11086 41380 11092
rect 41144 10804 41196 10810
rect 41144 10746 41196 10752
rect 41340 10742 41368 11086
rect 41708 11082 41736 11494
rect 41696 11076 41748 11082
rect 41696 11018 41748 11024
rect 40776 10736 40828 10742
rect 40776 10678 40828 10684
rect 41328 10736 41380 10742
rect 41328 10678 41380 10684
rect 39580 10056 39632 10062
rect 39580 9998 39632 10004
rect 40684 10056 40736 10062
rect 40684 9998 40736 10004
rect 38936 9920 38988 9926
rect 38936 9862 38988 9868
rect 39120 9920 39172 9926
rect 39120 9862 39172 9868
rect 38948 9586 38976 9862
rect 39132 9586 39160 9862
rect 39592 9586 39620 9998
rect 40592 9920 40644 9926
rect 40592 9862 40644 9868
rect 40604 9654 40632 9862
rect 40592 9648 40644 9654
rect 40592 9590 40644 9596
rect 38936 9580 38988 9586
rect 38936 9522 38988 9528
rect 39120 9580 39172 9586
rect 39304 9580 39356 9586
rect 39172 9540 39304 9568
rect 39120 9522 39172 9528
rect 39304 9522 39356 9528
rect 39580 9580 39632 9586
rect 39580 9522 39632 9528
rect 39028 9376 39080 9382
rect 39028 9318 39080 9324
rect 39040 9178 39068 9318
rect 39028 9172 39080 9178
rect 39028 9114 39080 9120
rect 39132 9110 39160 9522
rect 39120 9104 39172 9110
rect 39120 9046 39172 9052
rect 39592 8838 39620 9522
rect 40132 9512 40184 9518
rect 40132 9454 40184 9460
rect 40040 9376 40092 9382
rect 40040 9318 40092 9324
rect 39580 8832 39632 8838
rect 39580 8774 39632 8780
rect 39396 7744 39448 7750
rect 39396 7686 39448 7692
rect 39408 7546 39436 7686
rect 39396 7540 39448 7546
rect 39396 7482 39448 7488
rect 39120 6996 39172 7002
rect 39120 6938 39172 6944
rect 39132 6458 39160 6938
rect 39592 6934 39620 8774
rect 39948 8424 40000 8430
rect 39948 8366 40000 8372
rect 39960 7206 39988 8366
rect 40052 7410 40080 9318
rect 40144 9042 40172 9454
rect 40696 9178 40724 9998
rect 40684 9172 40736 9178
rect 40684 9114 40736 9120
rect 40132 9036 40184 9042
rect 40132 8978 40184 8984
rect 40144 7410 40172 8978
rect 40684 8900 40736 8906
rect 40684 8842 40736 8848
rect 40696 8634 40724 8842
rect 40684 8628 40736 8634
rect 40684 8570 40736 8576
rect 40788 8566 40816 10678
rect 41604 10668 41656 10674
rect 41604 10610 41656 10616
rect 41328 10600 41380 10606
rect 41328 10542 41380 10548
rect 41340 10062 41368 10542
rect 41328 10056 41380 10062
rect 41328 9998 41380 10004
rect 41340 9674 41368 9998
rect 41340 9646 41460 9674
rect 41432 9330 41460 9646
rect 41616 9586 41644 10610
rect 41708 9586 41736 11018
rect 41892 10674 41920 11494
rect 41880 10668 41932 10674
rect 41880 10610 41932 10616
rect 42248 10600 42300 10606
rect 42248 10542 42300 10548
rect 42156 10464 42208 10470
rect 42156 10406 42208 10412
rect 42168 10146 42196 10406
rect 42260 10266 42288 10542
rect 42248 10260 42300 10266
rect 42248 10202 42300 10208
rect 42444 10198 42472 11630
rect 42524 11008 42576 11014
rect 42524 10950 42576 10956
rect 42076 10130 42196 10146
rect 42432 10192 42484 10198
rect 42432 10134 42484 10140
rect 42064 10124 42196 10130
rect 42116 10118 42196 10124
rect 42064 10066 42116 10072
rect 42536 10062 42564 10950
rect 42812 10130 42840 12582
rect 42996 12434 43024 13262
rect 44192 12918 44220 14758
rect 44560 13802 44588 16458
rect 44640 16448 44692 16454
rect 44640 16390 44692 16396
rect 44732 16448 44784 16454
rect 44732 16390 44784 16396
rect 44652 16250 44680 16390
rect 44640 16244 44692 16250
rect 44640 16186 44692 16192
rect 44652 15502 44680 16186
rect 44744 16182 44772 16390
rect 44928 16250 44956 16934
rect 45020 16522 45048 18566
rect 45480 18290 45508 19654
rect 45652 18624 45704 18630
rect 45652 18566 45704 18572
rect 45664 18426 45692 18566
rect 45652 18420 45704 18426
rect 45652 18362 45704 18368
rect 45284 18284 45336 18290
rect 45284 18226 45336 18232
rect 45468 18284 45520 18290
rect 45468 18226 45520 18232
rect 45296 17882 45324 18226
rect 45652 18148 45704 18154
rect 45652 18090 45704 18096
rect 45284 17876 45336 17882
rect 45284 17818 45336 17824
rect 45664 17202 45692 18090
rect 45652 17196 45704 17202
rect 45652 17138 45704 17144
rect 45928 16992 45980 16998
rect 45928 16934 45980 16940
rect 45940 16794 45968 16934
rect 45928 16788 45980 16794
rect 45928 16730 45980 16736
rect 45376 16584 45428 16590
rect 45376 16526 45428 16532
rect 45742 16552 45798 16561
rect 45008 16516 45060 16522
rect 45008 16458 45060 16464
rect 45192 16448 45244 16454
rect 45192 16390 45244 16396
rect 44916 16244 44968 16250
rect 44916 16186 44968 16192
rect 44732 16176 44784 16182
rect 44732 16118 44784 16124
rect 44928 15706 44956 16186
rect 44916 15700 44968 15706
rect 44916 15642 44968 15648
rect 44732 15564 44784 15570
rect 44732 15506 44784 15512
rect 44640 15496 44692 15502
rect 44640 15438 44692 15444
rect 44744 15026 44772 15506
rect 45204 15162 45232 16390
rect 45388 15706 45416 16526
rect 45652 16516 45704 16522
rect 45742 16487 45798 16496
rect 45652 16458 45704 16464
rect 45664 15858 45692 16458
rect 45756 16182 45784 16487
rect 45744 16176 45796 16182
rect 45744 16118 45796 16124
rect 45744 15904 45796 15910
rect 45664 15852 45744 15858
rect 45664 15846 45796 15852
rect 45664 15830 45784 15846
rect 45376 15700 45428 15706
rect 45376 15642 45428 15648
rect 45192 15156 45244 15162
rect 45192 15098 45244 15104
rect 45664 15026 45692 15830
rect 45836 15360 45888 15366
rect 45836 15302 45888 15308
rect 44732 15020 44784 15026
rect 44732 14962 44784 14968
rect 45652 15020 45704 15026
rect 45652 14962 45704 14968
rect 44744 14074 44772 14962
rect 45560 14476 45612 14482
rect 45560 14418 45612 14424
rect 44732 14068 44784 14074
rect 44732 14010 44784 14016
rect 44824 13864 44876 13870
rect 44824 13806 44876 13812
rect 44548 13796 44600 13802
rect 44548 13738 44600 13744
rect 44364 13728 44416 13734
rect 44364 13670 44416 13676
rect 44180 12912 44232 12918
rect 44180 12854 44232 12860
rect 42996 12406 43116 12434
rect 43088 12306 43116 12406
rect 43076 12300 43128 12306
rect 43076 12242 43128 12248
rect 43352 12164 43404 12170
rect 43352 12106 43404 12112
rect 43364 11898 43392 12106
rect 43352 11892 43404 11898
rect 43352 11834 43404 11840
rect 43076 11076 43128 11082
rect 43076 11018 43128 11024
rect 43088 10810 43116 11018
rect 43168 11008 43220 11014
rect 43168 10950 43220 10956
rect 43076 10804 43128 10810
rect 43076 10746 43128 10752
rect 43180 10266 43208 10950
rect 44376 10810 44404 13670
rect 44836 13530 44864 13806
rect 45192 13728 45244 13734
rect 45192 13670 45244 13676
rect 44824 13524 44876 13530
rect 44824 13466 44876 13472
rect 44548 13252 44600 13258
rect 44548 13194 44600 13200
rect 44560 12986 44588 13194
rect 44548 12980 44600 12986
rect 44548 12922 44600 12928
rect 44916 12912 44968 12918
rect 44916 12854 44968 12860
rect 44732 12844 44784 12850
rect 44732 12786 44784 12792
rect 44744 12102 44772 12786
rect 44928 12238 44956 12854
rect 44916 12232 44968 12238
rect 44916 12174 44968 12180
rect 44732 12096 44784 12102
rect 44732 12038 44784 12044
rect 44824 12096 44876 12102
rect 44824 12038 44876 12044
rect 44744 11830 44772 12038
rect 44732 11824 44784 11830
rect 44732 11766 44784 11772
rect 44456 11756 44508 11762
rect 44456 11698 44508 11704
rect 44364 10804 44416 10810
rect 44364 10746 44416 10752
rect 43812 10464 43864 10470
rect 43812 10406 43864 10412
rect 43168 10260 43220 10266
rect 43168 10202 43220 10208
rect 43824 10130 43852 10406
rect 42800 10124 42852 10130
rect 42800 10066 42852 10072
rect 43812 10124 43864 10130
rect 43812 10066 43864 10072
rect 42248 10056 42300 10062
rect 42248 9998 42300 10004
rect 42524 10056 42576 10062
rect 42524 9998 42576 10004
rect 43352 10056 43404 10062
rect 43352 9998 43404 10004
rect 42260 9674 42288 9998
rect 43364 9722 43392 9998
rect 43904 9988 43956 9994
rect 43904 9930 43956 9936
rect 43916 9722 43944 9930
rect 42168 9646 42288 9674
rect 43352 9716 43404 9722
rect 43352 9658 43404 9664
rect 43904 9716 43956 9722
rect 43904 9658 43956 9664
rect 41604 9580 41656 9586
rect 41604 9522 41656 9528
rect 41696 9580 41748 9586
rect 41696 9522 41748 9528
rect 42168 9518 42196 9646
rect 43904 9580 43956 9586
rect 43904 9522 43956 9528
rect 41880 9512 41932 9518
rect 41800 9472 41880 9500
rect 41800 9382 41828 9472
rect 41880 9454 41932 9460
rect 42156 9512 42208 9518
rect 42156 9454 42208 9460
rect 41512 9376 41564 9382
rect 41432 9324 41512 9330
rect 41432 9318 41564 9324
rect 41788 9376 41840 9382
rect 41788 9318 41840 9324
rect 41880 9376 41932 9382
rect 41880 9318 41932 9324
rect 43260 9376 43312 9382
rect 43260 9318 43312 9324
rect 41432 9302 41552 9318
rect 41328 9036 41380 9042
rect 41328 8978 41380 8984
rect 40776 8560 40828 8566
rect 40776 8502 40828 8508
rect 41340 8430 41368 8978
rect 41328 8424 41380 8430
rect 41328 8366 41380 8372
rect 41432 7818 41460 9302
rect 41800 7886 41828 9318
rect 41892 8498 41920 9318
rect 43272 9178 43300 9318
rect 43260 9172 43312 9178
rect 43260 9114 43312 9120
rect 42984 8900 43036 8906
rect 42984 8842 43036 8848
rect 41972 8832 42024 8838
rect 41972 8774 42024 8780
rect 41984 8566 42012 8774
rect 41972 8560 42024 8566
rect 41972 8502 42024 8508
rect 42996 8498 43024 8842
rect 41880 8492 41932 8498
rect 41880 8434 41932 8440
rect 42064 8492 42116 8498
rect 42064 8434 42116 8440
rect 42984 8492 43036 8498
rect 42984 8434 43036 8440
rect 41788 7880 41840 7886
rect 41788 7822 41840 7828
rect 41420 7812 41472 7818
rect 41420 7754 41472 7760
rect 42076 7750 42104 8434
rect 42156 7880 42208 7886
rect 42156 7822 42208 7828
rect 42432 7880 42484 7886
rect 42432 7822 42484 7828
rect 43536 7880 43588 7886
rect 43536 7822 43588 7828
rect 41144 7744 41196 7750
rect 41144 7686 41196 7692
rect 42064 7744 42116 7750
rect 42064 7686 42116 7692
rect 41156 7410 41184 7686
rect 41328 7472 41380 7478
rect 41328 7414 41380 7420
rect 40040 7404 40092 7410
rect 40040 7346 40092 7352
rect 40132 7404 40184 7410
rect 40132 7346 40184 7352
rect 41144 7404 41196 7410
rect 41144 7346 41196 7352
rect 39948 7200 40000 7206
rect 39948 7142 40000 7148
rect 39580 6928 39632 6934
rect 39580 6870 39632 6876
rect 39592 6798 39620 6870
rect 39960 6798 39988 7142
rect 39580 6792 39632 6798
rect 39580 6734 39632 6740
rect 39948 6792 40000 6798
rect 39948 6734 40000 6740
rect 38844 6452 38896 6458
rect 38844 6394 38896 6400
rect 39120 6452 39172 6458
rect 39120 6394 39172 6400
rect 38936 6316 38988 6322
rect 38936 6258 38988 6264
rect 38948 5914 38976 6258
rect 38936 5908 38988 5914
rect 38936 5850 38988 5856
rect 39132 5370 39160 6394
rect 39304 6316 39356 6322
rect 39304 6258 39356 6264
rect 39316 5574 39344 6258
rect 39396 5704 39448 5710
rect 39396 5646 39448 5652
rect 39212 5568 39264 5574
rect 39212 5510 39264 5516
rect 39304 5568 39356 5574
rect 39304 5510 39356 5516
rect 39120 5364 39172 5370
rect 39120 5306 39172 5312
rect 38660 4616 38712 4622
rect 38660 4558 38712 4564
rect 39028 4480 39080 4486
rect 39028 4422 39080 4428
rect 39040 4282 39068 4422
rect 38384 4276 38436 4282
rect 38384 4218 38436 4224
rect 38476 4276 38528 4282
rect 38614 4276 38666 4282
rect 38528 4236 38614 4264
rect 38476 4218 38528 4224
rect 38614 4218 38666 4224
rect 39028 4276 39080 4282
rect 39028 4218 39080 4224
rect 38384 4140 38436 4146
rect 38384 4082 38436 4088
rect 38292 4004 38344 4010
rect 38292 3946 38344 3952
rect 38304 3602 38332 3946
rect 38396 3670 38424 4082
rect 38566 4040 38622 4049
rect 38566 3975 38622 3984
rect 38580 3942 38608 3975
rect 38568 3936 38620 3942
rect 38568 3878 38620 3884
rect 38384 3664 38436 3670
rect 38384 3606 38436 3612
rect 38292 3596 38344 3602
rect 38292 3538 38344 3544
rect 38200 3460 38252 3466
rect 38200 3402 38252 3408
rect 38304 3194 38332 3538
rect 38292 3188 38344 3194
rect 38292 3130 38344 3136
rect 37648 3120 37700 3126
rect 37648 3062 37700 3068
rect 37660 2990 37688 3062
rect 39040 3058 39068 4218
rect 39224 4078 39252 5510
rect 39212 4072 39264 4078
rect 39212 4014 39264 4020
rect 39316 3534 39344 5510
rect 39408 4758 39436 5646
rect 39592 5234 39620 6734
rect 40224 6656 40276 6662
rect 40224 6598 40276 6604
rect 40592 6656 40644 6662
rect 40592 6598 40644 6604
rect 40236 5710 40264 6598
rect 40604 6322 40632 6598
rect 40408 6316 40460 6322
rect 40408 6258 40460 6264
rect 40592 6316 40644 6322
rect 40592 6258 40644 6264
rect 40420 5778 40448 6258
rect 41236 6248 41288 6254
rect 41236 6190 41288 6196
rect 40868 6112 40920 6118
rect 40868 6054 40920 6060
rect 40880 5914 40908 6054
rect 40500 5908 40552 5914
rect 40500 5850 40552 5856
rect 40868 5908 40920 5914
rect 40868 5850 40920 5856
rect 40408 5772 40460 5778
rect 40408 5714 40460 5720
rect 40224 5704 40276 5710
rect 40276 5664 40356 5692
rect 40224 5646 40276 5652
rect 39672 5568 39724 5574
rect 39672 5510 39724 5516
rect 39488 5228 39540 5234
rect 39488 5170 39540 5176
rect 39580 5228 39632 5234
rect 39580 5170 39632 5176
rect 39500 4826 39528 5170
rect 39488 4820 39540 4826
rect 39488 4762 39540 4768
rect 39396 4752 39448 4758
rect 39396 4694 39448 4700
rect 39408 4282 39436 4694
rect 39592 4690 39620 5170
rect 39684 5030 39712 5510
rect 40328 5030 40356 5664
rect 40512 5370 40540 5850
rect 41248 5846 41276 6190
rect 41236 5840 41288 5846
rect 41236 5782 41288 5788
rect 40684 5636 40736 5642
rect 40684 5578 40736 5584
rect 41144 5636 41196 5642
rect 41144 5578 41196 5584
rect 40696 5370 40724 5578
rect 40960 5568 41012 5574
rect 40960 5510 41012 5516
rect 40500 5364 40552 5370
rect 40500 5306 40552 5312
rect 40684 5364 40736 5370
rect 40684 5306 40736 5312
rect 40972 5234 41000 5510
rect 40960 5228 41012 5234
rect 40960 5170 41012 5176
rect 41156 5166 41184 5578
rect 41248 5234 41276 5782
rect 41340 5778 41368 7414
rect 42076 6934 42104 7686
rect 42064 6928 42116 6934
rect 42064 6870 42116 6876
rect 42168 6798 42196 7822
rect 42444 7546 42472 7822
rect 42800 7744 42852 7750
rect 42800 7686 42852 7692
rect 42432 7540 42484 7546
rect 42432 7482 42484 7488
rect 42432 7404 42484 7410
rect 42432 7346 42484 7352
rect 42524 7404 42576 7410
rect 42524 7346 42576 7352
rect 42444 6866 42472 7346
rect 42536 7002 42564 7346
rect 42524 6996 42576 7002
rect 42524 6938 42576 6944
rect 42432 6860 42484 6866
rect 42432 6802 42484 6808
rect 42812 6798 42840 7686
rect 43548 7546 43576 7822
rect 43536 7540 43588 7546
rect 43536 7482 43588 7488
rect 42156 6792 42208 6798
rect 42156 6734 42208 6740
rect 42800 6792 42852 6798
rect 42800 6734 42852 6740
rect 41512 6452 41564 6458
rect 41512 6394 41564 6400
rect 41420 6248 41472 6254
rect 41420 6190 41472 6196
rect 41328 5772 41380 5778
rect 41328 5714 41380 5720
rect 41236 5228 41288 5234
rect 41236 5170 41288 5176
rect 41144 5160 41196 5166
rect 41144 5102 41196 5108
rect 39672 5024 39724 5030
rect 39672 4966 39724 4972
rect 40316 5024 40368 5030
rect 40316 4966 40368 4972
rect 40776 5024 40828 5030
rect 40776 4966 40828 4972
rect 39580 4684 39632 4690
rect 39580 4626 39632 4632
rect 39396 4276 39448 4282
rect 39396 4218 39448 4224
rect 39396 4140 39448 4146
rect 39396 4082 39448 4088
rect 39408 3738 39436 4082
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 39316 3058 39344 3470
rect 39396 3392 39448 3398
rect 39396 3334 39448 3340
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 39028 3052 39080 3058
rect 39028 2994 39080 3000
rect 39304 3052 39356 3058
rect 39304 2994 39356 3000
rect 37556 2984 37608 2990
rect 37556 2926 37608 2932
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 38672 2650 38700 2994
rect 39120 2848 39172 2854
rect 39172 2796 39252 2802
rect 39120 2790 39252 2796
rect 39132 2774 39252 2790
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 38292 2440 38344 2446
rect 38292 2382 38344 2388
rect 38028 870 38148 898
rect 38028 800 38056 870
rect 35544 734 35848 762
rect 38014 0 38070 800
rect 38120 762 38148 870
rect 38304 762 38332 2382
rect 39224 2378 39252 2774
rect 39408 2446 39436 3334
rect 39684 2514 39712 4966
rect 40040 4548 40092 4554
rect 40040 4490 40092 4496
rect 40132 4548 40184 4554
rect 40132 4490 40184 4496
rect 39948 4072 40000 4078
rect 39948 4014 40000 4020
rect 39960 3738 39988 4014
rect 40052 3942 40080 4490
rect 40144 4214 40172 4490
rect 40224 4480 40276 4486
rect 40224 4422 40276 4428
rect 40236 4282 40264 4422
rect 40224 4276 40276 4282
rect 40224 4218 40276 4224
rect 40328 4214 40356 4966
rect 40788 4826 40816 4966
rect 40776 4820 40828 4826
rect 40776 4762 40828 4768
rect 40500 4616 40552 4622
rect 40500 4558 40552 4564
rect 40408 4480 40460 4486
rect 40408 4422 40460 4428
rect 40132 4208 40184 4214
rect 40132 4150 40184 4156
rect 40316 4208 40368 4214
rect 40316 4150 40368 4156
rect 40040 3936 40092 3942
rect 40040 3878 40092 3884
rect 40052 3754 40080 3878
rect 39948 3732 40000 3738
rect 40052 3726 40172 3754
rect 39948 3674 40000 3680
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 40052 3126 40080 3538
rect 40040 3120 40092 3126
rect 40040 3062 40092 3068
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 39960 2650 39988 2926
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 39672 2508 39724 2514
rect 39672 2450 39724 2456
rect 40144 2446 40172 3726
rect 40420 3466 40448 4422
rect 40512 4214 40540 4558
rect 41340 4554 41368 5714
rect 41432 5574 41460 6190
rect 41420 5568 41472 5574
rect 41420 5510 41472 5516
rect 41524 5234 41552 6394
rect 43916 6390 43944 9522
rect 44272 9512 44324 9518
rect 44272 9454 44324 9460
rect 44284 9042 44312 9454
rect 44468 9382 44496 11698
rect 44836 11694 44864 12038
rect 44916 11756 44968 11762
rect 44916 11698 44968 11704
rect 44824 11688 44876 11694
rect 44824 11630 44876 11636
rect 44928 10810 44956 11698
rect 45100 11688 45152 11694
rect 45100 11630 45152 11636
rect 44916 10804 44968 10810
rect 44916 10746 44968 10752
rect 44640 10464 44692 10470
rect 44640 10406 44692 10412
rect 44652 10305 44680 10406
rect 44638 10296 44694 10305
rect 44928 10266 44956 10746
rect 45112 10606 45140 11630
rect 45204 10810 45232 13670
rect 45572 11218 45600 14418
rect 45664 14074 45692 14962
rect 45848 14278 45876 15302
rect 45836 14272 45888 14278
rect 45836 14214 45888 14220
rect 45652 14068 45704 14074
rect 45652 14010 45704 14016
rect 45744 13252 45796 13258
rect 45744 13194 45796 13200
rect 45756 12986 45784 13194
rect 45744 12980 45796 12986
rect 45744 12922 45796 12928
rect 45848 12850 45876 14214
rect 45836 12844 45888 12850
rect 45836 12786 45888 12792
rect 46032 11218 46060 19858
rect 46124 18970 46152 20402
rect 46216 19242 46244 20810
rect 46584 20806 46612 21082
rect 46664 20936 46716 20942
rect 46664 20878 46716 20884
rect 46572 20800 46624 20806
rect 46572 20742 46624 20748
rect 46480 20460 46532 20466
rect 46480 20402 46532 20408
rect 46492 19786 46520 20402
rect 46676 20058 46704 20878
rect 46756 20596 46808 20602
rect 46756 20538 46808 20544
rect 46664 20052 46716 20058
rect 46664 19994 46716 20000
rect 46664 19848 46716 19854
rect 46664 19790 46716 19796
rect 46480 19780 46532 19786
rect 46480 19722 46532 19728
rect 46388 19712 46440 19718
rect 46388 19654 46440 19660
rect 46400 19310 46428 19654
rect 46676 19514 46704 19790
rect 46664 19508 46716 19514
rect 46664 19450 46716 19456
rect 46388 19304 46440 19310
rect 46388 19246 46440 19252
rect 46572 19304 46624 19310
rect 46572 19246 46624 19252
rect 46204 19236 46256 19242
rect 46204 19178 46256 19184
rect 46400 18970 46428 19246
rect 46112 18964 46164 18970
rect 46112 18906 46164 18912
rect 46388 18964 46440 18970
rect 46388 18906 46440 18912
rect 46480 18624 46532 18630
rect 46480 18566 46532 18572
rect 46492 18290 46520 18566
rect 46584 18426 46612 19246
rect 46664 18896 46716 18902
rect 46664 18838 46716 18844
rect 46572 18420 46624 18426
rect 46572 18362 46624 18368
rect 46676 18290 46704 18838
rect 46768 18766 46796 20538
rect 46860 19378 46888 21508
rect 47032 21490 47084 21496
rect 47320 21146 47348 21558
rect 47504 21350 47532 21966
rect 47492 21344 47544 21350
rect 47492 21286 47544 21292
rect 47308 21140 47360 21146
rect 47308 21082 47360 21088
rect 47596 21010 47624 22510
rect 47964 22234 47992 22986
rect 47952 22228 48004 22234
rect 47952 22170 48004 22176
rect 47676 22024 47728 22030
rect 47674 21992 47676 22001
rect 47728 21992 47730 22001
rect 47674 21927 47730 21936
rect 47860 21888 47912 21894
rect 47860 21830 47912 21836
rect 47872 21690 47900 21830
rect 47860 21684 47912 21690
rect 47860 21626 47912 21632
rect 48056 21570 48084 23122
rect 49516 23112 49568 23118
rect 49516 23054 49568 23060
rect 49424 22976 49476 22982
rect 49424 22918 49476 22924
rect 49436 22642 49464 22918
rect 48872 22636 48924 22642
rect 48872 22578 48924 22584
rect 49424 22636 49476 22642
rect 49424 22578 49476 22584
rect 48320 22432 48372 22438
rect 48240 22392 48320 22420
rect 48136 22228 48188 22234
rect 48136 22170 48188 22176
rect 48148 21962 48176 22170
rect 48240 22030 48268 22392
rect 48320 22374 48372 22380
rect 48320 22160 48372 22166
rect 48320 22102 48372 22108
rect 48332 22030 48360 22102
rect 48884 22098 48912 22578
rect 48872 22092 48924 22098
rect 48872 22034 48924 22040
rect 48964 22092 49016 22098
rect 49528 22094 49556 23054
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 49528 22066 49648 22094
rect 48964 22034 49016 22040
rect 48228 22024 48280 22030
rect 48228 21966 48280 21972
rect 48320 22024 48372 22030
rect 48320 21966 48372 21972
rect 48410 21992 48466 22001
rect 48136 21956 48188 21962
rect 48410 21927 48412 21936
rect 48136 21898 48188 21904
rect 48464 21927 48466 21936
rect 48412 21898 48464 21904
rect 48596 21888 48648 21894
rect 48596 21830 48648 21836
rect 48608 21690 48636 21830
rect 48596 21684 48648 21690
rect 48596 21626 48648 21632
rect 47768 21548 47820 21554
rect 48056 21542 48268 21570
rect 47768 21490 47820 21496
rect 47584 21004 47636 21010
rect 47584 20946 47636 20952
rect 47780 20806 47808 21490
rect 48240 21486 48268 21542
rect 48228 21480 48280 21486
rect 48884 21434 48912 22034
rect 48976 21554 49004 22034
rect 49620 22030 49648 22066
rect 49608 22024 49660 22030
rect 49608 21966 49660 21972
rect 49700 22024 49752 22030
rect 49700 21966 49752 21972
rect 49240 21888 49292 21894
rect 49240 21830 49292 21836
rect 49252 21690 49280 21830
rect 49240 21684 49292 21690
rect 49240 21626 49292 21632
rect 48964 21548 49016 21554
rect 48964 21490 49016 21496
rect 48228 21422 48280 21428
rect 48792 21406 48912 21434
rect 48792 21146 48820 21406
rect 48872 21344 48924 21350
rect 48872 21286 48924 21292
rect 48320 21140 48372 21146
rect 48320 21082 48372 21088
rect 48780 21140 48832 21146
rect 48780 21082 48832 21088
rect 46940 20800 46992 20806
rect 46940 20742 46992 20748
rect 47768 20800 47820 20806
rect 47768 20742 47820 20748
rect 47860 20800 47912 20806
rect 47860 20742 47912 20748
rect 46952 20262 46980 20742
rect 47308 20528 47360 20534
rect 47308 20470 47360 20476
rect 46940 20256 46992 20262
rect 46940 20198 46992 20204
rect 47032 20256 47084 20262
rect 47032 20198 47084 20204
rect 47044 19854 47072 20198
rect 47032 19848 47084 19854
rect 47032 19790 47084 19796
rect 47124 19848 47176 19854
rect 47124 19790 47176 19796
rect 47032 19508 47084 19514
rect 47032 19450 47084 19456
rect 46848 19372 46900 19378
rect 46848 19314 46900 19320
rect 46940 19372 46992 19378
rect 46940 19314 46992 19320
rect 46756 18760 46808 18766
rect 46756 18702 46808 18708
rect 46952 18601 46980 19314
rect 46754 18592 46810 18601
rect 46754 18527 46810 18536
rect 46938 18592 46994 18601
rect 46938 18527 46994 18536
rect 46768 18290 46796 18527
rect 46848 18352 46900 18358
rect 46848 18294 46900 18300
rect 46938 18320 46994 18329
rect 46480 18284 46532 18290
rect 46480 18226 46532 18232
rect 46664 18284 46716 18290
rect 46664 18226 46716 18232
rect 46756 18284 46808 18290
rect 46756 18226 46808 18232
rect 46388 18080 46440 18086
rect 46388 18022 46440 18028
rect 46400 17610 46428 18022
rect 46480 17876 46532 17882
rect 46480 17818 46532 17824
rect 46388 17604 46440 17610
rect 46388 17546 46440 17552
rect 46492 17338 46520 17818
rect 46676 17678 46704 18226
rect 46860 17882 46888 18294
rect 46938 18255 46994 18264
rect 46952 18086 46980 18255
rect 46940 18080 46992 18086
rect 46940 18022 46992 18028
rect 46848 17876 46900 17882
rect 46848 17818 46900 17824
rect 46952 17678 46980 18022
rect 46664 17672 46716 17678
rect 46664 17614 46716 17620
rect 46756 17672 46808 17678
rect 46756 17614 46808 17620
rect 46940 17672 46992 17678
rect 46940 17614 46992 17620
rect 46480 17332 46532 17338
rect 46480 17274 46532 17280
rect 46388 17196 46440 17202
rect 46388 17138 46440 17144
rect 46204 16992 46256 16998
rect 46204 16934 46256 16940
rect 46216 16794 46244 16934
rect 46204 16788 46256 16794
rect 46204 16730 46256 16736
rect 46400 16096 46428 17138
rect 46572 17060 46624 17066
rect 46572 17002 46624 17008
rect 46584 16114 46612 17002
rect 46676 16658 46704 17614
rect 46664 16652 46716 16658
rect 46664 16594 46716 16600
rect 46768 16590 46796 17614
rect 47044 17338 47072 19450
rect 47136 18408 47164 19790
rect 47320 19514 47348 20470
rect 47768 20460 47820 20466
rect 47768 20402 47820 20408
rect 47492 20256 47544 20262
rect 47492 20198 47544 20204
rect 47504 19990 47532 20198
rect 47492 19984 47544 19990
rect 47492 19926 47544 19932
rect 47400 19780 47452 19786
rect 47452 19740 47624 19768
rect 47400 19722 47452 19728
rect 47308 19508 47360 19514
rect 47308 19450 47360 19456
rect 47320 19378 47348 19450
rect 47308 19372 47360 19378
rect 47308 19314 47360 19320
rect 47216 19168 47268 19174
rect 47216 19110 47268 19116
rect 47400 19168 47452 19174
rect 47400 19110 47452 19116
rect 47228 18970 47256 19110
rect 47216 18964 47268 18970
rect 47216 18906 47268 18912
rect 47412 18426 47440 19110
rect 47596 18426 47624 19740
rect 47780 19378 47808 20402
rect 47872 20330 47900 20742
rect 48332 20466 48360 21082
rect 48884 21010 48912 21286
rect 48976 21146 49004 21490
rect 49332 21480 49384 21486
rect 49332 21422 49384 21428
rect 49344 21146 49372 21422
rect 48964 21140 49016 21146
rect 48964 21082 49016 21088
rect 49332 21140 49384 21146
rect 49332 21082 49384 21088
rect 49712 21010 49740 21966
rect 49792 21888 49844 21894
rect 49792 21830 49844 21836
rect 49804 21622 49832 21830
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 49792 21616 49844 21622
rect 49792 21558 49844 21564
rect 68204 21457 68232 60658
rect 68374 60616 68430 60625
rect 68374 60551 68376 60560
rect 68428 60551 68430 60560
rect 68376 60522 68428 60528
rect 68468 57928 68520 57934
rect 68466 57896 68468 57905
rect 68520 57896 68522 57905
rect 68466 57831 68522 57840
rect 68466 55176 68522 55185
rect 68466 55111 68468 55120
rect 68520 55111 68522 55120
rect 68468 55082 68520 55088
rect 68468 52488 68520 52494
rect 68466 52456 68468 52465
rect 68520 52456 68522 52465
rect 68466 52391 68522 52400
rect 68468 49768 68520 49774
rect 68466 49736 68468 49745
rect 68520 49736 68522 49745
rect 68466 49671 68522 49680
rect 68468 47048 68520 47054
rect 68466 47016 68468 47025
rect 68520 47016 68522 47025
rect 68466 46951 68522 46960
rect 68466 44296 68522 44305
rect 68466 44231 68468 44240
rect 68520 44231 68522 44240
rect 68468 44202 68520 44208
rect 68468 41608 68520 41614
rect 68466 41576 68468 41585
rect 68520 41576 68522 41585
rect 68466 41511 68522 41520
rect 68468 36168 68520 36174
rect 68466 36136 68468 36145
rect 68520 36136 68522 36145
rect 68466 36071 68522 36080
rect 68744 33516 68796 33522
rect 68744 33458 68796 33464
rect 68756 33425 68784 33458
rect 68742 33416 68798 33425
rect 68742 33351 68798 33360
rect 68376 33312 68428 33318
rect 68376 33254 68428 33260
rect 68388 21593 68416 33254
rect 68468 30728 68520 30734
rect 68466 30696 68468 30705
rect 68520 30696 68522 30705
rect 68466 30631 68522 30640
rect 68466 27976 68522 27985
rect 68466 27911 68468 27920
rect 68520 27911 68522 27920
rect 68468 27882 68520 27888
rect 68468 25288 68520 25294
rect 68466 25256 68468 25265
rect 68520 25256 68522 25265
rect 68466 25191 68522 25200
rect 68466 22536 68522 22545
rect 68466 22471 68468 22480
rect 68520 22471 68522 22480
rect 68468 22442 68520 22448
rect 68374 21584 68430 21593
rect 68374 21519 68430 21528
rect 68190 21448 68246 21457
rect 68190 21383 68246 21392
rect 50068 21344 50120 21350
rect 50068 21286 50120 21292
rect 50712 21344 50764 21350
rect 50712 21286 50764 21292
rect 50804 21344 50856 21350
rect 50804 21286 50856 21292
rect 48872 21004 48924 21010
rect 48872 20946 48924 20952
rect 49700 21004 49752 21010
rect 49700 20946 49752 20952
rect 48596 20868 48648 20874
rect 48596 20810 48648 20816
rect 48504 20800 48556 20806
rect 48504 20742 48556 20748
rect 48320 20460 48372 20466
rect 48320 20402 48372 20408
rect 47860 20324 47912 20330
rect 47860 20266 47912 20272
rect 47952 20256 48004 20262
rect 47952 20198 48004 20204
rect 47964 19922 47992 20198
rect 48332 19990 48360 20402
rect 48516 20398 48544 20742
rect 48504 20392 48556 20398
rect 48504 20334 48556 20340
rect 48516 20058 48544 20334
rect 48608 20262 48636 20810
rect 48872 20800 48924 20806
rect 48872 20742 48924 20748
rect 49148 20800 49200 20806
rect 49148 20742 49200 20748
rect 48884 20482 48912 20742
rect 49160 20602 49188 20742
rect 49148 20596 49200 20602
rect 49148 20538 49200 20544
rect 48792 20454 48912 20482
rect 49160 20466 49188 20538
rect 49148 20460 49200 20466
rect 48792 20398 48820 20454
rect 49148 20402 49200 20408
rect 48780 20392 48832 20398
rect 48780 20334 48832 20340
rect 48596 20256 48648 20262
rect 48596 20198 48648 20204
rect 48504 20052 48556 20058
rect 48504 19994 48556 20000
rect 48320 19984 48372 19990
rect 48320 19926 48372 19932
rect 47952 19916 48004 19922
rect 47952 19858 48004 19864
rect 48792 19446 48820 20334
rect 49608 20256 49660 20262
rect 49608 20198 49660 20204
rect 49620 19854 49648 20198
rect 49608 19848 49660 19854
rect 49608 19790 49660 19796
rect 49712 19786 49740 20946
rect 49792 20868 49844 20874
rect 49792 20810 49844 20816
rect 49884 20868 49936 20874
rect 49884 20810 49936 20816
rect 49976 20868 50028 20874
rect 49976 20810 50028 20816
rect 49804 19786 49832 20810
rect 49896 20466 49924 20810
rect 49988 20602 50016 20810
rect 49976 20596 50028 20602
rect 49976 20538 50028 20544
rect 49884 20460 49936 20466
rect 49884 20402 49936 20408
rect 49988 20058 50016 20538
rect 49976 20052 50028 20058
rect 49976 19994 50028 20000
rect 49988 19854 50016 19994
rect 50080 19854 50108 21286
rect 50724 21010 50752 21286
rect 50816 21078 50844 21286
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 50804 21072 50856 21078
rect 50804 21014 50856 21020
rect 50712 21004 50764 21010
rect 50712 20946 50764 20952
rect 50436 20936 50488 20942
rect 50172 20884 50436 20890
rect 50172 20878 50488 20884
rect 50172 20862 50476 20878
rect 50172 20534 50200 20862
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50160 20528 50212 20534
rect 50160 20470 50212 20476
rect 50804 20460 50856 20466
rect 50804 20402 50856 20408
rect 50528 20052 50580 20058
rect 50528 19994 50580 20000
rect 50540 19922 50568 19994
rect 50528 19916 50580 19922
rect 50528 19858 50580 19864
rect 49976 19848 50028 19854
rect 49976 19790 50028 19796
rect 50068 19848 50120 19854
rect 50068 19790 50120 19796
rect 49700 19780 49752 19786
rect 49700 19722 49752 19728
rect 49792 19780 49844 19786
rect 49792 19722 49844 19728
rect 48780 19440 48832 19446
rect 48780 19382 48832 19388
rect 47768 19372 47820 19378
rect 47768 19314 47820 19320
rect 47676 18692 47728 18698
rect 47676 18634 47728 18640
rect 47400 18420 47452 18426
rect 47136 18380 47256 18408
rect 47122 18320 47178 18329
rect 47122 18255 47178 18264
rect 47136 18222 47164 18255
rect 47124 18216 47176 18222
rect 47124 18158 47176 18164
rect 47032 17332 47084 17338
rect 47032 17274 47084 17280
rect 46756 16584 46808 16590
rect 46756 16526 46808 16532
rect 46480 16108 46532 16114
rect 46400 16068 46480 16096
rect 46480 16050 46532 16056
rect 46572 16108 46624 16114
rect 46572 16050 46624 16056
rect 46296 15904 46348 15910
rect 46296 15846 46348 15852
rect 46308 15706 46336 15846
rect 46296 15700 46348 15706
rect 46296 15642 46348 15648
rect 46492 15473 46520 16050
rect 46768 15706 46796 16526
rect 46756 15700 46808 15706
rect 46756 15642 46808 15648
rect 46478 15464 46534 15473
rect 46478 15399 46534 15408
rect 46492 14482 46520 15399
rect 46768 15026 46796 15642
rect 46572 15020 46624 15026
rect 46572 14962 46624 14968
rect 46756 15020 46808 15026
rect 46756 14962 46808 14968
rect 46584 14618 46612 14962
rect 47228 14618 47256 18380
rect 47400 18362 47452 18368
rect 47584 18420 47636 18426
rect 47584 18362 47636 18368
rect 47596 18290 47624 18362
rect 47584 18284 47636 18290
rect 47584 18226 47636 18232
rect 47596 17746 47624 18226
rect 47688 18086 47716 18634
rect 47780 18358 47808 19314
rect 47952 19168 48004 19174
rect 47952 19110 48004 19116
rect 47768 18352 47820 18358
rect 47964 18329 47992 19110
rect 49712 18766 49740 19722
rect 49804 19378 49832 19722
rect 49988 19378 50016 19790
rect 49792 19372 49844 19378
rect 49792 19314 49844 19320
rect 49976 19372 50028 19378
rect 49976 19314 50028 19320
rect 48872 18760 48924 18766
rect 48872 18702 48924 18708
rect 49700 18760 49752 18766
rect 49700 18702 49752 18708
rect 48228 18692 48280 18698
rect 48228 18634 48280 18640
rect 47768 18294 47820 18300
rect 47950 18320 48006 18329
rect 47780 18170 47808 18294
rect 47950 18255 48006 18264
rect 47952 18216 48004 18222
rect 47780 18164 47952 18170
rect 47780 18158 48004 18164
rect 47780 18142 47992 18158
rect 47676 18080 47728 18086
rect 47676 18022 47728 18028
rect 47584 17740 47636 17746
rect 47584 17682 47636 17688
rect 48240 17134 48268 18634
rect 48780 18624 48832 18630
rect 48778 18592 48780 18601
rect 48832 18592 48834 18601
rect 48778 18527 48834 18536
rect 48884 18222 48912 18702
rect 48964 18624 49016 18630
rect 48964 18566 49016 18572
rect 48976 18290 49004 18566
rect 50080 18426 50108 19790
rect 50160 19712 50212 19718
rect 50160 19654 50212 19660
rect 50620 19712 50672 19718
rect 50620 19654 50672 19660
rect 50172 19514 50200 19654
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50160 19508 50212 19514
rect 50160 19450 50212 19456
rect 50632 18834 50660 19654
rect 50816 19310 50844 20402
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 68468 19848 68520 19854
rect 68466 19816 68468 19825
rect 68520 19816 68522 19825
rect 51080 19780 51132 19786
rect 68466 19751 68522 19760
rect 51080 19722 51132 19728
rect 50804 19304 50856 19310
rect 50804 19246 50856 19252
rect 50816 18970 50844 19246
rect 51092 18970 51120 19722
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 50804 18964 50856 18970
rect 50804 18906 50856 18912
rect 51080 18964 51132 18970
rect 51080 18906 51132 18912
rect 50816 18834 50844 18906
rect 50620 18828 50672 18834
rect 50620 18770 50672 18776
rect 50804 18828 50856 18834
rect 50804 18770 50856 18776
rect 50160 18624 50212 18630
rect 50160 18566 50212 18572
rect 50712 18624 50764 18630
rect 50712 18566 50764 18572
rect 50068 18420 50120 18426
rect 50068 18362 50120 18368
rect 48964 18284 49016 18290
rect 48964 18226 49016 18232
rect 48872 18216 48924 18222
rect 48872 18158 48924 18164
rect 49976 18216 50028 18222
rect 49976 18158 50028 18164
rect 49988 17882 50016 18158
rect 49976 17876 50028 17882
rect 49976 17818 50028 17824
rect 49240 17740 49292 17746
rect 49240 17682 49292 17688
rect 48412 17536 48464 17542
rect 48412 17478 48464 17484
rect 48780 17536 48832 17542
rect 48780 17478 48832 17484
rect 48872 17536 48924 17542
rect 48872 17478 48924 17484
rect 47308 17128 47360 17134
rect 47308 17070 47360 17076
rect 48228 17128 48280 17134
rect 48228 17070 48280 17076
rect 46572 14612 46624 14618
rect 46572 14554 46624 14560
rect 47216 14612 47268 14618
rect 47216 14554 47268 14560
rect 47320 14550 47348 17070
rect 48240 15910 48268 17070
rect 48424 16590 48452 17478
rect 48504 17128 48556 17134
rect 48504 17070 48556 17076
rect 48516 16794 48544 17070
rect 48792 16794 48820 17478
rect 48504 16788 48556 16794
rect 48504 16730 48556 16736
rect 48780 16788 48832 16794
rect 48780 16730 48832 16736
rect 48780 16652 48832 16658
rect 48780 16594 48832 16600
rect 48412 16584 48464 16590
rect 48412 16526 48464 16532
rect 48504 16108 48556 16114
rect 48504 16050 48556 16056
rect 48228 15904 48280 15910
rect 48228 15846 48280 15852
rect 48240 15706 48268 15846
rect 48228 15700 48280 15706
rect 48228 15642 48280 15648
rect 47400 15496 47452 15502
rect 47400 15438 47452 15444
rect 47412 14550 47440 15438
rect 48516 15366 48544 16050
rect 48504 15360 48556 15366
rect 48504 15302 48556 15308
rect 47584 14952 47636 14958
rect 47584 14894 47636 14900
rect 47492 14816 47544 14822
rect 47492 14758 47544 14764
rect 47504 14618 47532 14758
rect 47596 14618 47624 14894
rect 48320 14816 48372 14822
rect 48320 14758 48372 14764
rect 47492 14612 47544 14618
rect 47492 14554 47544 14560
rect 47584 14612 47636 14618
rect 47584 14554 47636 14560
rect 47308 14544 47360 14550
rect 47308 14486 47360 14492
rect 47400 14544 47452 14550
rect 47400 14486 47452 14492
rect 46480 14476 46532 14482
rect 46480 14418 46532 14424
rect 46756 14476 46808 14482
rect 46756 14418 46808 14424
rect 46388 13728 46440 13734
rect 46388 13670 46440 13676
rect 46480 13728 46532 13734
rect 46480 13670 46532 13676
rect 46112 13388 46164 13394
rect 46112 13330 46164 13336
rect 46124 12714 46152 13330
rect 46400 12782 46428 13670
rect 46492 12850 46520 13670
rect 46768 13326 46796 14418
rect 48228 14272 48280 14278
rect 48228 14214 48280 14220
rect 47216 13932 47268 13938
rect 47216 13874 47268 13880
rect 47032 13728 47084 13734
rect 47032 13670 47084 13676
rect 46756 13320 46808 13326
rect 46756 13262 46808 13268
rect 46480 12844 46532 12850
rect 46480 12786 46532 12792
rect 46388 12776 46440 12782
rect 46388 12718 46440 12724
rect 46112 12708 46164 12714
rect 46112 12650 46164 12656
rect 46124 12306 46152 12650
rect 46112 12300 46164 12306
rect 46112 12242 46164 12248
rect 46124 11762 46152 12242
rect 46112 11756 46164 11762
rect 46112 11698 46164 11704
rect 47044 11286 47072 13670
rect 47228 13462 47256 13874
rect 48136 13864 48188 13870
rect 48136 13806 48188 13812
rect 47952 13728 48004 13734
rect 47952 13670 48004 13676
rect 47964 13462 47992 13670
rect 48148 13462 48176 13806
rect 48240 13530 48268 14214
rect 48228 13524 48280 13530
rect 48228 13466 48280 13472
rect 47216 13456 47268 13462
rect 47216 13398 47268 13404
rect 47952 13456 48004 13462
rect 47952 13398 48004 13404
rect 48136 13456 48188 13462
rect 48136 13398 48188 13404
rect 47964 13326 47992 13398
rect 47952 13320 48004 13326
rect 47952 13262 48004 13268
rect 48228 13320 48280 13326
rect 48228 13262 48280 13268
rect 47308 13184 47360 13190
rect 47308 13126 47360 13132
rect 47320 12434 47348 13126
rect 48240 12986 48268 13262
rect 48332 13258 48360 14758
rect 48412 13932 48464 13938
rect 48412 13874 48464 13880
rect 48320 13252 48372 13258
rect 48320 13194 48372 13200
rect 48228 12980 48280 12986
rect 48228 12922 48280 12928
rect 48228 12776 48280 12782
rect 48228 12718 48280 12724
rect 48240 12442 48268 12718
rect 47136 12406 47348 12434
rect 48228 12436 48280 12442
rect 47136 12306 47164 12406
rect 48228 12378 48280 12384
rect 47124 12300 47176 12306
rect 47124 12242 47176 12248
rect 47124 12164 47176 12170
rect 47124 12106 47176 12112
rect 47136 11898 47164 12106
rect 47124 11892 47176 11898
rect 47124 11834 47176 11840
rect 47768 11824 47820 11830
rect 47768 11766 47820 11772
rect 47216 11756 47268 11762
rect 47216 11698 47268 11704
rect 47032 11280 47084 11286
rect 47032 11222 47084 11228
rect 45560 11212 45612 11218
rect 45560 11154 45612 11160
rect 46020 11212 46072 11218
rect 46020 11154 46072 11160
rect 45192 10804 45244 10810
rect 45192 10746 45244 10752
rect 45572 10606 45600 11154
rect 46388 11144 46440 11150
rect 46388 11086 46440 11092
rect 45836 11076 45888 11082
rect 45836 11018 45888 11024
rect 45100 10600 45152 10606
rect 45100 10542 45152 10548
rect 45560 10600 45612 10606
rect 45560 10542 45612 10548
rect 44638 10231 44694 10240
rect 44916 10260 44968 10266
rect 44916 10202 44968 10208
rect 45112 9586 45140 10542
rect 45572 10266 45600 10542
rect 45560 10260 45612 10266
rect 45560 10202 45612 10208
rect 45560 10124 45612 10130
rect 45560 10066 45612 10072
rect 45572 9654 45600 10066
rect 45560 9648 45612 9654
rect 45560 9590 45612 9596
rect 45100 9580 45152 9586
rect 45100 9522 45152 9528
rect 44456 9376 44508 9382
rect 44456 9318 44508 9324
rect 44272 9036 44324 9042
rect 44272 8978 44324 8984
rect 45112 8974 45140 9522
rect 45652 9512 45704 9518
rect 45652 9454 45704 9460
rect 45468 9444 45520 9450
rect 45468 9386 45520 9392
rect 45192 9376 45244 9382
rect 45192 9318 45244 9324
rect 45204 8974 45232 9318
rect 45100 8968 45152 8974
rect 45100 8910 45152 8916
rect 45192 8968 45244 8974
rect 45192 8910 45244 8916
rect 45376 8832 45428 8838
rect 45376 8774 45428 8780
rect 44732 8492 44784 8498
rect 44732 8434 44784 8440
rect 44744 8294 44772 8434
rect 44732 8288 44784 8294
rect 44732 8230 44784 8236
rect 45388 7449 45416 8774
rect 45480 8498 45508 9386
rect 45664 9042 45692 9454
rect 45652 9036 45704 9042
rect 45652 8978 45704 8984
rect 45560 8968 45612 8974
rect 45560 8910 45612 8916
rect 45468 8492 45520 8498
rect 45468 8434 45520 8440
rect 45572 8362 45600 8910
rect 45744 8492 45796 8498
rect 45744 8434 45796 8440
rect 45560 8356 45612 8362
rect 45560 8298 45612 8304
rect 45756 8090 45784 8434
rect 45848 8090 45876 11018
rect 46400 10266 46428 11086
rect 47228 11082 47256 11698
rect 47584 11688 47636 11694
rect 47584 11630 47636 11636
rect 47216 11076 47268 11082
rect 47216 11018 47268 11024
rect 46388 10260 46440 10266
rect 46388 10202 46440 10208
rect 46020 10056 46072 10062
rect 46020 9998 46072 10004
rect 45928 9920 45980 9926
rect 45928 9862 45980 9868
rect 45744 8084 45796 8090
rect 45744 8026 45796 8032
rect 45836 8084 45888 8090
rect 45836 8026 45888 8032
rect 45940 7478 45968 9862
rect 46032 9722 46060 9998
rect 46940 9988 46992 9994
rect 46940 9930 46992 9936
rect 46480 9920 46532 9926
rect 46480 9862 46532 9868
rect 46020 9716 46072 9722
rect 46020 9658 46072 9664
rect 46032 8498 46060 9658
rect 46492 9586 46520 9862
rect 46756 9648 46808 9654
rect 46756 9590 46808 9596
rect 46480 9580 46532 9586
rect 46480 9522 46532 9528
rect 46572 9580 46624 9586
rect 46572 9522 46624 9528
rect 46584 8566 46612 9522
rect 46768 9450 46796 9590
rect 46756 9444 46808 9450
rect 46756 9386 46808 9392
rect 46664 9376 46716 9382
rect 46664 9318 46716 9324
rect 46572 8560 46624 8566
rect 46572 8502 46624 8508
rect 46020 8492 46072 8498
rect 46020 8434 46072 8440
rect 46204 8492 46256 8498
rect 46204 8434 46256 8440
rect 46032 8362 46060 8434
rect 46020 8356 46072 8362
rect 46020 8298 46072 8304
rect 46112 8016 46164 8022
rect 46112 7958 46164 7964
rect 46020 7744 46072 7750
rect 46020 7686 46072 7692
rect 46032 7546 46060 7686
rect 46020 7540 46072 7546
rect 46020 7482 46072 7488
rect 45928 7472 45980 7478
rect 45374 7440 45430 7449
rect 45928 7414 45980 7420
rect 45374 7375 45430 7384
rect 45388 6730 45416 7375
rect 45940 7002 45968 7414
rect 46124 7206 46152 7958
rect 46216 7818 46244 8434
rect 46676 7886 46704 9318
rect 46756 8900 46808 8906
rect 46756 8842 46808 8848
rect 46768 8498 46796 8842
rect 46952 8634 46980 9930
rect 47228 9586 47256 11018
rect 47596 10674 47624 11630
rect 47780 11286 47808 11766
rect 47860 11688 47912 11694
rect 47860 11630 47912 11636
rect 47872 11354 47900 11630
rect 47860 11348 47912 11354
rect 47860 11290 47912 11296
rect 47768 11280 47820 11286
rect 47768 11222 47820 11228
rect 48332 11218 48360 13194
rect 48424 12918 48452 13874
rect 48516 13308 48544 15302
rect 48792 15094 48820 16594
rect 48780 15088 48832 15094
rect 48780 15030 48832 15036
rect 48596 14952 48648 14958
rect 48688 14952 48740 14958
rect 48596 14894 48648 14900
rect 48686 14920 48688 14929
rect 48740 14920 48742 14929
rect 48608 14278 48636 14894
rect 48686 14855 48742 14864
rect 48700 14822 48728 14855
rect 48688 14816 48740 14822
rect 48688 14758 48740 14764
rect 48884 14550 48912 17478
rect 49252 16998 49280 17682
rect 50172 17678 50200 18566
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50724 17678 50752 18566
rect 50816 18426 50844 18770
rect 50804 18420 50856 18426
rect 50804 18362 50856 18368
rect 51080 18284 51132 18290
rect 51080 18226 51132 18232
rect 51092 17882 51120 18226
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 51080 17876 51132 17882
rect 51080 17818 51132 17824
rect 50160 17672 50212 17678
rect 50160 17614 50212 17620
rect 50712 17672 50764 17678
rect 50712 17614 50764 17620
rect 50068 17536 50120 17542
rect 50068 17478 50120 17484
rect 50080 17202 50108 17478
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50068 17196 50120 17202
rect 50068 17138 50120 17144
rect 68466 17096 68522 17105
rect 49792 17060 49844 17066
rect 68466 17031 68468 17040
rect 49792 17002 49844 17008
rect 68520 17031 68522 17040
rect 68468 17002 68520 17008
rect 49240 16992 49292 16998
rect 49240 16934 49292 16940
rect 49252 16658 49280 16934
rect 49240 16652 49292 16658
rect 49240 16594 49292 16600
rect 49804 16522 49832 17002
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 51816 16584 51868 16590
rect 51816 16526 51868 16532
rect 49792 16516 49844 16522
rect 49792 16458 49844 16464
rect 49700 16448 49752 16454
rect 49700 16390 49752 16396
rect 48964 15904 49016 15910
rect 48964 15846 49016 15852
rect 48976 15162 49004 15846
rect 48964 15156 49016 15162
rect 48964 15098 49016 15104
rect 49148 14952 49200 14958
rect 49148 14894 49200 14900
rect 49160 14618 49188 14894
rect 49712 14618 49740 16390
rect 49804 15502 49832 16458
rect 51448 16448 51500 16454
rect 51448 16390 51500 16396
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 51460 16182 51488 16390
rect 51828 16250 51856 16526
rect 52368 16448 52420 16454
rect 52368 16390 52420 16396
rect 52736 16448 52788 16454
rect 52736 16390 52788 16396
rect 51816 16244 51868 16250
rect 51816 16186 51868 16192
rect 51448 16176 51500 16182
rect 51448 16118 51500 16124
rect 50436 16040 50488 16046
rect 51828 15994 51856 16186
rect 50436 15982 50488 15988
rect 50448 15706 50476 15982
rect 51736 15966 51856 15994
rect 50436 15700 50488 15706
rect 50436 15642 50488 15648
rect 49792 15496 49844 15502
rect 49792 15438 49844 15444
rect 49804 14822 49832 15438
rect 51632 15428 51684 15434
rect 51632 15370 51684 15376
rect 49884 15360 49936 15366
rect 49884 15302 49936 15308
rect 49896 15094 49924 15302
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 51644 15094 51672 15370
rect 51736 15162 51764 15966
rect 52276 15904 52328 15910
rect 52276 15846 52328 15852
rect 52000 15700 52052 15706
rect 52000 15642 52052 15648
rect 51816 15496 51868 15502
rect 51816 15438 51868 15444
rect 51724 15156 51776 15162
rect 51724 15098 51776 15104
rect 49884 15088 49936 15094
rect 49884 15030 49936 15036
rect 51264 15088 51316 15094
rect 51264 15030 51316 15036
rect 51632 15088 51684 15094
rect 51632 15030 51684 15036
rect 49792 14816 49844 14822
rect 49792 14758 49844 14764
rect 50712 14816 50764 14822
rect 50712 14758 50764 14764
rect 48964 14612 49016 14618
rect 48964 14554 49016 14560
rect 49148 14612 49200 14618
rect 49148 14554 49200 14560
rect 49700 14612 49752 14618
rect 49700 14554 49752 14560
rect 48688 14544 48740 14550
rect 48688 14486 48740 14492
rect 48872 14544 48924 14550
rect 48872 14486 48924 14492
rect 48700 14346 48728 14486
rect 48872 14408 48924 14414
rect 48872 14350 48924 14356
rect 48688 14340 48740 14346
rect 48688 14282 48740 14288
rect 48596 14272 48648 14278
rect 48596 14214 48648 14220
rect 48700 13938 48728 14282
rect 48884 13938 48912 14350
rect 48688 13932 48740 13938
rect 48688 13874 48740 13880
rect 48872 13932 48924 13938
rect 48872 13874 48924 13880
rect 48780 13728 48832 13734
rect 48780 13670 48832 13676
rect 48792 13530 48820 13670
rect 48780 13524 48832 13530
rect 48780 13466 48832 13472
rect 48596 13320 48648 13326
rect 48516 13280 48596 13308
rect 48596 13262 48648 13268
rect 48792 13190 48820 13466
rect 48976 13410 49004 14554
rect 49620 14470 49832 14498
rect 49620 14074 49648 14470
rect 49804 14414 49832 14470
rect 49700 14408 49752 14414
rect 49700 14350 49752 14356
rect 49792 14408 49844 14414
rect 49792 14350 49844 14356
rect 49712 14074 49740 14350
rect 50160 14340 50212 14346
rect 50160 14282 50212 14288
rect 50620 14340 50672 14346
rect 50620 14282 50672 14288
rect 49608 14068 49660 14074
rect 49608 14010 49660 14016
rect 49700 14068 49752 14074
rect 49700 14010 49752 14016
rect 49148 13932 49200 13938
rect 49148 13874 49200 13880
rect 49240 13932 49292 13938
rect 49240 13874 49292 13880
rect 49160 13462 49188 13874
rect 48884 13382 49004 13410
rect 49148 13456 49200 13462
rect 49148 13398 49200 13404
rect 48884 13326 48912 13382
rect 48872 13320 48924 13326
rect 48872 13262 48924 13268
rect 48780 13184 48832 13190
rect 48780 13126 48832 13132
rect 48964 13184 49016 13190
rect 48964 13126 49016 13132
rect 48412 12912 48464 12918
rect 48412 12854 48464 12860
rect 48976 12782 49004 13126
rect 49160 12850 49188 13398
rect 49252 13326 49280 13874
rect 49424 13864 49476 13870
rect 49424 13806 49476 13812
rect 49240 13320 49292 13326
rect 49240 13262 49292 13268
rect 49332 13320 49384 13326
rect 49332 13262 49384 13268
rect 49148 12844 49200 12850
rect 49148 12786 49200 12792
rect 48964 12776 49016 12782
rect 48964 12718 49016 12724
rect 49160 12434 49188 12786
rect 49344 12782 49372 13262
rect 49332 12776 49384 12782
rect 49332 12718 49384 12724
rect 49436 12434 49464 13806
rect 49620 12646 49648 14010
rect 49792 14000 49844 14006
rect 49792 13942 49844 13948
rect 49804 13530 49832 13942
rect 50172 13802 50200 14282
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50252 13932 50304 13938
rect 50252 13874 50304 13880
rect 50160 13796 50212 13802
rect 50160 13738 50212 13744
rect 49792 13524 49844 13530
rect 49792 13466 49844 13472
rect 50264 13326 50292 13874
rect 50632 13394 50660 14282
rect 50724 13870 50752 14758
rect 51276 14618 51304 15030
rect 51448 14952 51500 14958
rect 51448 14894 51500 14900
rect 51264 14612 51316 14618
rect 51264 14554 51316 14560
rect 50988 14408 51040 14414
rect 50988 14350 51040 14356
rect 51276 14362 51304 14554
rect 51460 14414 51488 14894
rect 51540 14816 51592 14822
rect 51828 14804 51856 15438
rect 52012 15366 52040 15642
rect 52092 15428 52144 15434
rect 52092 15370 52144 15376
rect 52184 15428 52236 15434
rect 52184 15370 52236 15376
rect 52000 15360 52052 15366
rect 52000 15302 52052 15308
rect 52104 15026 52132 15370
rect 52092 15020 52144 15026
rect 52092 14962 52144 14968
rect 52196 14929 52224 15370
rect 52288 15094 52316 15846
rect 52380 15706 52408 16390
rect 52368 15700 52420 15706
rect 52368 15642 52420 15648
rect 52552 15632 52604 15638
rect 52552 15574 52604 15580
rect 52460 15360 52512 15366
rect 52460 15302 52512 15308
rect 52276 15088 52328 15094
rect 52276 15030 52328 15036
rect 52472 15026 52500 15302
rect 52564 15026 52592 15574
rect 52644 15496 52696 15502
rect 52644 15438 52696 15444
rect 52460 15020 52512 15026
rect 52460 14962 52512 14968
rect 52552 15020 52604 15026
rect 52552 14962 52604 14968
rect 52182 14920 52238 14929
rect 52182 14855 52238 14864
rect 51592 14776 51856 14804
rect 52000 14816 52052 14822
rect 51540 14758 51592 14764
rect 52000 14758 52052 14764
rect 52012 14618 52040 14758
rect 52000 14612 52052 14618
rect 52000 14554 52052 14560
rect 51448 14408 51500 14414
rect 50804 14340 50856 14346
rect 50804 14282 50856 14288
rect 50816 14074 50844 14282
rect 50804 14068 50856 14074
rect 50804 14010 50856 14016
rect 50712 13864 50764 13870
rect 50712 13806 50764 13812
rect 51000 13462 51028 14350
rect 51276 14334 51396 14362
rect 51448 14350 51500 14356
rect 51264 14272 51316 14278
rect 51264 14214 51316 14220
rect 51276 14006 51304 14214
rect 51264 14000 51316 14006
rect 51264 13942 51316 13948
rect 51172 13864 51224 13870
rect 51172 13806 51224 13812
rect 50988 13456 51040 13462
rect 50988 13398 51040 13404
rect 50620 13388 50672 13394
rect 50620 13330 50672 13336
rect 50896 13388 50948 13394
rect 50896 13330 50948 13336
rect 50252 13320 50304 13326
rect 50252 13262 50304 13268
rect 49700 13252 49752 13258
rect 49700 13194 49752 13200
rect 49712 12782 49740 13194
rect 49976 13184 50028 13190
rect 49976 13126 50028 13132
rect 50068 13184 50120 13190
rect 50068 13126 50120 13132
rect 49988 12782 50016 13126
rect 50080 12850 50108 13126
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50908 12850 50936 13330
rect 50068 12844 50120 12850
rect 50068 12786 50120 12792
rect 50528 12844 50580 12850
rect 50528 12786 50580 12792
rect 50896 12844 50948 12850
rect 50896 12786 50948 12792
rect 49700 12776 49752 12782
rect 49700 12718 49752 12724
rect 49976 12776 50028 12782
rect 49976 12718 50028 12724
rect 49608 12640 49660 12646
rect 49608 12582 49660 12588
rect 49160 12406 49372 12434
rect 49436 12406 49648 12434
rect 49344 12170 49372 12406
rect 49332 12164 49384 12170
rect 49332 12106 49384 12112
rect 49344 11898 49372 12106
rect 49332 11892 49384 11898
rect 49332 11834 49384 11840
rect 48320 11212 48372 11218
rect 48320 11154 48372 11160
rect 49344 11150 49372 11834
rect 49620 11778 49648 12406
rect 49988 12238 50016 12718
rect 50540 12306 50568 12786
rect 50528 12300 50580 12306
rect 50528 12242 50580 12248
rect 49976 12232 50028 12238
rect 49976 12174 50028 12180
rect 49884 11824 49936 11830
rect 49620 11772 49884 11778
rect 49620 11766 49936 11772
rect 49620 11750 49924 11766
rect 49620 11626 49648 11750
rect 49608 11620 49660 11626
rect 49608 11562 49660 11568
rect 49516 11552 49568 11558
rect 49516 11494 49568 11500
rect 49332 11144 49384 11150
rect 49332 11086 49384 11092
rect 49240 11008 49292 11014
rect 49240 10950 49292 10956
rect 49252 10674 49280 10950
rect 49528 10742 49556 11494
rect 49620 11082 49648 11562
rect 49988 11218 50016 12174
rect 51000 12170 51028 13398
rect 51184 13326 51212 13806
rect 51368 13734 51396 14334
rect 51356 13728 51408 13734
rect 51356 13670 51408 13676
rect 51460 13530 51488 14350
rect 51632 14272 51684 14278
rect 51632 14214 51684 14220
rect 51448 13524 51500 13530
rect 51448 13466 51500 13472
rect 51644 13462 51672 14214
rect 51816 13864 51868 13870
rect 51816 13806 51868 13812
rect 51724 13796 51776 13802
rect 51724 13738 51776 13744
rect 51736 13530 51764 13738
rect 51724 13524 51776 13530
rect 51724 13466 51776 13472
rect 51632 13456 51684 13462
rect 51632 13398 51684 13404
rect 51172 13320 51224 13326
rect 51172 13262 51224 13268
rect 51356 13320 51408 13326
rect 51356 13262 51408 13268
rect 51540 13320 51592 13326
rect 51540 13262 51592 13268
rect 51368 12986 51396 13262
rect 51448 13252 51500 13258
rect 51448 13194 51500 13200
rect 51356 12980 51408 12986
rect 51356 12922 51408 12928
rect 51264 12776 51316 12782
rect 51264 12718 51316 12724
rect 51276 12442 51304 12718
rect 51460 12442 51488 13194
rect 51552 12782 51580 13262
rect 51644 12918 51672 13398
rect 51632 12912 51684 12918
rect 51632 12854 51684 12860
rect 51540 12776 51592 12782
rect 51828 12730 51856 13806
rect 52000 13320 52052 13326
rect 52000 13262 52052 13268
rect 51540 12718 51592 12724
rect 51736 12702 51856 12730
rect 51264 12436 51316 12442
rect 51264 12378 51316 12384
rect 51448 12436 51500 12442
rect 51736 12434 51764 12702
rect 51816 12640 51868 12646
rect 51868 12588 51948 12594
rect 51816 12582 51948 12588
rect 51828 12566 51948 12582
rect 51736 12406 51856 12434
rect 51448 12378 51500 12384
rect 50988 12164 51040 12170
rect 50988 12106 51040 12112
rect 50160 12096 50212 12102
rect 50160 12038 50212 12044
rect 50620 12096 50672 12102
rect 50620 12038 50672 12044
rect 50172 11898 50200 12038
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50160 11892 50212 11898
rect 50160 11834 50212 11840
rect 50344 11824 50396 11830
rect 50342 11792 50344 11801
rect 50528 11824 50580 11830
rect 50396 11792 50398 11801
rect 50528 11766 50580 11772
rect 50342 11727 50398 11736
rect 50436 11688 50488 11694
rect 50540 11676 50568 11766
rect 50488 11648 50568 11676
rect 50436 11630 50488 11636
rect 50632 11354 50660 12038
rect 51000 11830 51028 12106
rect 51276 11914 51304 12378
rect 51460 12306 51488 12378
rect 51448 12300 51500 12306
rect 51448 12242 51500 12248
rect 51448 12096 51500 12102
rect 51448 12038 51500 12044
rect 51276 11886 51396 11914
rect 51460 11898 51488 12038
rect 50988 11824 51040 11830
rect 50988 11766 51040 11772
rect 50620 11348 50672 11354
rect 50620 11290 50672 11296
rect 49976 11212 50028 11218
rect 49976 11154 50028 11160
rect 49608 11076 49660 11082
rect 49608 11018 49660 11024
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 51000 10810 51028 11766
rect 51264 11552 51316 11558
rect 51264 11494 51316 11500
rect 51276 11354 51304 11494
rect 51368 11354 51396 11886
rect 51448 11892 51500 11898
rect 51448 11834 51500 11840
rect 51540 11756 51592 11762
rect 51540 11698 51592 11704
rect 51552 11642 51580 11698
rect 51552 11626 51764 11642
rect 51552 11620 51776 11626
rect 51552 11614 51724 11620
rect 51724 11562 51776 11568
rect 51828 11558 51856 12406
rect 51920 11762 51948 12566
rect 51908 11756 51960 11762
rect 51908 11698 51960 11704
rect 51816 11552 51868 11558
rect 51816 11494 51868 11500
rect 51264 11348 51316 11354
rect 51264 11290 51316 11296
rect 51356 11348 51408 11354
rect 51356 11290 51408 11296
rect 52012 11218 52040 13262
rect 52196 12850 52224 14855
rect 52472 14414 52500 14962
rect 52564 14414 52592 14962
rect 52656 14618 52684 15438
rect 52644 14612 52696 14618
rect 52644 14554 52696 14560
rect 52748 14414 52776 16390
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 54484 15496 54536 15502
rect 54484 15438 54536 15444
rect 53932 15360 53984 15366
rect 53932 15302 53984 15308
rect 53944 15162 53972 15302
rect 54496 15162 54524 15438
rect 53932 15156 53984 15162
rect 53932 15098 53984 15104
rect 54484 15156 54536 15162
rect 54484 15098 54536 15104
rect 53472 15088 53524 15094
rect 53472 15030 53524 15036
rect 53484 14618 53512 15030
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 53472 14612 53524 14618
rect 53472 14554 53524 14560
rect 52460 14408 52512 14414
rect 52460 14350 52512 14356
rect 52552 14408 52604 14414
rect 52552 14350 52604 14356
rect 52736 14408 52788 14414
rect 68468 14408 68520 14414
rect 52736 14350 52788 14356
rect 68466 14376 68468 14385
rect 68520 14376 68522 14385
rect 52564 13938 52592 14350
rect 53472 14340 53524 14346
rect 68466 14311 68522 14320
rect 53472 14282 53524 14288
rect 52552 13932 52604 13938
rect 52552 13874 52604 13880
rect 53484 12850 53512 14282
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 53564 13252 53616 13258
rect 53564 13194 53616 13200
rect 53576 12986 53604 13194
rect 53748 13184 53800 13190
rect 53748 13126 53800 13132
rect 53760 12986 53788 13126
rect 53564 12980 53616 12986
rect 53564 12922 53616 12928
rect 53748 12980 53800 12986
rect 53748 12922 53800 12928
rect 52184 12844 52236 12850
rect 52184 12786 52236 12792
rect 53472 12844 53524 12850
rect 53472 12786 53524 12792
rect 52092 12164 52144 12170
rect 52092 12106 52144 12112
rect 52104 11830 52132 12106
rect 52196 11898 52224 12786
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 52184 11892 52236 11898
rect 52184 11834 52236 11840
rect 52092 11824 52144 11830
rect 52196 11801 52224 11834
rect 52092 11766 52144 11772
rect 52182 11792 52238 11801
rect 52182 11727 52238 11736
rect 52276 11756 52328 11762
rect 52276 11698 52328 11704
rect 52288 11218 52316 11698
rect 68466 11656 68522 11665
rect 68466 11591 68468 11600
rect 68520 11591 68522 11600
rect 68468 11562 68520 11568
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 52000 11212 52052 11218
rect 52000 11154 52052 11160
rect 52276 11212 52328 11218
rect 52276 11154 52328 11160
rect 51448 11076 51500 11082
rect 51448 11018 51500 11024
rect 51460 10810 51488 11018
rect 50988 10804 51040 10810
rect 50988 10746 51040 10752
rect 51448 10804 51500 10810
rect 51448 10746 51500 10752
rect 49516 10736 49568 10742
rect 49516 10678 49568 10684
rect 47584 10668 47636 10674
rect 47584 10610 47636 10616
rect 49240 10668 49292 10674
rect 49240 10610 49292 10616
rect 51080 10668 51132 10674
rect 51080 10610 51132 10616
rect 47596 10130 47624 10610
rect 47584 10124 47636 10130
rect 47584 10066 47636 10072
rect 48044 9988 48096 9994
rect 48044 9930 48096 9936
rect 47216 9580 47268 9586
rect 47216 9522 47268 9528
rect 47860 9580 47912 9586
rect 47860 9522 47912 9528
rect 47952 9580 48004 9586
rect 47952 9522 48004 9528
rect 47308 9376 47360 9382
rect 47308 9318 47360 9324
rect 47676 9376 47728 9382
rect 47676 9318 47728 9324
rect 47032 9036 47084 9042
rect 47032 8978 47084 8984
rect 46940 8628 46992 8634
rect 46940 8570 46992 8576
rect 46756 8492 46808 8498
rect 46756 8434 46808 8440
rect 46388 7880 46440 7886
rect 46388 7822 46440 7828
rect 46664 7880 46716 7886
rect 46664 7822 46716 7828
rect 46204 7812 46256 7818
rect 46204 7754 46256 7760
rect 46112 7200 46164 7206
rect 46164 7160 46244 7188
rect 46112 7142 46164 7148
rect 45928 6996 45980 7002
rect 45928 6938 45980 6944
rect 45940 6798 45968 6938
rect 45928 6792 45980 6798
rect 45928 6734 45980 6740
rect 46112 6792 46164 6798
rect 46112 6734 46164 6740
rect 44272 6724 44324 6730
rect 44272 6666 44324 6672
rect 45376 6724 45428 6730
rect 45376 6666 45428 6672
rect 46020 6724 46072 6730
rect 46020 6666 46072 6672
rect 44284 6458 44312 6666
rect 44272 6452 44324 6458
rect 44272 6394 44324 6400
rect 43904 6384 43956 6390
rect 43904 6326 43956 6332
rect 43916 5710 43944 6326
rect 43904 5704 43956 5710
rect 43904 5646 43956 5652
rect 41972 5636 42024 5642
rect 41972 5578 42024 5584
rect 41984 5370 42012 5578
rect 41972 5364 42024 5370
rect 41972 5306 42024 5312
rect 41512 5228 41564 5234
rect 41512 5170 41564 5176
rect 42432 5160 42484 5166
rect 42432 5102 42484 5108
rect 43720 5160 43772 5166
rect 43720 5102 43772 5108
rect 42444 4826 42472 5102
rect 43732 4826 43760 5102
rect 42432 4820 42484 4826
rect 42432 4762 42484 4768
rect 43720 4820 43772 4826
rect 43720 4762 43772 4768
rect 43916 4622 43944 5646
rect 45388 5370 45416 6666
rect 45836 6248 45888 6254
rect 45836 6190 45888 6196
rect 45848 5778 45876 6190
rect 46032 6186 46060 6666
rect 46124 6390 46152 6734
rect 46216 6730 46244 7160
rect 46204 6724 46256 6730
rect 46204 6666 46256 6672
rect 46216 6390 46244 6666
rect 46112 6384 46164 6390
rect 46112 6326 46164 6332
rect 46204 6384 46256 6390
rect 46256 6344 46336 6372
rect 46204 6326 46256 6332
rect 46020 6180 46072 6186
rect 46020 6122 46072 6128
rect 45836 5772 45888 5778
rect 45836 5714 45888 5720
rect 45376 5364 45428 5370
rect 45376 5306 45428 5312
rect 46032 5302 46060 6122
rect 46124 5846 46152 6326
rect 46204 6112 46256 6118
rect 46204 6054 46256 6060
rect 46216 5914 46244 6054
rect 46204 5908 46256 5914
rect 46204 5850 46256 5856
rect 46112 5840 46164 5846
rect 46112 5782 46164 5788
rect 44456 5296 44508 5302
rect 44456 5238 44508 5244
rect 46020 5296 46072 5302
rect 46020 5238 46072 5244
rect 44468 4826 44496 5238
rect 46124 5166 46152 5782
rect 46308 5778 46336 6344
rect 46400 5914 46428 7822
rect 46676 7392 46704 7822
rect 46768 7410 46796 8434
rect 47044 8430 47072 8978
rect 47320 8906 47348 9318
rect 47688 9178 47716 9318
rect 47872 9178 47900 9522
rect 47676 9172 47728 9178
rect 47676 9114 47728 9120
rect 47860 9172 47912 9178
rect 47860 9114 47912 9120
rect 47308 8900 47360 8906
rect 47308 8842 47360 8848
rect 47964 8634 47992 9522
rect 48056 9518 48084 9930
rect 48964 9648 49016 9654
rect 48964 9590 49016 9596
rect 48044 9512 48096 9518
rect 48044 9454 48096 9460
rect 48056 9178 48084 9454
rect 48044 9172 48096 9178
rect 48044 9114 48096 9120
rect 48228 9172 48280 9178
rect 48228 9114 48280 9120
rect 47952 8628 48004 8634
rect 47952 8570 48004 8576
rect 47032 8424 47084 8430
rect 47032 8366 47084 8372
rect 46584 7364 46704 7392
rect 46756 7404 46808 7410
rect 46480 7200 46532 7206
rect 46480 7142 46532 7148
rect 46492 6934 46520 7142
rect 46480 6928 46532 6934
rect 46480 6870 46532 6876
rect 46584 6322 46612 7364
rect 46756 7346 46808 7352
rect 46664 7200 46716 7206
rect 46664 7142 46716 7148
rect 46848 7200 46900 7206
rect 46848 7142 46900 7148
rect 46676 6390 46704 7142
rect 46756 6792 46808 6798
rect 46756 6734 46808 6740
rect 46664 6384 46716 6390
rect 46664 6326 46716 6332
rect 46572 6316 46624 6322
rect 46572 6258 46624 6264
rect 46768 6254 46796 6734
rect 46756 6248 46808 6254
rect 46756 6190 46808 6196
rect 46572 6180 46624 6186
rect 46572 6122 46624 6128
rect 46388 5908 46440 5914
rect 46388 5850 46440 5856
rect 46296 5772 46348 5778
rect 46296 5714 46348 5720
rect 46480 5364 46532 5370
rect 46480 5306 46532 5312
rect 46492 5234 46520 5306
rect 46584 5234 46612 6122
rect 46768 5914 46796 6190
rect 46756 5908 46808 5914
rect 46756 5850 46808 5856
rect 46860 5574 46888 7142
rect 47044 6798 47072 8366
rect 47964 8090 47992 8570
rect 48056 8566 48084 9114
rect 48240 8838 48268 9114
rect 48976 8974 49004 9590
rect 49252 9586 49280 10610
rect 50160 10056 50212 10062
rect 50160 9998 50212 10004
rect 50068 9920 50120 9926
rect 50068 9862 50120 9868
rect 49240 9580 49292 9586
rect 49240 9522 49292 9528
rect 49148 9376 49200 9382
rect 49148 9318 49200 9324
rect 49160 9178 49188 9318
rect 49056 9172 49108 9178
rect 49056 9114 49108 9120
rect 49148 9172 49200 9178
rect 49148 9114 49200 9120
rect 48596 8968 48648 8974
rect 48596 8910 48648 8916
rect 48780 8968 48832 8974
rect 48780 8910 48832 8916
rect 48872 8968 48924 8974
rect 48872 8910 48924 8916
rect 48964 8968 49016 8974
rect 48964 8910 49016 8916
rect 48228 8832 48280 8838
rect 48228 8774 48280 8780
rect 48044 8560 48096 8566
rect 48044 8502 48096 8508
rect 47952 8084 48004 8090
rect 47952 8026 48004 8032
rect 47768 7948 47820 7954
rect 47768 7890 47820 7896
rect 47676 7880 47728 7886
rect 47676 7822 47728 7828
rect 47688 7546 47716 7822
rect 47780 7750 47808 7890
rect 48240 7834 48268 8774
rect 48608 8634 48636 8910
rect 48792 8634 48820 8910
rect 48884 8820 48912 8910
rect 49068 8906 49096 9114
rect 50080 8974 50108 9862
rect 50172 9722 50200 9998
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50160 9716 50212 9722
rect 50160 9658 50212 9664
rect 51092 9586 51120 10610
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 51080 9580 51132 9586
rect 51080 9522 51132 9528
rect 51448 9512 51500 9518
rect 51448 9454 51500 9460
rect 49792 8968 49844 8974
rect 49712 8916 49792 8922
rect 49712 8910 49844 8916
rect 50068 8968 50120 8974
rect 50068 8910 50120 8916
rect 49056 8900 49108 8906
rect 49056 8842 49108 8848
rect 49712 8894 49832 8910
rect 48964 8832 49016 8838
rect 48884 8792 48964 8820
rect 48596 8628 48648 8634
rect 48596 8570 48648 8576
rect 48780 8628 48832 8634
rect 48780 8570 48832 8576
rect 48884 8498 48912 8792
rect 48964 8774 49016 8780
rect 49332 8628 49384 8634
rect 49332 8570 49384 8576
rect 48872 8492 48924 8498
rect 48872 8434 48924 8440
rect 49344 8294 49372 8570
rect 49712 8566 49740 8894
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 49700 8560 49752 8566
rect 49700 8502 49752 8508
rect 49332 8288 49384 8294
rect 49332 8230 49384 8236
rect 49344 7954 49372 8230
rect 49332 7948 49384 7954
rect 49332 7890 49384 7896
rect 48056 7806 48268 7834
rect 48412 7812 48464 7818
rect 47768 7744 47820 7750
rect 47768 7686 47820 7692
rect 47676 7540 47728 7546
rect 47676 7482 47728 7488
rect 47780 7342 47808 7686
rect 48056 7410 48084 7806
rect 48412 7754 48464 7760
rect 49516 7812 49568 7818
rect 49516 7754 49568 7760
rect 48136 7744 48188 7750
rect 48136 7686 48188 7692
rect 48320 7744 48372 7750
rect 48320 7686 48372 7692
rect 48148 7478 48176 7686
rect 48332 7546 48360 7686
rect 48424 7546 48452 7754
rect 48596 7744 48648 7750
rect 48596 7686 48648 7692
rect 49148 7744 49200 7750
rect 49148 7686 49200 7692
rect 48608 7546 48636 7686
rect 49160 7546 49188 7686
rect 48320 7540 48372 7546
rect 48320 7482 48372 7488
rect 48412 7540 48464 7546
rect 48412 7482 48464 7488
rect 48596 7540 48648 7546
rect 48596 7482 48648 7488
rect 49148 7540 49200 7546
rect 49148 7482 49200 7488
rect 49528 7478 49556 7754
rect 48136 7472 48188 7478
rect 48134 7440 48136 7449
rect 49516 7472 49568 7478
rect 48188 7440 48190 7449
rect 48044 7404 48096 7410
rect 49516 7414 49568 7420
rect 49712 7410 49740 8502
rect 51460 8498 51488 9454
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 68468 8968 68520 8974
rect 68466 8936 68468 8945
rect 68520 8936 68522 8945
rect 68466 8871 68522 8880
rect 51448 8492 51500 8498
rect 51448 8434 51500 8440
rect 49792 8424 49844 8430
rect 49792 8366 49844 8372
rect 49804 8090 49832 8366
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 49792 8084 49844 8090
rect 49792 8026 49844 8032
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 48134 7375 48190 7384
rect 49700 7404 49752 7410
rect 48044 7346 48096 7352
rect 49700 7346 49752 7352
rect 47768 7336 47820 7342
rect 47768 7278 47820 7284
rect 47032 6792 47084 6798
rect 47032 6734 47084 6740
rect 46940 5772 46992 5778
rect 46940 5714 46992 5720
rect 46848 5568 46900 5574
rect 46848 5510 46900 5516
rect 46860 5370 46888 5510
rect 46848 5364 46900 5370
rect 46848 5306 46900 5312
rect 46860 5234 46888 5306
rect 46952 5234 46980 5714
rect 47044 5710 47072 6734
rect 48056 6338 48084 7346
rect 49792 7268 49844 7274
rect 49792 7210 49844 7216
rect 49056 7200 49108 7206
rect 49056 7142 49108 7148
rect 49068 7002 49096 7142
rect 49804 7002 49832 7210
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 49056 6996 49108 7002
rect 49056 6938 49108 6944
rect 49792 6996 49844 7002
rect 49792 6938 49844 6944
rect 48780 6724 48832 6730
rect 48780 6666 48832 6672
rect 48792 6458 48820 6666
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 48780 6452 48832 6458
rect 48780 6394 48832 6400
rect 47964 6322 48084 6338
rect 47952 6316 48084 6322
rect 48004 6310 48084 6316
rect 48320 6316 48372 6322
rect 47952 6258 48004 6264
rect 48320 6258 48372 6264
rect 47400 6112 47452 6118
rect 47400 6054 47452 6060
rect 47412 5778 47440 6054
rect 47400 5772 47452 5778
rect 47400 5714 47452 5720
rect 47032 5704 47084 5710
rect 47032 5646 47084 5652
rect 48332 5658 48360 6258
rect 68466 6216 68522 6225
rect 68466 6151 68468 6160
rect 68520 6151 68522 6160
rect 68468 6122 68520 6128
rect 48872 6112 48924 6118
rect 48872 6054 48924 6060
rect 48884 5914 48912 6054
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 48872 5908 48924 5914
rect 48872 5850 48924 5856
rect 48412 5704 48464 5710
rect 48332 5652 48412 5658
rect 48332 5646 48464 5652
rect 46480 5228 46532 5234
rect 46480 5170 46532 5176
rect 46572 5228 46624 5234
rect 46572 5170 46624 5176
rect 46848 5228 46900 5234
rect 46848 5170 46900 5176
rect 46940 5228 46992 5234
rect 46940 5170 46992 5176
rect 46112 5160 46164 5166
rect 46112 5102 46164 5108
rect 45100 5024 45152 5030
rect 45100 4966 45152 4972
rect 45284 5024 45336 5030
rect 45284 4966 45336 4972
rect 45928 5024 45980 5030
rect 45928 4966 45980 4972
rect 44456 4820 44508 4826
rect 44456 4762 44508 4768
rect 45112 4690 45140 4966
rect 45296 4826 45324 4966
rect 45940 4826 45968 4966
rect 45284 4820 45336 4826
rect 45284 4762 45336 4768
rect 45928 4820 45980 4826
rect 45928 4762 45980 4768
rect 47044 4690 47072 5646
rect 48332 5630 48452 5646
rect 47584 5228 47636 5234
rect 47584 5170 47636 5176
rect 45100 4684 45152 4690
rect 45100 4626 45152 4632
rect 47032 4684 47084 4690
rect 47032 4626 47084 4632
rect 47596 4622 47624 5170
rect 48332 4622 48360 5630
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 43904 4616 43956 4622
rect 43904 4558 43956 4564
rect 47584 4616 47636 4622
rect 47584 4558 47636 4564
rect 48320 4616 48372 4622
rect 48320 4558 48372 4564
rect 41328 4548 41380 4554
rect 41328 4490 41380 4496
rect 40500 4208 40552 4214
rect 40500 4150 40552 4156
rect 40592 4072 40644 4078
rect 40592 4014 40644 4020
rect 40408 3460 40460 3466
rect 40408 3402 40460 3408
rect 40604 2582 40632 4014
rect 41340 3602 41368 4490
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41432 3670 41460 3878
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 41420 3664 41472 3670
rect 41420 3606 41472 3612
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 68468 3528 68520 3534
rect 68466 3496 68468 3505
rect 68520 3496 68522 3505
rect 68466 3431 68522 3440
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 40684 3120 40736 3126
rect 40684 3062 40736 3068
rect 40696 2650 40724 3062
rect 48320 2848 48372 2854
rect 48320 2790 48372 2796
rect 40684 2644 40736 2650
rect 40684 2586 40736 2592
rect 40592 2576 40644 2582
rect 40592 2518 40644 2524
rect 48332 2446 48360 2790
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 40132 2440 40184 2446
rect 40132 2382 40184 2388
rect 43168 2440 43220 2446
rect 43168 2382 43220 2388
rect 45744 2440 45796 2446
rect 45744 2382 45796 2388
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 50896 2440 50948 2446
rect 50896 2382 50948 2388
rect 53472 2440 53524 2446
rect 53472 2382 53524 2388
rect 56048 2440 56100 2446
rect 56048 2382 56100 2388
rect 58624 2440 58676 2446
rect 58624 2382 58676 2388
rect 66352 2440 66404 2446
rect 66352 2382 66404 2388
rect 68468 2440 68520 2446
rect 68468 2382 68520 2388
rect 68652 2440 68704 2446
rect 68652 2382 68704 2388
rect 39212 2372 39264 2378
rect 39212 2314 39264 2320
rect 43180 800 43208 2382
rect 45756 800 45784 2382
rect 48320 2304 48372 2310
rect 48320 2246 48372 2252
rect 48332 800 48360 2246
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50908 800 50936 2382
rect 53484 800 53512 2382
rect 56060 800 56088 2382
rect 58636 800 58664 2382
rect 66364 800 66392 2382
rect 68480 1306 68508 2382
rect 68296 1278 68508 1306
rect 68296 800 68324 1278
rect 38120 734 38332 762
rect 40590 0 40646 800
rect 43166 0 43222 800
rect 45742 0 45798 800
rect 48318 0 48374 800
rect 50894 0 50950 800
rect 53470 0 53526 800
rect 56046 0 56102 800
rect 58622 0 58678 800
rect 61198 0 61254 800
rect 63774 0 63830 800
rect 66350 0 66406 800
rect 68282 0 68338 800
rect 68664 785 68692 2382
rect 68650 776 68706 785
rect 68650 711 68706 720
<< via2 >>
rect 938 67360 994 67416
rect 19580 67482 19636 67484
rect 19660 67482 19716 67484
rect 19740 67482 19796 67484
rect 19820 67482 19876 67484
rect 19580 67430 19626 67482
rect 19626 67430 19636 67482
rect 19660 67430 19690 67482
rect 19690 67430 19702 67482
rect 19702 67430 19716 67482
rect 19740 67430 19754 67482
rect 19754 67430 19766 67482
rect 19766 67430 19796 67482
rect 19820 67430 19830 67482
rect 19830 67430 19876 67482
rect 19580 67428 19636 67430
rect 19660 67428 19716 67430
rect 19740 67428 19796 67430
rect 19820 67428 19876 67430
rect 50300 67482 50356 67484
rect 50380 67482 50436 67484
rect 50460 67482 50516 67484
rect 50540 67482 50596 67484
rect 50300 67430 50346 67482
rect 50346 67430 50356 67482
rect 50380 67430 50410 67482
rect 50410 67430 50422 67482
rect 50422 67430 50436 67482
rect 50460 67430 50474 67482
rect 50474 67430 50486 67482
rect 50486 67430 50516 67482
rect 50540 67430 50550 67482
rect 50550 67430 50596 67482
rect 50300 67428 50356 67430
rect 50380 67428 50436 67430
rect 50460 67428 50516 67430
rect 50540 67428 50596 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 19580 66394 19636 66396
rect 19660 66394 19716 66396
rect 19740 66394 19796 66396
rect 19820 66394 19876 66396
rect 19580 66342 19626 66394
rect 19626 66342 19636 66394
rect 19660 66342 19690 66394
rect 19690 66342 19702 66394
rect 19702 66342 19716 66394
rect 19740 66342 19754 66394
rect 19754 66342 19766 66394
rect 19766 66342 19796 66394
rect 19820 66342 19830 66394
rect 19830 66342 19876 66394
rect 19580 66340 19636 66342
rect 19660 66340 19716 66342
rect 19740 66340 19796 66342
rect 19820 66340 19876 66342
rect 50300 66394 50356 66396
rect 50380 66394 50436 66396
rect 50460 66394 50516 66396
rect 50540 66394 50596 66396
rect 50300 66342 50346 66394
rect 50346 66342 50356 66394
rect 50380 66342 50410 66394
rect 50410 66342 50422 66394
rect 50422 66342 50436 66394
rect 50460 66342 50474 66394
rect 50474 66342 50486 66394
rect 50486 66342 50516 66394
rect 50540 66342 50550 66394
rect 50550 66342 50596 66394
rect 50300 66340 50356 66342
rect 50380 66340 50436 66342
rect 50460 66340 50516 66342
rect 50540 66340 50596 66342
rect 68466 66020 68522 66056
rect 68466 66000 68468 66020
rect 68468 66000 68520 66020
rect 68520 66000 68522 66020
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 19580 65306 19636 65308
rect 19660 65306 19716 65308
rect 19740 65306 19796 65308
rect 19820 65306 19876 65308
rect 19580 65254 19626 65306
rect 19626 65254 19636 65306
rect 19660 65254 19690 65306
rect 19690 65254 19702 65306
rect 19702 65254 19716 65306
rect 19740 65254 19754 65306
rect 19754 65254 19766 65306
rect 19766 65254 19796 65306
rect 19820 65254 19830 65306
rect 19830 65254 19876 65306
rect 19580 65252 19636 65254
rect 19660 65252 19716 65254
rect 19740 65252 19796 65254
rect 19820 65252 19876 65254
rect 50300 65306 50356 65308
rect 50380 65306 50436 65308
rect 50460 65306 50516 65308
rect 50540 65306 50596 65308
rect 50300 65254 50346 65306
rect 50346 65254 50356 65306
rect 50380 65254 50410 65306
rect 50410 65254 50422 65306
rect 50422 65254 50436 65306
rect 50460 65254 50474 65306
rect 50474 65254 50486 65306
rect 50486 65254 50516 65306
rect 50540 65254 50550 65306
rect 50550 65254 50596 65306
rect 50300 65252 50356 65254
rect 50380 65252 50436 65254
rect 50460 65252 50516 65254
rect 50540 65252 50596 65254
rect 1582 64776 1638 64832
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 34940 64762 34996 64764
rect 35020 64762 35076 64764
rect 35100 64762 35156 64764
rect 35180 64762 35236 64764
rect 34940 64710 34986 64762
rect 34986 64710 34996 64762
rect 35020 64710 35050 64762
rect 35050 64710 35062 64762
rect 35062 64710 35076 64762
rect 35100 64710 35114 64762
rect 35114 64710 35126 64762
rect 35126 64710 35156 64762
rect 35180 64710 35190 64762
rect 35190 64710 35236 64762
rect 34940 64708 34996 64710
rect 35020 64708 35076 64710
rect 35100 64708 35156 64710
rect 35180 64708 35236 64710
rect 65660 64762 65716 64764
rect 65740 64762 65796 64764
rect 65820 64762 65876 64764
rect 65900 64762 65956 64764
rect 65660 64710 65706 64762
rect 65706 64710 65716 64762
rect 65740 64710 65770 64762
rect 65770 64710 65782 64762
rect 65782 64710 65796 64762
rect 65820 64710 65834 64762
rect 65834 64710 65846 64762
rect 65846 64710 65876 64762
rect 65900 64710 65910 64762
rect 65910 64710 65956 64762
rect 65660 64708 65716 64710
rect 65740 64708 65796 64710
rect 65820 64708 65876 64710
rect 65900 64708 65956 64710
rect 19580 64218 19636 64220
rect 19660 64218 19716 64220
rect 19740 64218 19796 64220
rect 19820 64218 19876 64220
rect 19580 64166 19626 64218
rect 19626 64166 19636 64218
rect 19660 64166 19690 64218
rect 19690 64166 19702 64218
rect 19702 64166 19716 64218
rect 19740 64166 19754 64218
rect 19754 64166 19766 64218
rect 19766 64166 19796 64218
rect 19820 64166 19830 64218
rect 19830 64166 19876 64218
rect 19580 64164 19636 64166
rect 19660 64164 19716 64166
rect 19740 64164 19796 64166
rect 19820 64164 19876 64166
rect 50300 64218 50356 64220
rect 50380 64218 50436 64220
rect 50460 64218 50516 64220
rect 50540 64218 50596 64220
rect 50300 64166 50346 64218
rect 50346 64166 50356 64218
rect 50380 64166 50410 64218
rect 50410 64166 50422 64218
rect 50422 64166 50436 64218
rect 50460 64166 50474 64218
rect 50474 64166 50486 64218
rect 50486 64166 50516 64218
rect 50540 64166 50550 64218
rect 50550 64166 50596 64218
rect 50300 64164 50356 64166
rect 50380 64164 50436 64166
rect 50460 64164 50516 64166
rect 50540 64164 50596 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 34940 63674 34996 63676
rect 35020 63674 35076 63676
rect 35100 63674 35156 63676
rect 35180 63674 35236 63676
rect 34940 63622 34986 63674
rect 34986 63622 34996 63674
rect 35020 63622 35050 63674
rect 35050 63622 35062 63674
rect 35062 63622 35076 63674
rect 35100 63622 35114 63674
rect 35114 63622 35126 63674
rect 35126 63622 35156 63674
rect 35180 63622 35190 63674
rect 35190 63622 35236 63674
rect 34940 63620 34996 63622
rect 35020 63620 35076 63622
rect 35100 63620 35156 63622
rect 35180 63620 35236 63622
rect 65660 63674 65716 63676
rect 65740 63674 65796 63676
rect 65820 63674 65876 63676
rect 65900 63674 65956 63676
rect 65660 63622 65706 63674
rect 65706 63622 65716 63674
rect 65740 63622 65770 63674
rect 65770 63622 65782 63674
rect 65782 63622 65796 63674
rect 65820 63622 65834 63674
rect 65834 63622 65846 63674
rect 65846 63622 65876 63674
rect 65900 63622 65910 63674
rect 65910 63622 65956 63674
rect 65660 63620 65716 63622
rect 65740 63620 65796 63622
rect 65820 63620 65876 63622
rect 65900 63620 65956 63622
rect 68466 63316 68468 63336
rect 68468 63316 68520 63336
rect 68520 63316 68522 63336
rect 68466 63280 68522 63316
rect 19580 63130 19636 63132
rect 19660 63130 19716 63132
rect 19740 63130 19796 63132
rect 19820 63130 19876 63132
rect 19580 63078 19626 63130
rect 19626 63078 19636 63130
rect 19660 63078 19690 63130
rect 19690 63078 19702 63130
rect 19702 63078 19716 63130
rect 19740 63078 19754 63130
rect 19754 63078 19766 63130
rect 19766 63078 19796 63130
rect 19820 63078 19830 63130
rect 19830 63078 19876 63130
rect 19580 63076 19636 63078
rect 19660 63076 19716 63078
rect 19740 63076 19796 63078
rect 19820 63076 19876 63078
rect 50300 63130 50356 63132
rect 50380 63130 50436 63132
rect 50460 63130 50516 63132
rect 50540 63130 50596 63132
rect 50300 63078 50346 63130
rect 50346 63078 50356 63130
rect 50380 63078 50410 63130
rect 50410 63078 50422 63130
rect 50422 63078 50436 63130
rect 50460 63078 50474 63130
rect 50474 63078 50486 63130
rect 50486 63078 50516 63130
rect 50540 63078 50550 63130
rect 50550 63078 50596 63130
rect 50300 63076 50356 63078
rect 50380 63076 50436 63078
rect 50460 63076 50516 63078
rect 50540 63076 50596 63078
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 34940 62586 34996 62588
rect 35020 62586 35076 62588
rect 35100 62586 35156 62588
rect 35180 62586 35236 62588
rect 34940 62534 34986 62586
rect 34986 62534 34996 62586
rect 35020 62534 35050 62586
rect 35050 62534 35062 62586
rect 35062 62534 35076 62586
rect 35100 62534 35114 62586
rect 35114 62534 35126 62586
rect 35126 62534 35156 62586
rect 35180 62534 35190 62586
rect 35190 62534 35236 62586
rect 34940 62532 34996 62534
rect 35020 62532 35076 62534
rect 35100 62532 35156 62534
rect 35180 62532 35236 62534
rect 65660 62586 65716 62588
rect 65740 62586 65796 62588
rect 65820 62586 65876 62588
rect 65900 62586 65956 62588
rect 65660 62534 65706 62586
rect 65706 62534 65716 62586
rect 65740 62534 65770 62586
rect 65770 62534 65782 62586
rect 65782 62534 65796 62586
rect 65820 62534 65834 62586
rect 65834 62534 65846 62586
rect 65846 62534 65876 62586
rect 65900 62534 65910 62586
rect 65910 62534 65956 62586
rect 65660 62532 65716 62534
rect 65740 62532 65796 62534
rect 65820 62532 65876 62534
rect 65900 62532 65956 62534
rect 19580 62042 19636 62044
rect 19660 62042 19716 62044
rect 19740 62042 19796 62044
rect 19820 62042 19876 62044
rect 19580 61990 19626 62042
rect 19626 61990 19636 62042
rect 19660 61990 19690 62042
rect 19690 61990 19702 62042
rect 19702 61990 19716 62042
rect 19740 61990 19754 62042
rect 19754 61990 19766 62042
rect 19766 61990 19796 62042
rect 19820 61990 19830 62042
rect 19830 61990 19876 62042
rect 19580 61988 19636 61990
rect 19660 61988 19716 61990
rect 19740 61988 19796 61990
rect 19820 61988 19876 61990
rect 50300 62042 50356 62044
rect 50380 62042 50436 62044
rect 50460 62042 50516 62044
rect 50540 62042 50596 62044
rect 50300 61990 50346 62042
rect 50346 61990 50356 62042
rect 50380 61990 50410 62042
rect 50410 61990 50422 62042
rect 50422 61990 50436 62042
rect 50460 61990 50474 62042
rect 50474 61990 50486 62042
rect 50486 61990 50516 62042
rect 50540 61990 50550 62042
rect 50550 61990 50596 62042
rect 50300 61988 50356 61990
rect 50380 61988 50436 61990
rect 50460 61988 50516 61990
rect 50540 61988 50596 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 65660 61498 65716 61500
rect 65740 61498 65796 61500
rect 65820 61498 65876 61500
rect 65900 61498 65956 61500
rect 65660 61446 65706 61498
rect 65706 61446 65716 61498
rect 65740 61446 65770 61498
rect 65770 61446 65782 61498
rect 65782 61446 65796 61498
rect 65820 61446 65834 61498
rect 65834 61446 65846 61498
rect 65846 61446 65876 61498
rect 65900 61446 65910 61498
rect 65910 61446 65956 61498
rect 65660 61444 65716 61446
rect 65740 61444 65796 61446
rect 65820 61444 65876 61446
rect 65900 61444 65956 61446
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 65660 60410 65716 60412
rect 65740 60410 65796 60412
rect 65820 60410 65876 60412
rect 65900 60410 65956 60412
rect 65660 60358 65706 60410
rect 65706 60358 65716 60410
rect 65740 60358 65770 60410
rect 65770 60358 65782 60410
rect 65782 60358 65796 60410
rect 65820 60358 65834 60410
rect 65834 60358 65846 60410
rect 65846 60358 65876 60410
rect 65900 60358 65910 60410
rect 65910 60358 65956 60410
rect 65660 60356 65716 60358
rect 65740 60356 65796 60358
rect 65820 60356 65876 60358
rect 65900 60356 65956 60358
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 65660 59322 65716 59324
rect 65740 59322 65796 59324
rect 65820 59322 65876 59324
rect 65900 59322 65956 59324
rect 65660 59270 65706 59322
rect 65706 59270 65716 59322
rect 65740 59270 65770 59322
rect 65770 59270 65782 59322
rect 65782 59270 65796 59322
rect 65820 59270 65834 59322
rect 65834 59270 65846 59322
rect 65846 59270 65876 59322
rect 65900 59270 65910 59322
rect 65910 59270 65956 59322
rect 65660 59268 65716 59270
rect 65740 59268 65796 59270
rect 65820 59268 65876 59270
rect 65900 59268 65956 59270
rect 1582 59200 1638 59256
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 65660 58234 65716 58236
rect 65740 58234 65796 58236
rect 65820 58234 65876 58236
rect 65900 58234 65956 58236
rect 65660 58182 65706 58234
rect 65706 58182 65716 58234
rect 65740 58182 65770 58234
rect 65770 58182 65782 58234
rect 65782 58182 65796 58234
rect 65820 58182 65834 58234
rect 65834 58182 65846 58234
rect 65846 58182 65876 58234
rect 65900 58182 65910 58234
rect 65910 58182 65956 58234
rect 65660 58180 65716 58182
rect 65740 58180 65796 58182
rect 65820 58180 65876 58182
rect 65900 58180 65956 58182
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 1582 56480 1638 56536
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 938 51040 994 51096
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 938 48320 994 48376
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 938 45600 994 45656
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 938 42880 994 42936
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 938 37440 994 37496
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 938 34720 994 34776
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 938 32000 994 32056
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 938 29280 994 29336
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 938 26560 994 26616
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 938 23840 994 23896
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 938 21120 994 21176
rect 938 18400 994 18456
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 938 15680 994 15736
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 938 12960 994 13016
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 938 10240 994 10296
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 938 7520 994 7576
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 31390 18692 31446 18728
rect 31390 18672 31392 18692
rect 31392 18672 31444 18692
rect 31444 18672 31446 18692
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 28814 6316 28870 6352
rect 28814 6296 28816 6316
rect 28816 6296 28868 6316
rect 28868 6296 28870 6316
rect 27710 3304 27766 3360
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 938 2080 994 2136
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 29458 5364 29514 5400
rect 29458 5344 29460 5364
rect 29460 5344 29512 5364
rect 29512 5344 29514 5364
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 42706 21548 42762 21584
rect 42706 21528 42708 21548
rect 42708 21528 42760 21548
rect 42760 21528 42762 21548
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 36818 18536 36874 18592
rect 30838 6296 30894 6352
rect 30838 5344 30894 5400
rect 33506 9424 33562 9480
rect 34426 15408 34482 15464
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 37922 18708 37924 18728
rect 37924 18708 37976 18728
rect 37976 18708 37978 18728
rect 37922 18672 37978 18708
rect 38474 18536 38530 18592
rect 38198 16516 38254 16552
rect 38198 16496 38200 16516
rect 38200 16496 38252 16516
rect 38252 16496 38254 16516
rect 37462 13776 37518 13832
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 39210 15428 39266 15464
rect 39210 15408 39212 15428
rect 39212 15408 39264 15428
rect 39264 15408 39266 15428
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38198 9460 38200 9480
rect 38200 9460 38252 9480
rect 38252 9460 38254 9480
rect 38198 9424 38254 9460
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38106 4004 38162 4040
rect 38106 3984 38108 4004
rect 38108 3984 38160 4004
rect 38160 3984 38162 4004
rect 45282 21392 45338 21448
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 41326 18284 41382 18320
rect 41326 18264 41328 18284
rect 41328 18264 41380 18284
rect 41380 18264 41382 18284
rect 41050 16108 41106 16144
rect 41050 16088 41052 16108
rect 41052 16088 41104 16108
rect 41104 16088 41106 16108
rect 44178 16088 44234 16144
rect 40590 10240 40646 10296
rect 45742 16496 45798 16552
rect 38566 3984 38622 4040
rect 44638 10240 44694 10296
rect 47674 21972 47676 21992
rect 47676 21972 47728 21992
rect 47728 21972 47730 21992
rect 47674 21936 47730 21972
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 48410 21956 48466 21992
rect 48410 21936 48412 21956
rect 48412 21936 48464 21956
rect 48464 21936 48466 21956
rect 46754 18536 46810 18592
rect 46938 18536 46994 18592
rect 46938 18264 46994 18320
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 68374 60580 68430 60616
rect 68374 60560 68376 60580
rect 68376 60560 68428 60580
rect 68428 60560 68430 60580
rect 68466 57876 68468 57896
rect 68468 57876 68520 57896
rect 68520 57876 68522 57896
rect 68466 57840 68522 57876
rect 68466 55140 68522 55176
rect 68466 55120 68468 55140
rect 68468 55120 68520 55140
rect 68520 55120 68522 55140
rect 68466 52436 68468 52456
rect 68468 52436 68520 52456
rect 68520 52436 68522 52456
rect 68466 52400 68522 52436
rect 68466 49716 68468 49736
rect 68468 49716 68520 49736
rect 68520 49716 68522 49736
rect 68466 49680 68522 49716
rect 68466 46996 68468 47016
rect 68468 46996 68520 47016
rect 68520 46996 68522 47016
rect 68466 46960 68522 46996
rect 68466 44260 68522 44296
rect 68466 44240 68468 44260
rect 68468 44240 68520 44260
rect 68520 44240 68522 44260
rect 68466 41556 68468 41576
rect 68468 41556 68520 41576
rect 68520 41556 68522 41576
rect 68466 41520 68522 41556
rect 68466 36116 68468 36136
rect 68468 36116 68520 36136
rect 68520 36116 68522 36136
rect 68466 36080 68522 36116
rect 68742 33360 68798 33416
rect 68466 30676 68468 30696
rect 68468 30676 68520 30696
rect 68520 30676 68522 30696
rect 68466 30640 68522 30676
rect 68466 27940 68522 27976
rect 68466 27920 68468 27940
rect 68468 27920 68520 27940
rect 68520 27920 68522 27940
rect 68466 25236 68468 25256
rect 68468 25236 68520 25256
rect 68520 25236 68522 25256
rect 68466 25200 68522 25236
rect 68466 22500 68522 22536
rect 68466 22480 68468 22500
rect 68468 22480 68520 22500
rect 68520 22480 68522 22500
rect 68374 21528 68430 21584
rect 68190 21392 68246 21448
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 47122 18264 47178 18320
rect 46478 15408 46534 15464
rect 47950 18264 48006 18320
rect 48778 18572 48780 18592
rect 48780 18572 48832 18592
rect 48832 18572 48834 18592
rect 48778 18536 48834 18572
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 68466 19796 68468 19816
rect 68468 19796 68520 19816
rect 68520 19796 68522 19816
rect 68466 19760 68522 19796
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 45374 7384 45430 7440
rect 48686 14900 48688 14920
rect 48688 14900 48740 14920
rect 48740 14900 48742 14920
rect 48686 14864 48742 14900
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 68466 17060 68522 17096
rect 68466 17040 68468 17060
rect 68468 17040 68520 17060
rect 68520 17040 68522 17060
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 52182 14864 52238 14920
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50342 11772 50344 11792
rect 50344 11772 50396 11792
rect 50396 11772 50398 11792
rect 50342 11736 50398 11772
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 68466 14356 68468 14376
rect 68468 14356 68520 14376
rect 68520 14356 68522 14376
rect 68466 14320 68522 14356
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 52182 11736 52238 11792
rect 68466 11620 68522 11656
rect 68466 11600 68468 11620
rect 68468 11600 68520 11620
rect 68520 11600 68522 11620
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 48134 7420 48136 7440
rect 48136 7420 48188 7440
rect 48188 7420 48190 7440
rect 48134 7384 48190 7420
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 68466 8916 68468 8936
rect 68468 8916 68520 8936
rect 68520 8916 68522 8936
rect 68466 8880 68522 8916
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 68466 6180 68522 6216
rect 68466 6160 68468 6180
rect 68468 6160 68520 6180
rect 68520 6160 68522 6180
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 68466 3476 68468 3496
rect 68468 3476 68520 3496
rect 68520 3476 68522 3496
rect 68466 3440 68522 3476
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 68650 720 68706 776
<< metal3 >>
rect 69200 68688 70000 68808
rect 19570 67488 19886 67489
rect 0 67418 800 67448
rect 19570 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19886 67488
rect 19570 67423 19886 67424
rect 50290 67488 50606 67489
rect 50290 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50606 67488
rect 50290 67423 50606 67424
rect 933 67418 999 67421
rect 0 67416 999 67418
rect 0 67360 938 67416
rect 994 67360 999 67416
rect 0 67358 999 67360
rect 0 67328 800 67358
rect 933 67355 999 67358
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 19570 66400 19886 66401
rect 19570 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19886 66400
rect 19570 66335 19886 66336
rect 50290 66400 50606 66401
rect 50290 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50606 66400
rect 50290 66335 50606 66336
rect 68461 66058 68527 66061
rect 69200 66058 70000 66088
rect 68461 66056 70000 66058
rect 68461 66000 68466 66056
rect 68522 66000 70000 66056
rect 68461 65998 70000 66000
rect 68461 65995 68527 65998
rect 69200 65968 70000 65998
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 19570 65312 19886 65313
rect 19570 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19886 65312
rect 19570 65247 19886 65248
rect 50290 65312 50606 65313
rect 50290 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50606 65312
rect 50290 65247 50606 65248
rect 1577 64834 1643 64837
rect 798 64832 1643 64834
rect 798 64776 1582 64832
rect 1638 64776 1643 64832
rect 798 64774 1643 64776
rect 798 64728 858 64774
rect 1577 64771 1643 64774
rect 0 64638 858 64728
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 34930 64768 35246 64769
rect 34930 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35246 64768
rect 34930 64703 35246 64704
rect 65650 64768 65966 64769
rect 65650 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65966 64768
rect 65650 64703 65966 64704
rect 0 64608 800 64638
rect 19570 64224 19886 64225
rect 19570 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19886 64224
rect 19570 64159 19886 64160
rect 50290 64224 50606 64225
rect 50290 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50606 64224
rect 50290 64159 50606 64160
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 34930 63680 35246 63681
rect 34930 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35246 63680
rect 34930 63615 35246 63616
rect 65650 63680 65966 63681
rect 65650 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65966 63680
rect 65650 63615 65966 63616
rect 68461 63338 68527 63341
rect 69200 63338 70000 63368
rect 68461 63336 70000 63338
rect 68461 63280 68466 63336
rect 68522 63280 70000 63336
rect 68461 63278 70000 63280
rect 68461 63275 68527 63278
rect 69200 63248 70000 63278
rect 19570 63136 19886 63137
rect 19570 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19886 63136
rect 19570 63071 19886 63072
rect 50290 63136 50606 63137
rect 50290 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50606 63136
rect 50290 63071 50606 63072
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 34930 62592 35246 62593
rect 34930 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35246 62592
rect 34930 62527 35246 62528
rect 65650 62592 65966 62593
rect 65650 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65966 62592
rect 65650 62527 65966 62528
rect 19570 62048 19886 62049
rect 0 61888 800 62008
rect 19570 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19886 62048
rect 19570 61983 19886 61984
rect 50290 62048 50606 62049
rect 50290 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50606 62048
rect 50290 61983 50606 61984
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 34930 61439 35246 61440
rect 65650 61504 65966 61505
rect 65650 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65966 61504
rect 65650 61439 65966 61440
rect 19570 60960 19886 60961
rect 19570 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19886 60960
rect 19570 60895 19886 60896
rect 50290 60960 50606 60961
rect 50290 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50606 60960
rect 50290 60895 50606 60896
rect 68369 60618 68435 60621
rect 69200 60618 70000 60648
rect 68369 60616 70000 60618
rect 68369 60560 68374 60616
rect 68430 60560 70000 60616
rect 68369 60558 70000 60560
rect 68369 60555 68435 60558
rect 69200 60528 70000 60558
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 34930 60351 35246 60352
rect 65650 60416 65966 60417
rect 65650 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65966 60416
rect 65650 60351 65966 60352
rect 19570 59872 19886 59873
rect 19570 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19886 59872
rect 19570 59807 19886 59808
rect 50290 59872 50606 59873
rect 50290 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50606 59872
rect 50290 59807 50606 59808
rect 4210 59328 4526 59329
rect 0 59258 800 59288
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 34930 59328 35246 59329
rect 34930 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35246 59328
rect 34930 59263 35246 59264
rect 65650 59328 65966 59329
rect 65650 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65966 59328
rect 65650 59263 65966 59264
rect 1577 59258 1643 59261
rect 0 59256 1643 59258
rect 0 59200 1582 59256
rect 1638 59200 1643 59256
rect 0 59198 1643 59200
rect 0 59168 800 59198
rect 1577 59195 1643 59198
rect 19570 58784 19886 58785
rect 19570 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19886 58784
rect 19570 58719 19886 58720
rect 50290 58784 50606 58785
rect 50290 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50606 58784
rect 50290 58719 50606 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 34930 58240 35246 58241
rect 34930 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35246 58240
rect 34930 58175 35246 58176
rect 65650 58240 65966 58241
rect 65650 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65966 58240
rect 65650 58175 65966 58176
rect 68461 57898 68527 57901
rect 69200 57898 70000 57928
rect 68461 57896 70000 57898
rect 68461 57840 68466 57896
rect 68522 57840 70000 57896
rect 68461 57838 70000 57840
rect 68461 57835 68527 57838
rect 69200 57808 70000 57838
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 19570 56608 19886 56609
rect 0 56538 800 56568
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 1577 56538 1643 56541
rect 0 56536 1643 56538
rect 0 56480 1582 56536
rect 1638 56480 1643 56536
rect 0 56478 1643 56480
rect 0 56448 800 56478
rect 1577 56475 1643 56478
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 65650 55999 65966 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 68461 55178 68527 55181
rect 69200 55178 70000 55208
rect 68461 55176 70000 55178
rect 68461 55120 68466 55176
rect 68522 55120 70000 55176
rect 68461 55118 70000 55120
rect 68461 55115 68527 55118
rect 69200 55088 70000 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 0 53728 800 53848
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 65650 53823 65966 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 68461 52458 68527 52461
rect 69200 52458 70000 52488
rect 68461 52456 70000 52458
rect 68461 52400 68466 52456
rect 68522 52400 70000 52456
rect 68461 52398 70000 52400
rect 68461 52395 68527 52398
rect 69200 52368 70000 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 19570 51168 19886 51169
rect 0 51098 800 51128
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 933 51098 999 51101
rect 0 51096 999 51098
rect 0 51040 938 51096
rect 994 51040 999 51096
rect 0 51038 999 51040
rect 0 51008 800 51038
rect 933 51035 999 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 68461 49738 68527 49741
rect 69200 49738 70000 49768
rect 68461 49736 70000 49738
rect 68461 49680 68466 49736
rect 68522 49680 70000 49736
rect 68461 49678 70000 49680
rect 68461 49675 68527 49678
rect 69200 49648 70000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 0 48378 800 48408
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 65650 48383 65966 48384
rect 933 48378 999 48381
rect 0 48376 999 48378
rect 0 48320 938 48376
rect 994 48320 999 48376
rect 0 48318 999 48320
rect 0 48288 800 48318
rect 933 48315 999 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 68461 47018 68527 47021
rect 69200 47018 70000 47048
rect 68461 47016 70000 47018
rect 68461 46960 68466 47016
rect 68522 46960 70000 47016
rect 68461 46958 70000 46960
rect 68461 46955 68527 46958
rect 69200 46928 70000 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 65650 46207 65966 46208
rect 19570 45728 19886 45729
rect 0 45658 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 933 45658 999 45661
rect 0 45656 999 45658
rect 0 45600 938 45656
rect 994 45600 999 45656
rect 0 45598 999 45600
rect 0 45568 800 45598
rect 933 45595 999 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 68461 44298 68527 44301
rect 69200 44298 70000 44328
rect 68461 44296 70000 44298
rect 68461 44240 68466 44296
rect 68522 44240 70000 44296
rect 68461 44238 70000 44240
rect 68461 44235 68527 44238
rect 69200 44208 70000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 65650 44031 65966 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 0 42938 800 42968
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 65650 42943 65966 42944
rect 933 42938 999 42941
rect 0 42936 999 42938
rect 0 42880 938 42936
rect 994 42880 999 42936
rect 0 42878 999 42880
rect 0 42848 800 42878
rect 933 42875 999 42878
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 68461 41578 68527 41581
rect 69200 41578 70000 41608
rect 68461 41576 70000 41578
rect 68461 41520 68466 41576
rect 68522 41520 70000 41576
rect 68461 41518 70000 41520
rect 68461 41515 68527 41518
rect 69200 41488 70000 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 19570 40288 19886 40289
rect 0 40128 800 40248
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 69200 38768 70000 38888
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 933 37498 999 37501
rect 0 37496 999 37498
rect 0 37440 938 37496
rect 994 37440 999 37496
rect 0 37438 999 37440
rect 0 37408 800 37438
rect 933 37435 999 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 68461 36138 68527 36141
rect 69200 36138 70000 36168
rect 68461 36136 70000 36138
rect 68461 36080 68466 36136
rect 68522 36080 70000 36136
rect 68461 36078 70000 36080
rect 68461 36075 68527 36078
rect 69200 36048 70000 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 19570 34848 19886 34849
rect 0 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 933 34778 999 34781
rect 0 34776 999 34778
rect 0 34720 938 34776
rect 994 34720 999 34776
rect 0 34718 999 34720
rect 0 34688 800 34718
rect 933 34715 999 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 68737 33418 68803 33421
rect 69200 33418 70000 33448
rect 68737 33416 70000 33418
rect 68737 33360 68742 33416
rect 68798 33360 70000 33416
rect 68737 33358 70000 33360
rect 68737 33355 68803 33358
rect 69200 33328 70000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 933 32058 999 32061
rect 0 32056 999 32058
rect 0 32000 938 32056
rect 994 32000 999 32056
rect 0 31998 999 32000
rect 0 31968 800 31998
rect 933 31995 999 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 68461 30698 68527 30701
rect 69200 30698 70000 30728
rect 68461 30696 70000 30698
rect 68461 30640 68466 30696
rect 68522 30640 70000 30696
rect 68461 30638 70000 30640
rect 68461 30635 68527 30638
rect 69200 30608 70000 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 19570 29408 19886 29409
rect 0 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 933 29338 999 29341
rect 0 29336 999 29338
rect 0 29280 938 29336
rect 994 29280 999 29336
rect 0 29278 999 29280
rect 0 29248 800 29278
rect 933 29275 999 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 68461 27978 68527 27981
rect 69200 27978 70000 28008
rect 68461 27976 70000 27978
rect 68461 27920 68466 27976
rect 68522 27920 70000 27976
rect 68461 27918 70000 27920
rect 68461 27915 68527 27918
rect 69200 27888 70000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 933 26618 999 26621
rect 0 26616 999 26618
rect 0 26560 938 26616
rect 994 26560 999 26616
rect 0 26558 999 26560
rect 0 26528 800 26558
rect 933 26555 999 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 68461 25258 68527 25261
rect 69200 25258 70000 25288
rect 68461 25256 70000 25258
rect 68461 25200 68466 25256
rect 68522 25200 70000 25256
rect 68461 25198 70000 25200
rect 68461 25195 68527 25198
rect 69200 25168 70000 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 19570 23968 19886 23969
rect 0 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 933 23898 999 23901
rect 0 23896 999 23898
rect 0 23840 938 23896
rect 994 23840 999 23896
rect 0 23838 999 23840
rect 0 23808 800 23838
rect 933 23835 999 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 68461 22538 68527 22541
rect 69200 22538 70000 22568
rect 68461 22536 70000 22538
rect 68461 22480 68466 22536
rect 68522 22480 70000 22536
rect 68461 22478 70000 22480
rect 68461 22475 68527 22478
rect 69200 22448 70000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 47669 21994 47735 21997
rect 48405 21994 48471 21997
rect 47669 21992 48471 21994
rect 47669 21936 47674 21992
rect 47730 21936 48410 21992
rect 48466 21936 48471 21992
rect 47669 21934 48471 21936
rect 47669 21931 47735 21934
rect 48405 21931 48471 21934
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 42701 21586 42767 21589
rect 68369 21586 68435 21589
rect 42701 21584 68435 21586
rect 42701 21528 42706 21584
rect 42762 21528 68374 21584
rect 68430 21528 68435 21584
rect 42701 21526 68435 21528
rect 42701 21523 42767 21526
rect 68369 21523 68435 21526
rect 45277 21450 45343 21453
rect 68185 21450 68251 21453
rect 45277 21448 68251 21450
rect 45277 21392 45282 21448
rect 45338 21392 68190 21448
rect 68246 21392 68251 21448
rect 45277 21390 68251 21392
rect 45277 21387 45343 21390
rect 68185 21387 68251 21390
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 68461 19818 68527 19821
rect 69200 19818 70000 19848
rect 68461 19816 70000 19818
rect 68461 19760 68466 19816
rect 68522 19760 70000 19816
rect 68461 19758 70000 19760
rect 68461 19755 68527 19758
rect 69200 19728 70000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 31385 18730 31451 18733
rect 37917 18730 37983 18733
rect 31385 18728 37983 18730
rect 31385 18672 31390 18728
rect 31446 18672 37922 18728
rect 37978 18672 37983 18728
rect 31385 18670 37983 18672
rect 31385 18667 31451 18670
rect 37917 18667 37983 18670
rect 36813 18594 36879 18597
rect 38469 18594 38535 18597
rect 36813 18592 38535 18594
rect 36813 18536 36818 18592
rect 36874 18536 38474 18592
rect 38530 18536 38535 18592
rect 36813 18534 38535 18536
rect 36813 18531 36879 18534
rect 38469 18531 38535 18534
rect 46749 18594 46815 18597
rect 46933 18594 46999 18597
rect 48773 18594 48839 18597
rect 46749 18592 48839 18594
rect 46749 18536 46754 18592
rect 46810 18536 46938 18592
rect 46994 18536 48778 18592
rect 48834 18536 48839 18592
rect 46749 18534 48839 18536
rect 46749 18531 46815 18534
rect 46933 18531 46999 18534
rect 48773 18531 48839 18534
rect 19570 18528 19886 18529
rect 0 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 41321 18322 41387 18325
rect 46933 18322 46999 18325
rect 41321 18320 46999 18322
rect 41321 18264 41326 18320
rect 41382 18264 46938 18320
rect 46994 18264 46999 18320
rect 41321 18262 46999 18264
rect 41321 18259 41387 18262
rect 46933 18259 46999 18262
rect 47117 18322 47183 18325
rect 47945 18322 48011 18325
rect 47117 18320 48011 18322
rect 47117 18264 47122 18320
rect 47178 18264 47950 18320
rect 48006 18264 48011 18320
rect 47117 18262 48011 18264
rect 47117 18259 47183 18262
rect 47945 18259 48011 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 68461 17098 68527 17101
rect 69200 17098 70000 17128
rect 68461 17096 70000 17098
rect 68461 17040 68466 17096
rect 68522 17040 70000 17096
rect 68461 17038 70000 17040
rect 68461 17035 68527 17038
rect 69200 17008 70000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 38193 16554 38259 16557
rect 45737 16554 45803 16557
rect 38193 16552 45803 16554
rect 38193 16496 38198 16552
rect 38254 16496 45742 16552
rect 45798 16496 45803 16552
rect 38193 16494 45803 16496
rect 38193 16491 38259 16494
rect 45737 16491 45803 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 41045 16146 41111 16149
rect 44173 16146 44239 16149
rect 41045 16144 44239 16146
rect 41045 16088 41050 16144
rect 41106 16088 44178 16144
rect 44234 16088 44239 16144
rect 41045 16086 44239 16088
rect 41045 16083 41111 16086
rect 44173 16083 44239 16086
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 34421 15466 34487 15469
rect 39205 15466 39271 15469
rect 46473 15466 46539 15469
rect 34421 15464 46539 15466
rect 34421 15408 34426 15464
rect 34482 15408 39210 15464
rect 39266 15408 46478 15464
rect 46534 15408 46539 15464
rect 34421 15406 46539 15408
rect 34421 15403 34487 15406
rect 39205 15403 39271 15406
rect 46473 15403 46539 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 48681 14922 48747 14925
rect 52177 14922 52243 14925
rect 48681 14920 52243 14922
rect 48681 14864 48686 14920
rect 48742 14864 52182 14920
rect 52238 14864 52243 14920
rect 48681 14862 52243 14864
rect 48681 14859 48747 14862
rect 52177 14859 52243 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 68461 14378 68527 14381
rect 69200 14378 70000 14408
rect 68461 14376 70000 14378
rect 68461 14320 68466 14376
rect 68522 14320 70000 14376
rect 68461 14318 70000 14320
rect 68461 14315 68527 14318
rect 69200 14288 70000 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 37457 13834 37523 13837
rect 37590 13834 37596 13836
rect 37457 13832 37596 13834
rect 37457 13776 37462 13832
rect 37518 13776 37596 13832
rect 37457 13774 37596 13776
rect 37457 13771 37523 13774
rect 37590 13772 37596 13774
rect 37660 13772 37666 13836
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 19570 13088 19886 13089
rect 0 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 50337 11794 50403 11797
rect 52177 11794 52243 11797
rect 50337 11792 52243 11794
rect 50337 11736 50342 11792
rect 50398 11736 52182 11792
rect 52238 11736 52243 11792
rect 50337 11734 52243 11736
rect 50337 11731 50403 11734
rect 52177 11731 52243 11734
rect 68461 11658 68527 11661
rect 69200 11658 70000 11688
rect 68461 11656 70000 11658
rect 68461 11600 68466 11656
rect 68522 11600 70000 11656
rect 68461 11598 70000 11600
rect 68461 11595 68527 11598
rect 69200 11568 70000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10208 800 10238
rect 933 10235 999 10238
rect 40585 10298 40651 10301
rect 44633 10298 44699 10301
rect 40585 10296 44699 10298
rect 40585 10240 40590 10296
rect 40646 10240 44638 10296
rect 44694 10240 44699 10296
rect 40585 10238 44699 10240
rect 40585 10235 40651 10238
rect 44633 10235 44699 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 33501 9482 33567 9485
rect 38193 9482 38259 9485
rect 33501 9480 38259 9482
rect 33501 9424 33506 9480
rect 33562 9424 38198 9480
rect 38254 9424 38259 9480
rect 33501 9422 38259 9424
rect 33501 9419 33567 9422
rect 38193 9419 38259 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 68461 8938 68527 8941
rect 69200 8938 70000 8968
rect 68461 8936 70000 8938
rect 68461 8880 68466 8936
rect 68522 8880 70000 8936
rect 68461 8878 70000 8880
rect 68461 8875 68527 8878
rect 69200 8848 70000 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 45369 7442 45435 7445
rect 48129 7442 48195 7445
rect 45369 7440 48195 7442
rect 45369 7384 45374 7440
rect 45430 7384 48134 7440
rect 48190 7384 48195 7440
rect 45369 7382 48195 7384
rect 45369 7379 45435 7382
rect 48129 7379 48195 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 28809 6354 28875 6357
rect 30833 6354 30899 6357
rect 28809 6352 30899 6354
rect 28809 6296 28814 6352
rect 28870 6296 30838 6352
rect 30894 6296 30899 6352
rect 28809 6294 30899 6296
rect 28809 6291 28875 6294
rect 30833 6291 30899 6294
rect 68461 6218 68527 6221
rect 69200 6218 70000 6248
rect 68461 6216 70000 6218
rect 68461 6160 68466 6216
rect 68522 6160 70000 6216
rect 68461 6158 70000 6160
rect 68461 6155 68527 6158
rect 69200 6128 70000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 29453 5402 29519 5405
rect 30833 5402 30899 5405
rect 29453 5400 30899 5402
rect 29453 5344 29458 5400
rect 29514 5344 30838 5400
rect 30894 5344 30899 5400
rect 29453 5342 30899 5344
rect 29453 5339 29519 5342
rect 30833 5339 30899 5342
rect 4210 4928 4526 4929
rect 0 4768 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 38101 4042 38167 4045
rect 38561 4042 38627 4045
rect 38101 4040 38627 4042
rect 38101 3984 38106 4040
rect 38162 3984 38566 4040
rect 38622 3984 38627 4040
rect 38101 3982 38627 3984
rect 38101 3979 38167 3982
rect 38561 3979 38627 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 68461 3498 68527 3501
rect 69200 3498 70000 3528
rect 68461 3496 70000 3498
rect 68461 3440 68466 3496
rect 68522 3440 70000 3496
rect 68461 3438 70000 3440
rect 68461 3435 68527 3438
rect 69200 3408 70000 3438
rect 27705 3362 27771 3365
rect 37590 3362 37596 3364
rect 27705 3360 37596 3362
rect 27705 3304 27710 3360
rect 27766 3304 37596 3360
rect 27705 3302 37596 3304
rect 27705 3299 27771 3302
rect 37590 3300 37596 3302
rect 37660 3300 37666 3364
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 19570 2208 19886 2209
rect 0 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 933 2138 999 2141
rect 0 2136 999 2138
rect 0 2080 938 2136
rect 994 2080 999 2136
rect 0 2078 999 2080
rect 0 2048 800 2078
rect 933 2075 999 2078
rect 68645 778 68711 781
rect 69200 778 70000 808
rect 68645 776 70000 778
rect 68645 720 68650 776
rect 68706 720 70000 776
rect 68645 718 70000 720
rect 68645 715 68711 718
rect 69200 688 70000 718
<< via3 >>
rect 19576 67484 19640 67488
rect 19576 67428 19580 67484
rect 19580 67428 19636 67484
rect 19636 67428 19640 67484
rect 19576 67424 19640 67428
rect 19656 67484 19720 67488
rect 19656 67428 19660 67484
rect 19660 67428 19716 67484
rect 19716 67428 19720 67484
rect 19656 67424 19720 67428
rect 19736 67484 19800 67488
rect 19736 67428 19740 67484
rect 19740 67428 19796 67484
rect 19796 67428 19800 67484
rect 19736 67424 19800 67428
rect 19816 67484 19880 67488
rect 19816 67428 19820 67484
rect 19820 67428 19876 67484
rect 19876 67428 19880 67484
rect 19816 67424 19880 67428
rect 50296 67484 50360 67488
rect 50296 67428 50300 67484
rect 50300 67428 50356 67484
rect 50356 67428 50360 67484
rect 50296 67424 50360 67428
rect 50376 67484 50440 67488
rect 50376 67428 50380 67484
rect 50380 67428 50436 67484
rect 50436 67428 50440 67484
rect 50376 67424 50440 67428
rect 50456 67484 50520 67488
rect 50456 67428 50460 67484
rect 50460 67428 50516 67484
rect 50516 67428 50520 67484
rect 50456 67424 50520 67428
rect 50536 67484 50600 67488
rect 50536 67428 50540 67484
rect 50540 67428 50596 67484
rect 50596 67428 50600 67484
rect 50536 67424 50600 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 19576 66396 19640 66400
rect 19576 66340 19580 66396
rect 19580 66340 19636 66396
rect 19636 66340 19640 66396
rect 19576 66336 19640 66340
rect 19656 66396 19720 66400
rect 19656 66340 19660 66396
rect 19660 66340 19716 66396
rect 19716 66340 19720 66396
rect 19656 66336 19720 66340
rect 19736 66396 19800 66400
rect 19736 66340 19740 66396
rect 19740 66340 19796 66396
rect 19796 66340 19800 66396
rect 19736 66336 19800 66340
rect 19816 66396 19880 66400
rect 19816 66340 19820 66396
rect 19820 66340 19876 66396
rect 19876 66340 19880 66396
rect 19816 66336 19880 66340
rect 50296 66396 50360 66400
rect 50296 66340 50300 66396
rect 50300 66340 50356 66396
rect 50356 66340 50360 66396
rect 50296 66336 50360 66340
rect 50376 66396 50440 66400
rect 50376 66340 50380 66396
rect 50380 66340 50436 66396
rect 50436 66340 50440 66396
rect 50376 66336 50440 66340
rect 50456 66396 50520 66400
rect 50456 66340 50460 66396
rect 50460 66340 50516 66396
rect 50516 66340 50520 66396
rect 50456 66336 50520 66340
rect 50536 66396 50600 66400
rect 50536 66340 50540 66396
rect 50540 66340 50596 66396
rect 50596 66340 50600 66396
rect 50536 66336 50600 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 19576 65308 19640 65312
rect 19576 65252 19580 65308
rect 19580 65252 19636 65308
rect 19636 65252 19640 65308
rect 19576 65248 19640 65252
rect 19656 65308 19720 65312
rect 19656 65252 19660 65308
rect 19660 65252 19716 65308
rect 19716 65252 19720 65308
rect 19656 65248 19720 65252
rect 19736 65308 19800 65312
rect 19736 65252 19740 65308
rect 19740 65252 19796 65308
rect 19796 65252 19800 65308
rect 19736 65248 19800 65252
rect 19816 65308 19880 65312
rect 19816 65252 19820 65308
rect 19820 65252 19876 65308
rect 19876 65252 19880 65308
rect 19816 65248 19880 65252
rect 50296 65308 50360 65312
rect 50296 65252 50300 65308
rect 50300 65252 50356 65308
rect 50356 65252 50360 65308
rect 50296 65248 50360 65252
rect 50376 65308 50440 65312
rect 50376 65252 50380 65308
rect 50380 65252 50436 65308
rect 50436 65252 50440 65308
rect 50376 65248 50440 65252
rect 50456 65308 50520 65312
rect 50456 65252 50460 65308
rect 50460 65252 50516 65308
rect 50516 65252 50520 65308
rect 50456 65248 50520 65252
rect 50536 65308 50600 65312
rect 50536 65252 50540 65308
rect 50540 65252 50596 65308
rect 50596 65252 50600 65308
rect 50536 65248 50600 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 34936 64764 35000 64768
rect 34936 64708 34940 64764
rect 34940 64708 34996 64764
rect 34996 64708 35000 64764
rect 34936 64704 35000 64708
rect 35016 64764 35080 64768
rect 35016 64708 35020 64764
rect 35020 64708 35076 64764
rect 35076 64708 35080 64764
rect 35016 64704 35080 64708
rect 35096 64764 35160 64768
rect 35096 64708 35100 64764
rect 35100 64708 35156 64764
rect 35156 64708 35160 64764
rect 35096 64704 35160 64708
rect 35176 64764 35240 64768
rect 35176 64708 35180 64764
rect 35180 64708 35236 64764
rect 35236 64708 35240 64764
rect 35176 64704 35240 64708
rect 65656 64764 65720 64768
rect 65656 64708 65660 64764
rect 65660 64708 65716 64764
rect 65716 64708 65720 64764
rect 65656 64704 65720 64708
rect 65736 64764 65800 64768
rect 65736 64708 65740 64764
rect 65740 64708 65796 64764
rect 65796 64708 65800 64764
rect 65736 64704 65800 64708
rect 65816 64764 65880 64768
rect 65816 64708 65820 64764
rect 65820 64708 65876 64764
rect 65876 64708 65880 64764
rect 65816 64704 65880 64708
rect 65896 64764 65960 64768
rect 65896 64708 65900 64764
rect 65900 64708 65956 64764
rect 65956 64708 65960 64764
rect 65896 64704 65960 64708
rect 19576 64220 19640 64224
rect 19576 64164 19580 64220
rect 19580 64164 19636 64220
rect 19636 64164 19640 64220
rect 19576 64160 19640 64164
rect 19656 64220 19720 64224
rect 19656 64164 19660 64220
rect 19660 64164 19716 64220
rect 19716 64164 19720 64220
rect 19656 64160 19720 64164
rect 19736 64220 19800 64224
rect 19736 64164 19740 64220
rect 19740 64164 19796 64220
rect 19796 64164 19800 64220
rect 19736 64160 19800 64164
rect 19816 64220 19880 64224
rect 19816 64164 19820 64220
rect 19820 64164 19876 64220
rect 19876 64164 19880 64220
rect 19816 64160 19880 64164
rect 50296 64220 50360 64224
rect 50296 64164 50300 64220
rect 50300 64164 50356 64220
rect 50356 64164 50360 64220
rect 50296 64160 50360 64164
rect 50376 64220 50440 64224
rect 50376 64164 50380 64220
rect 50380 64164 50436 64220
rect 50436 64164 50440 64220
rect 50376 64160 50440 64164
rect 50456 64220 50520 64224
rect 50456 64164 50460 64220
rect 50460 64164 50516 64220
rect 50516 64164 50520 64220
rect 50456 64160 50520 64164
rect 50536 64220 50600 64224
rect 50536 64164 50540 64220
rect 50540 64164 50596 64220
rect 50596 64164 50600 64220
rect 50536 64160 50600 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 34936 63676 35000 63680
rect 34936 63620 34940 63676
rect 34940 63620 34996 63676
rect 34996 63620 35000 63676
rect 34936 63616 35000 63620
rect 35016 63676 35080 63680
rect 35016 63620 35020 63676
rect 35020 63620 35076 63676
rect 35076 63620 35080 63676
rect 35016 63616 35080 63620
rect 35096 63676 35160 63680
rect 35096 63620 35100 63676
rect 35100 63620 35156 63676
rect 35156 63620 35160 63676
rect 35096 63616 35160 63620
rect 35176 63676 35240 63680
rect 35176 63620 35180 63676
rect 35180 63620 35236 63676
rect 35236 63620 35240 63676
rect 35176 63616 35240 63620
rect 65656 63676 65720 63680
rect 65656 63620 65660 63676
rect 65660 63620 65716 63676
rect 65716 63620 65720 63676
rect 65656 63616 65720 63620
rect 65736 63676 65800 63680
rect 65736 63620 65740 63676
rect 65740 63620 65796 63676
rect 65796 63620 65800 63676
rect 65736 63616 65800 63620
rect 65816 63676 65880 63680
rect 65816 63620 65820 63676
rect 65820 63620 65876 63676
rect 65876 63620 65880 63676
rect 65816 63616 65880 63620
rect 65896 63676 65960 63680
rect 65896 63620 65900 63676
rect 65900 63620 65956 63676
rect 65956 63620 65960 63676
rect 65896 63616 65960 63620
rect 19576 63132 19640 63136
rect 19576 63076 19580 63132
rect 19580 63076 19636 63132
rect 19636 63076 19640 63132
rect 19576 63072 19640 63076
rect 19656 63132 19720 63136
rect 19656 63076 19660 63132
rect 19660 63076 19716 63132
rect 19716 63076 19720 63132
rect 19656 63072 19720 63076
rect 19736 63132 19800 63136
rect 19736 63076 19740 63132
rect 19740 63076 19796 63132
rect 19796 63076 19800 63132
rect 19736 63072 19800 63076
rect 19816 63132 19880 63136
rect 19816 63076 19820 63132
rect 19820 63076 19876 63132
rect 19876 63076 19880 63132
rect 19816 63072 19880 63076
rect 50296 63132 50360 63136
rect 50296 63076 50300 63132
rect 50300 63076 50356 63132
rect 50356 63076 50360 63132
rect 50296 63072 50360 63076
rect 50376 63132 50440 63136
rect 50376 63076 50380 63132
rect 50380 63076 50436 63132
rect 50436 63076 50440 63132
rect 50376 63072 50440 63076
rect 50456 63132 50520 63136
rect 50456 63076 50460 63132
rect 50460 63076 50516 63132
rect 50516 63076 50520 63132
rect 50456 63072 50520 63076
rect 50536 63132 50600 63136
rect 50536 63076 50540 63132
rect 50540 63076 50596 63132
rect 50596 63076 50600 63132
rect 50536 63072 50600 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 34936 62588 35000 62592
rect 34936 62532 34940 62588
rect 34940 62532 34996 62588
rect 34996 62532 35000 62588
rect 34936 62528 35000 62532
rect 35016 62588 35080 62592
rect 35016 62532 35020 62588
rect 35020 62532 35076 62588
rect 35076 62532 35080 62588
rect 35016 62528 35080 62532
rect 35096 62588 35160 62592
rect 35096 62532 35100 62588
rect 35100 62532 35156 62588
rect 35156 62532 35160 62588
rect 35096 62528 35160 62532
rect 35176 62588 35240 62592
rect 35176 62532 35180 62588
rect 35180 62532 35236 62588
rect 35236 62532 35240 62588
rect 35176 62528 35240 62532
rect 65656 62588 65720 62592
rect 65656 62532 65660 62588
rect 65660 62532 65716 62588
rect 65716 62532 65720 62588
rect 65656 62528 65720 62532
rect 65736 62588 65800 62592
rect 65736 62532 65740 62588
rect 65740 62532 65796 62588
rect 65796 62532 65800 62588
rect 65736 62528 65800 62532
rect 65816 62588 65880 62592
rect 65816 62532 65820 62588
rect 65820 62532 65876 62588
rect 65876 62532 65880 62588
rect 65816 62528 65880 62532
rect 65896 62588 65960 62592
rect 65896 62532 65900 62588
rect 65900 62532 65956 62588
rect 65956 62532 65960 62588
rect 65896 62528 65960 62532
rect 19576 62044 19640 62048
rect 19576 61988 19580 62044
rect 19580 61988 19636 62044
rect 19636 61988 19640 62044
rect 19576 61984 19640 61988
rect 19656 62044 19720 62048
rect 19656 61988 19660 62044
rect 19660 61988 19716 62044
rect 19716 61988 19720 62044
rect 19656 61984 19720 61988
rect 19736 62044 19800 62048
rect 19736 61988 19740 62044
rect 19740 61988 19796 62044
rect 19796 61988 19800 62044
rect 19736 61984 19800 61988
rect 19816 62044 19880 62048
rect 19816 61988 19820 62044
rect 19820 61988 19876 62044
rect 19876 61988 19880 62044
rect 19816 61984 19880 61988
rect 50296 62044 50360 62048
rect 50296 61988 50300 62044
rect 50300 61988 50356 62044
rect 50356 61988 50360 62044
rect 50296 61984 50360 61988
rect 50376 62044 50440 62048
rect 50376 61988 50380 62044
rect 50380 61988 50436 62044
rect 50436 61988 50440 62044
rect 50376 61984 50440 61988
rect 50456 62044 50520 62048
rect 50456 61988 50460 62044
rect 50460 61988 50516 62044
rect 50516 61988 50520 62044
rect 50456 61984 50520 61988
rect 50536 62044 50600 62048
rect 50536 61988 50540 62044
rect 50540 61988 50596 62044
rect 50596 61988 50600 62044
rect 50536 61984 50600 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 65656 61500 65720 61504
rect 65656 61444 65660 61500
rect 65660 61444 65716 61500
rect 65716 61444 65720 61500
rect 65656 61440 65720 61444
rect 65736 61500 65800 61504
rect 65736 61444 65740 61500
rect 65740 61444 65796 61500
rect 65796 61444 65800 61500
rect 65736 61440 65800 61444
rect 65816 61500 65880 61504
rect 65816 61444 65820 61500
rect 65820 61444 65876 61500
rect 65876 61444 65880 61500
rect 65816 61440 65880 61444
rect 65896 61500 65960 61504
rect 65896 61444 65900 61500
rect 65900 61444 65956 61500
rect 65956 61444 65960 61500
rect 65896 61440 65960 61444
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 65656 60412 65720 60416
rect 65656 60356 65660 60412
rect 65660 60356 65716 60412
rect 65716 60356 65720 60412
rect 65656 60352 65720 60356
rect 65736 60412 65800 60416
rect 65736 60356 65740 60412
rect 65740 60356 65796 60412
rect 65796 60356 65800 60412
rect 65736 60352 65800 60356
rect 65816 60412 65880 60416
rect 65816 60356 65820 60412
rect 65820 60356 65876 60412
rect 65876 60356 65880 60412
rect 65816 60352 65880 60356
rect 65896 60412 65960 60416
rect 65896 60356 65900 60412
rect 65900 60356 65956 60412
rect 65956 60356 65960 60412
rect 65896 60352 65960 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 65656 59324 65720 59328
rect 65656 59268 65660 59324
rect 65660 59268 65716 59324
rect 65716 59268 65720 59324
rect 65656 59264 65720 59268
rect 65736 59324 65800 59328
rect 65736 59268 65740 59324
rect 65740 59268 65796 59324
rect 65796 59268 65800 59324
rect 65736 59264 65800 59268
rect 65816 59324 65880 59328
rect 65816 59268 65820 59324
rect 65820 59268 65876 59324
rect 65876 59268 65880 59324
rect 65816 59264 65880 59268
rect 65896 59324 65960 59328
rect 65896 59268 65900 59324
rect 65900 59268 65956 59324
rect 65956 59268 65960 59324
rect 65896 59264 65960 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 65656 58236 65720 58240
rect 65656 58180 65660 58236
rect 65660 58180 65716 58236
rect 65716 58180 65720 58236
rect 65656 58176 65720 58180
rect 65736 58236 65800 58240
rect 65736 58180 65740 58236
rect 65740 58180 65796 58236
rect 65796 58180 65800 58236
rect 65736 58176 65800 58180
rect 65816 58236 65880 58240
rect 65816 58180 65820 58236
rect 65820 58180 65876 58236
rect 65876 58180 65880 58236
rect 65816 58176 65880 58180
rect 65896 58236 65960 58240
rect 65896 58180 65900 58236
rect 65900 58180 65956 58236
rect 65956 58180 65960 58236
rect 65896 58176 65960 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 37596 13772 37660 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 37596 3300 37660 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 66944 4528 67504
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 65856 4528 66880
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 67488 19888 67504
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 66400 19888 67424
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 65312 19888 66336
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 64224 19888 65248
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 63136 19888 64160
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 62048 19888 63072
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 60960 19888 61984
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 66944 35248 67504
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 65856 35248 66880
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 64768 35248 65792
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 63680 35248 64704
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 62592 35248 63616
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 61504 35248 62528
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 50288 67488 50608 67504
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 66400 50608 67424
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 65312 50608 66336
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 64224 50608 65248
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 63136 50608 64160
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 62048 50608 63072
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 60960 50608 61984
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 37595 13836 37661 13837
rect 37595 13772 37596 13836
rect 37660 13772 37661 13836
rect 37595 13771 37661 13772
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 37598 3365 37658 13771
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 37595 3364 37661 3365
rect 37595 3300 37596 3364
rect 37660 3300 37661 3364
rect 37595 3299 37661 3300
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 66944 65968 67504
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 65856 65968 66880
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 64768 65968 65792
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 63680 65968 64704
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 62592 65968 63616
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 61504 65968 62528
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 60416 65968 61440
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 59328 65968 60352
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 58240 65968 59264
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 57152 65968 58176
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__or4b_1  _0611_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0612_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47840 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0613_
timestamp 1688980957
transform 1 0 46736 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0614_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46276 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0615_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46460 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0616_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 48576 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0617_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 48852 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0618_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47012 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0619_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47196 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0620_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46092 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0621_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 45816 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0622_
timestamp 1688980957
transform 1 0 46828 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0623_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46460 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0624_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46184 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0625_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0626_
timestamp 1688980957
transform 1 0 46920 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1688980957
transform 1 0 46828 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0628_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47288 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0629_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46000 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0630_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0631_
timestamp 1688980957
transform 1 0 48392 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0632_
timestamp 1688980957
transform 1 0 47840 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1688980957
transform 1 0 48760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0634_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 50140 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0635_
timestamp 1688980957
transform 1 0 49220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0636_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 50048 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0637_
timestamp 1688980957
transform 1 0 50140 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0638_
timestamp 1688980957
transform 1 0 49312 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0639_
timestamp 1688980957
transform 1 0 47564 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0640_
timestamp 1688980957
transform 1 0 48668 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0641_
timestamp 1688980957
transform 1 0 46736 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform 1 0 50140 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1688980957
transform 1 0 49220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0644_
timestamp 1688980957
transform 1 0 45172 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0645_
timestamp 1688980957
transform 1 0 44712 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _0646_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 45816 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0647_
timestamp 1688980957
transform 1 0 45540 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0648_
timestamp 1688980957
transform 1 0 48024 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0649_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44988 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0650_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46276 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0651_
timestamp 1688980957
transform 1 0 45816 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0652_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0653_
timestamp 1688980957
transform 1 0 49036 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0654_
timestamp 1688980957
transform 1 0 50600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0655_
timestamp 1688980957
transform 1 0 49680 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0656_
timestamp 1688980957
transform 1 0 49036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0657_
timestamp 1688980957
transform 1 0 48392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0658_
timestamp 1688980957
transform 1 0 49496 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0659_
timestamp 1688980957
transform 1 0 51060 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0660_
timestamp 1688980957
transform 1 0 50876 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0661_
timestamp 1688980957
transform 1 0 51244 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0662_
timestamp 1688980957
transform 1 0 52624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0663_
timestamp 1688980957
transform 1 0 48300 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0664_
timestamp 1688980957
transform 1 0 52164 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1688980957
transform 1 0 52348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0666_
timestamp 1688980957
transform 1 0 51704 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0667_
timestamp 1688980957
transform 1 0 51428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0668_
timestamp 1688980957
transform 1 0 48576 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0669_
timestamp 1688980957
transform 1 0 51980 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0670_
timestamp 1688980957
transform 1 0 51520 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0671_
timestamp 1688980957
transform 1 0 51888 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1688980957
transform 1 0 50692 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0673_
timestamp 1688980957
transform 1 0 49496 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0674_
timestamp 1688980957
transform 1 0 51336 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1688980957
transform 1 0 51520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0676_
timestamp 1688980957
transform 1 0 50140 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0677_
timestamp 1688980957
transform 1 0 49496 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0678_
timestamp 1688980957
transform 1 0 52716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0679_
timestamp 1688980957
transform 1 0 51980 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0680_
timestamp 1688980957
transform 1 0 51244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0681_
timestamp 1688980957
transform 1 0 48944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0682_
timestamp 1688980957
transform 1 0 47564 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0683_
timestamp 1688980957
transform 1 0 47932 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1688980957
transform 1 0 47288 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1688980957
transform 1 0 38732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0686_
timestamp 1688980957
transform 1 0 39560 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0687_
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0688_
timestamp 1688980957
transform 1 0 41124 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0689_
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0690_
timestamp 1688980957
transform 1 0 37812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0691_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38640 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0692_
timestamp 1688980957
transform 1 0 38916 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0693_
timestamp 1688980957
transform 1 0 39008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0694_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44896 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1688980957
transform 1 0 45724 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0696_
timestamp 1688980957
transform 1 0 45908 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1688980957
transform 1 0 47748 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0698_
timestamp 1688980957
transform 1 0 48208 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0699_
timestamp 1688980957
transform 1 0 49680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0700_
timestamp 1688980957
transform 1 0 45540 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0701_
timestamp 1688980957
transform 1 0 49220 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0702_
timestamp 1688980957
transform 1 0 48668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0703_
timestamp 1688980957
transform 1 0 48576 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0704_
timestamp 1688980957
transform 1 0 47656 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1688980957
transform 1 0 47472 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0706_
timestamp 1688980957
transform 1 0 49588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0707_
timestamp 1688980957
transform 1 0 45080 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0708_
timestamp 1688980957
transform 1 0 47748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1688980957
transform 1 0 48760 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0710_
timestamp 1688980957
transform 1 0 49588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0711_
timestamp 1688980957
transform 1 0 48208 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0712_
timestamp 1688980957
transform 1 0 49036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1688980957
transform 1 0 46368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0714_
timestamp 1688980957
transform 1 0 46460 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0715_
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0716_
timestamp 1688980957
transform 1 0 48300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0717_
timestamp 1688980957
transform 1 0 46828 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0718_
timestamp 1688980957
transform 1 0 46092 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0719_
timestamp 1688980957
transform 1 0 46644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0720_
timestamp 1688980957
transform 1 0 46552 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1688980957
transform 1 0 45264 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 1688980957
transform 1 0 43976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 1688980957
transform 1 0 33304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1688980957
transform 1 0 32844 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0727_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1688980957
transform 1 0 27692 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0729_
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0730_
timestamp 1688980957
transform 1 0 27140 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0732_
timestamp 1688980957
transform 1 0 33028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1688980957
transform 1 0 40388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0734_
timestamp 1688980957
transform 1 0 37628 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1688980957
transform 1 0 39376 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 1688980957
transform 1 0 39376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0737_
timestamp 1688980957
transform 1 0 40480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0738_
timestamp 1688980957
transform 1 0 40388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0739_
timestamp 1688980957
transform 1 0 39284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0740_
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0741_
timestamp 1688980957
transform 1 0 40020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1688980957
transform 1 0 40756 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 1688980957
transform 1 0 41308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0744_
timestamp 1688980957
transform 1 0 40572 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0745_
timestamp 1688980957
transform 1 0 40756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0746_
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0747_
timestamp 1688980957
transform 1 0 39284 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0748_
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0749_
timestamp 1688980957
transform 1 0 39100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0750_
timestamp 1688980957
transform 1 0 39100 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0751_
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0752_
timestamp 1688980957
transform 1 0 38272 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0753_
timestamp 1688980957
transform 1 0 37536 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1688980957
transform 1 0 36340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0755_
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0756_
timestamp 1688980957
transform 1 0 36248 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0757_
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0758_
timestamp 1688980957
transform 1 0 35880 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1688980957
transform 1 0 37536 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0760_
timestamp 1688980957
transform 1 0 36064 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0761_
timestamp 1688980957
transform 1 0 35880 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0762_
timestamp 1688980957
transform 1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0763_
timestamp 1688980957
transform 1 0 33580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1688980957
transform 1 0 33304 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0765_
timestamp 1688980957
transform 1 0 31556 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1688980957
transform 1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0767_
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0768_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0769_
timestamp 1688980957
transform 1 0 31004 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0770_
timestamp 1688980957
transform 1 0 31096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0771_
timestamp 1688980957
transform 1 0 33028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0772_
timestamp 1688980957
transform 1 0 28520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0773_
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0774_
timestamp 1688980957
transform 1 0 25668 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 1688980957
transform 1 0 26496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0776_
timestamp 1688980957
transform 1 0 27232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1688980957
transform 1 0 26404 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0778_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _0779_
timestamp 1688980957
transform 1 0 26956 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0780_
timestamp 1688980957
transform 1 0 26220 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1688980957
transform 1 0 26772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0782_
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0783_
timestamp 1688980957
transform 1 0 25760 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0784_
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0785_
timestamp 1688980957
transform 1 0 26128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0786_
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0787_
timestamp 1688980957
transform 1 0 25944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0788_
timestamp 1688980957
transform 1 0 24472 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1688980957
transform 1 0 25760 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0790_
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0791_
timestamp 1688980957
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1688980957
transform 1 0 24748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0793_
timestamp 1688980957
transform 1 0 25392 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0794_
timestamp 1688980957
transform 1 0 24380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0795_
timestamp 1688980957
transform 1 0 24840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0796_
timestamp 1688980957
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0797_
timestamp 1688980957
transform 1 0 24472 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0798_
timestamp 1688980957
transform 1 0 26496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0799_
timestamp 1688980957
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1688980957
transform 1 0 24748 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 1688980957
transform 1 0 23368 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0802_
timestamp 1688980957
transform 1 0 30544 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0803_
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0804_
timestamp 1688980957
transform 1 0 27968 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0805_
timestamp 1688980957
transform 1 0 28888 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1688980957
transform 1 0 31556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0807_
timestamp 1688980957
transform 1 0 31556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0808_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0809_
timestamp 1688980957
transform 1 0 28428 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0811_
timestamp 1688980957
transform 1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0812_
timestamp 1688980957
transform 1 0 28612 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 1688980957
transform 1 0 28336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1688980957
transform 1 0 28060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1688980957
transform 1 0 31556 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0816_
timestamp 1688980957
transform 1 0 28336 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1688980957
transform 1 0 27232 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0818_
timestamp 1688980957
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1688980957
transform 1 0 29348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0820_
timestamp 1688980957
transform 1 0 28888 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0821_
timestamp 1688980957
transform 1 0 27048 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0822_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0823_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28060 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1688980957
transform 1 0 29992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0825_
timestamp 1688980957
transform 1 0 30544 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0826_
timestamp 1688980957
transform 1 0 29808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1688980957
transform 1 0 32844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0828_
timestamp 1688980957
transform 1 0 32108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1688980957
transform 1 0 31188 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0830_
timestamp 1688980957
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0831_
timestamp 1688980957
transform 1 0 44988 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1688980957
transform 1 0 45356 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1688980957
transform 1 0 44620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0834_
timestamp 1688980957
transform 1 0 44988 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 1688980957
transform 1 0 46460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0836_
timestamp 1688980957
transform 1 0 46000 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0837_
timestamp 1688980957
transform 1 0 45540 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1688980957
transform 1 0 34960 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0839_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0840_
timestamp 1688980957
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0841_
timestamp 1688980957
transform 1 0 31004 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1688980957
transform 1 0 39652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0843_
timestamp 1688980957
transform 1 0 29900 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0844_
timestamp 1688980957
transform 1 0 44252 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0845_
timestamp 1688980957
transform 1 0 38640 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0846_
timestamp 1688980957
transform 1 0 39284 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0847_
timestamp 1688980957
transform 1 0 30544 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0848_
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1688980957
transform 1 0 33856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0851_
timestamp 1688980957
transform 1 0 33120 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1688980957
transform 1 0 43608 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0853_
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0854_
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0855_
timestamp 1688980957
transform 1 0 39744 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0856_
timestamp 1688980957
transform 1 0 39652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0857_
timestamp 1688980957
transform 1 0 38364 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0858_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0859_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43884 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0860_
timestamp 1688980957
transform 1 0 42412 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1688980957
transform 1 0 43884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1688980957
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1688980957
transform 1 0 34224 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0864_
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1688980957
transform 1 0 41952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0866_
timestamp 1688980957
transform 1 0 40204 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1688980957
transform 1 0 41308 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0868_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40940 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1688980957
transform 1 0 40664 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0870_
timestamp 1688980957
transform 1 0 42320 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0871_
timestamp 1688980957
transform 1 0 43056 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0872_
timestamp 1688980957
transform 1 0 38456 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0873_
timestamp 1688980957
transform 1 0 34224 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0874_
timestamp 1688980957
transform 1 0 33580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0875_
timestamp 1688980957
transform 1 0 38916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0876_
timestamp 1688980957
transform 1 0 36800 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0877_
timestamp 1688980957
transform 1 0 36340 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0879_
timestamp 1688980957
transform 1 0 43700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0880_
timestamp 1688980957
transform 1 0 45724 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0881_
timestamp 1688980957
transform 1 0 45080 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0882_
timestamp 1688980957
transform 1 0 43516 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0883_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27048 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0884_
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0885_
timestamp 1688980957
transform 1 0 30544 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0886_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28520 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0887_
timestamp 1688980957
transform 1 0 28520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0888_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 1688980957
transform 1 0 28980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0890_
timestamp 1688980957
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0891_
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1688980957
transform 1 0 32292 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0894_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33304 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0895_
timestamp 1688980957
transform 1 0 34224 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0896_
timestamp 1688980957
transform 1 0 31280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0897_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33120 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0898_
timestamp 1688980957
transform 1 0 37996 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1688980957
transform 1 0 37076 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_2  _0900_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37812 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0901_
timestamp 1688980957
transform 1 0 37996 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 1688980957
transform 1 0 36800 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0903_
timestamp 1688980957
transform 1 0 36340 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1688980957
transform 1 0 35052 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1688980957
transform 1 0 35512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0906_
timestamp 1688980957
transform 1 0 38548 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0907_
timestamp 1688980957
transform 1 0 37628 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0908_
timestamp 1688980957
transform 1 0 39100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0909_
timestamp 1688980957
transform 1 0 36248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0910_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0911_
timestamp 1688980957
transform 1 0 40664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1688980957
transform 1 0 39376 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0913_
timestamp 1688980957
transform 1 0 32016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1688980957
transform 1 0 29624 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0915_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 1688980957
transform 1 0 33856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1688980957
transform 1 0 32844 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0918_
timestamp 1688980957
transform 1 0 32660 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 1688980957
transform 1 0 40664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0920_
timestamp 1688980957
transform 1 0 41768 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0921_
timestamp 1688980957
transform 1 0 40572 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0922_
timestamp 1688980957
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0923_
timestamp 1688980957
transform 1 0 29808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0924_
timestamp 1688980957
transform 1 0 40296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1688980957
transform 1 0 39192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1688980957
transform 1 0 39468 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0927_
timestamp 1688980957
transform 1 0 39284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0928_
timestamp 1688980957
transform 1 0 34132 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp 1688980957
transform 1 0 26956 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0930_
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1688980957
transform 1 0 25944 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0932_
timestamp 1688980957
transform 1 0 36340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0933_
timestamp 1688980957
transform 1 0 37904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0934_
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0935_
timestamp 1688980957
transform 1 0 37720 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0936_
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0937_
timestamp 1688980957
transform 1 0 35052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 1688980957
transform 1 0 45172 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 1688980957
transform 1 0 44620 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1688980957
transform 1 0 37812 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0941_
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1688980957
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0944_
timestamp 1688980957
transform 1 0 44344 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp 1688980957
transform 1 0 43792 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 1688980957
transform 1 0 38640 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0947_
timestamp 1688980957
transform 1 0 33580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 1688980957
transform 1 0 33028 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0949_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 1688980957
transform 1 0 25392 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_1  _0951_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26036 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0952_
timestamp 1688980957
transform 1 0 28244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0953_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0954_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0955_
timestamp 1688980957
transform 1 0 37260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1688980957
transform 1 0 36064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0957_
timestamp 1688980957
transform 1 0 35788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0958_
timestamp 1688980957
transform 1 0 35512 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0959_
timestamp 1688980957
transform 1 0 36340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0960_
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0961_
timestamp 1688980957
transform 1 0 38180 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0962_
timestamp 1688980957
transform 1 0 51520 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1688980957
transform 1 0 47656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1688980957
transform 1 0 48208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0965_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 48300 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0966_
timestamp 1688980957
transform 1 0 49312 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0967_
timestamp 1688980957
transform 1 0 49864 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0968_
timestamp 1688980957
transform 1 0 49036 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _0969_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1688980957
transform 1 0 47288 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1688980957
transform 1 0 46736 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0972_
timestamp 1688980957
transform 1 0 46736 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0973_
timestamp 1688980957
transform 1 0 47472 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 1688980957
transform 1 0 47472 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0975_
timestamp 1688980957
transform 1 0 48484 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0976_
timestamp 1688980957
transform 1 0 47656 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _0977_
timestamp 1688980957
transform 1 0 46460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1688980957
transform 1 0 46552 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0979_
timestamp 1688980957
transform 1 0 44344 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _0980_
timestamp 1688980957
transform 1 0 46000 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0981_
timestamp 1688980957
transform 1 0 46368 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0982_
timestamp 1688980957
transform 1 0 45816 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0983_
timestamp 1688980957
transform 1 0 45632 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0984_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 45908 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0985_
timestamp 1688980957
transform 1 0 37352 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _0986_
timestamp 1688980957
transform 1 0 29716 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1688980957
transform 1 0 30912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0988_
timestamp 1688980957
transform 1 0 30544 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0989_
timestamp 1688980957
transform 1 0 29716 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _0990_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29992 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0991_
timestamp 1688980957
transform 1 0 30360 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _0992_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1688980957
transform 1 0 30820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 1688980957
transform 1 0 28704 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1688980957
transform 1 0 29532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0997_
timestamp 1688980957
transform 1 0 37812 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1688980957
transform 1 0 39376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp 1688980957
transform 1 0 43240 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1688980957
transform 1 0 42688 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 1688980957
transform 1 0 48392 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1688980957
transform 1 0 48208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1003_
timestamp 1688980957
transform 1 0 42964 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1688980957
transform 1 0 42412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1688980957
transform 1 0 31556 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1688980957
transform 1 0 33580 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1007_
timestamp 1688980957
transform 1 0 31556 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1009_
timestamp 1688980957
transform 1 0 39100 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _1011_
timestamp 1688980957
transform 1 0 40112 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1012_
timestamp 1688980957
transform 1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1013_
timestamp 1688980957
transform 1 0 28704 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1015_
timestamp 1688980957
transform 1 0 27784 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1688980957
transform 1 0 29348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1017_
timestamp 1688980957
transform 1 0 40296 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1688980957
transform 1 0 40020 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1019_
timestamp 1688980957
transform 1 0 41768 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1688980957
transform 1 0 41216 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1021_
timestamp 1688980957
transform 1 0 32844 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1688980957
transform 1 0 32568 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1023_
timestamp 1688980957
transform 1 0 33948 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1688980957
transform 1 0 34776 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1025_
timestamp 1688980957
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1688980957
transform 1 0 30820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1027_
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1028_
timestamp 1688980957
transform 1 0 38364 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1688980957
transform 1 0 39008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 1688980957
transform 1 0 35880 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1688980957
transform 1 0 37628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1032_
timestamp 1688980957
transform 1 0 43240 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1033_
timestamp 1688980957
transform 1 0 48116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1034_
timestamp 1688980957
transform 1 0 43792 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1035_
timestamp 1688980957
transform 1 0 37444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1036_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38548 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1037_
timestamp 1688980957
transform 1 0 40296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1038_
timestamp 1688980957
transform 1 0 39192 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1039_
timestamp 1688980957
transform 1 0 38732 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1040_
timestamp 1688980957
transform 1 0 37076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1041_
timestamp 1688980957
transform 1 0 36524 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1042_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1043_
timestamp 1688980957
transform 1 0 36800 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1044_
timestamp 1688980957
transform 1 0 37352 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1045_
timestamp 1688980957
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1046_
timestamp 1688980957
transform 1 0 37904 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1047_
timestamp 1688980957
transform 1 0 38640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1688980957
transform 1 0 35512 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1049_
timestamp 1688980957
transform 1 0 36064 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1050_
timestamp 1688980957
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1051_
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1052_
timestamp 1688980957
transform 1 0 34224 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1053_
timestamp 1688980957
transform 1 0 36064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1054_
timestamp 1688980957
transform 1 0 36064 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1055_
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1056_
timestamp 1688980957
transform 1 0 34684 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1057_
timestamp 1688980957
transform 1 0 36616 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1058_
timestamp 1688980957
transform 1 0 36524 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1059_
timestamp 1688980957
transform 1 0 37720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1060_
timestamp 1688980957
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1061_
timestamp 1688980957
transform 1 0 39284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1062_
timestamp 1688980957
transform 1 0 36064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1063_
timestamp 1688980957
transform 1 0 35696 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1688980957
transform 1 0 33948 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1065_
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1066_
timestamp 1688980957
transform 1 0 33580 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1067_
timestamp 1688980957
transform 1 0 31556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 1688980957
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1069_
timestamp 1688980957
transform 1 0 31280 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 1688980957
transform 1 0 32200 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1071_
timestamp 1688980957
transform 1 0 33764 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1072_
timestamp 1688980957
transform 1 0 32844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1073_
timestamp 1688980957
transform 1 0 38732 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1074_
timestamp 1688980957
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1075_
timestamp 1688980957
transform 1 0 47012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1076_
timestamp 1688980957
transform 1 0 46276 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1077_
timestamp 1688980957
transform 1 0 47012 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1078_
timestamp 1688980957
transform 1 0 33120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1079_
timestamp 1688980957
transform 1 0 33396 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1080_
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1081_
timestamp 1688980957
transform 1 0 28704 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1082_
timestamp 1688980957
transform 1 0 29072 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1083_
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1084_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1085_
timestamp 1688980957
transform 1 0 31004 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1086_
timestamp 1688980957
transform 1 0 30360 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1087_
timestamp 1688980957
transform 1 0 31464 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1088_
timestamp 1688980957
transform 1 0 32568 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1089_
timestamp 1688980957
transform 1 0 31280 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1090_
timestamp 1688980957
transform 1 0 33028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1091_
timestamp 1688980957
transform 1 0 32016 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _1092_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31280 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1094_
timestamp 1688980957
transform 1 0 29808 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1095_
timestamp 1688980957
transform 1 0 30728 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1096_
timestamp 1688980957
transform 1 0 30636 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1097_
timestamp 1688980957
transform 1 0 30084 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1098_
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1099_
timestamp 1688980957
transform 1 0 30268 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1688980957
transform 1 0 28704 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1101_
timestamp 1688980957
transform 1 0 28796 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1102_
timestamp 1688980957
transform 1 0 29348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1103_
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1104_
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1105_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1106_
timestamp 1688980957
transform 1 0 28336 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1107_
timestamp 1688980957
transform 1 0 29440 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1108_
timestamp 1688980957
transform 1 0 28796 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1688980957
transform 1 0 30452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1110_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 1688980957
transform 1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1112_
timestamp 1688980957
transform 1 0 27692 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1113_
timestamp 1688980957
transform 1 0 26956 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1114_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1688980957
transform 1 0 26128 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1116_
timestamp 1688980957
transform 1 0 26404 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1117_
timestamp 1688980957
transform 1 0 26312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1118_
timestamp 1688980957
transform 1 0 25392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1119_
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1120_
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1121_
timestamp 1688980957
transform 1 0 37444 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1688980957
transform 1 0 37996 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1123_
timestamp 1688980957
transform 1 0 43332 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1124_
timestamp 1688980957
transform 1 0 44344 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1688980957
transform 1 0 38088 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1688980957
transform 1 0 32936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1688980957
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1688980957
transform 1 0 28428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1688980957
transform 1 0 26404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1688980957
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1134_
timestamp 1688980957
transform 1 0 32568 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1688980957
transform 1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1137_
timestamp 1688980957
transform 1 0 31188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1138_
timestamp 1688980957
transform 1 0 31280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1688980957
transform 1 0 31556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1140_
timestamp 1688980957
transform 1 0 30452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1688980957
transform 1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 1688980957
transform 1 0 26496 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1688980957
transform 1 0 23552 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1688980957
transform 1 0 23460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1688980957
transform 1 0 23552 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1149_
timestamp 1688980957
transform 1 0 37996 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1150_
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1688980957
transform 1 0 31096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1152_
timestamp 1688980957
transform 1 0 27416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1153_
timestamp 1688980957
transform 1 0 27784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1155_
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1156_
timestamp 1688980957
transform 1 0 29624 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1157_
timestamp 1688980957
transform 1 0 30912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1158_
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1159_
timestamp 1688980957
transform 1 0 33764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1688980957
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1688980957
transform 1 0 34960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1163_
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1688980957
transform 1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1688980957
transform 1 0 41032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1688980957
transform 1 0 40572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1167_
timestamp 1688980957
transform 1 0 34684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1688980957
transform 1 0 42964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1688980957
transform 1 0 43516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1688980957
transform 1 0 40020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1171_
timestamp 1688980957
transform 1 0 35328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1172_
timestamp 1688980957
transform 1 0 36616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1688980957
transform 1 0 37260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1174_
timestamp 1688980957
transform 1 0 36064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1688980957
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1176_
timestamp 1688980957
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1177_
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1688980957
transform 1 0 26220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1179_
timestamp 1688980957
transform 1 0 25760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1688980957
transform 1 0 43884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1688980957
transform 1 0 44344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1688980957
transform 1 0 48944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1688980957
transform 1 0 47656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1688980957
transform 1 0 44160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1688980957
transform 1 0 48668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1186_
timestamp 1688980957
transform 1 0 42504 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1688980957
transform 1 0 51428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1688980957
transform 1 0 47196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1688980957
transform 1 0 51060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190_
timestamp 1688980957
transform 1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1191_
timestamp 1688980957
transform 1 0 41676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1192_
timestamp 1688980957
transform 1 0 41860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1688980957
transform 1 0 41492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1194_
timestamp 1688980957
transform 1 0 42044 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1195_
timestamp 1688980957
transform 1 0 40572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1196_
timestamp 1688980957
transform 1 0 35512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1197_
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198_
timestamp 1688980957
transform 1 0 36340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1199_
timestamp 1688980957
transform 1 0 34960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1688980957
transform 1 0 44436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1688980957
transform 1 0 47656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1688980957
transform 1 0 47012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1203_
timestamp 1688980957
transform 1 0 51336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1688980957
transform 1 0 51060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1205_
timestamp 1688980957
transform 1 0 43884 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1206_
timestamp 1688980957
transform 1 0 53452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1207_
timestamp 1688980957
transform 1 0 49772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1208_
timestamp 1688980957
transform 1 0 51244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp 1688980957
transform 1 0 52716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1688980957
transform 1 0 50048 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1211_
timestamp 1688980957
transform 1 0 46184 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1212_
timestamp 1688980957
transform 1 0 44988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1688980957
transform 1 0 41308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1688980957
transform 1 0 41032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1215_
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1216_
timestamp 1688980957
transform 1 0 41860 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1217_
timestamp 1688980957
transform 1 0 44436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1218_
timestamp 1688980957
transform 1 0 50508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1219_
timestamp 1688980957
transform 1 0 48944 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1220_
timestamp 1688980957
transform 1 0 50968 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1221_
timestamp 1688980957
transform 1 0 49588 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1222_
timestamp 1688980957
transform 1 0 49496 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1223_
timestamp 1688980957
transform 1 0 44988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1688980957
transform 1 0 44436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1688980957
transform 1 0 46644 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1226_
timestamp 1688980957
transform 1 0 43424 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1227_
timestamp 1688980957
transform 1 0 43240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1228_
timestamp 1688980957
transform 1 0 41032 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1229_
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1230_
timestamp 1688980957
transform 1 0 44160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1231_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1232_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30728 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp 1688980957
transform 1 0 27508 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 1688980957
transform 1 0 29716 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp 1688980957
transform 1 0 29440 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 1688980957
transform 1 0 27876 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp 1688980957
transform 1 0 35328 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1688980957
transform 1 0 34776 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1688980957
transform 1 0 35052 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1688980957
transform 1 0 37076 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 1688980957
transform 1 0 37812 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1688980957
transform 1 0 37444 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1688980957
transform 1 0 35236 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1688980957
transform 1 0 37168 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1688980957
transform 1 0 38824 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1688980957
transform 1 0 34040 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1688980957
transform 1 0 35420 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1688980957
transform 1 0 33948 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1688980957
transform 1 0 37352 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1688980957
transform 1 0 38548 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1688980957
transform 1 0 35328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 1688980957
transform 1 0 30728 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1688980957
transform 1 0 32200 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 1688980957
transform 1 0 33672 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1688980957
transform 1 0 46736 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1688980957
transform 1 0 45908 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1688980957
transform 1 0 42412 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1688980957
transform 1 0 40664 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1688980957
transform 1 0 40112 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1688980957
transform 1 0 39100 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1688980957
transform 1 0 39468 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1688980957
transform 1 0 29992 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1688980957
transform 1 0 31832 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1688980957
transform 1 0 32384 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1688980957
transform 1 0 30176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1688980957
transform 1 0 28152 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1688980957
transform 1 0 26036 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp 1688980957
transform 1 0 25576 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1688980957
transform 1 0 24932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1688980957
transform 1 0 25392 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1280_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 45448 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1281_
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1688980957
transform 1 0 44988 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1688980957
transform 1 0 41308 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1284_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1688980957
transform 1 0 33028 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1286_
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1688980957
transform 1 0 40848 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1289_
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1688980957
transform 1 0 42780 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1688980957
transform 1 0 27692 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1688980957
transform 1 0 28796 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1688980957
transform 1 0 31648 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1688980957
transform 1 0 34224 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1688980957
transform 1 0 32292 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1688980957
transform 1 0 35604 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1688980957
transform 1 0 35880 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1688980957
transform 1 0 32568 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1688980957
transform 1 0 29440 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1688980957
transform 1 0 31556 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1688980957
transform 1 0 33120 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1688980957
transform 1 0 32292 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1304_
timestamp 1688980957
transform 1 0 44436 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1305_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32200 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1306_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31004 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1307_
timestamp 1688980957
transform 1 0 31832 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1308_
timestamp 1688980957
transform 1 0 29348 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1309_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1310_
timestamp 1688980957
transform 1 0 25760 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1311_
timestamp 1688980957
transform 1 0 25392 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 1688980957
transform 1 0 25576 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 1688980957
transform 1 0 27600 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 1688980957
transform 1 0 30360 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1688980957
transform 1 0 30268 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1688980957
transform 1 0 28980 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1317_
timestamp 1688980957
transform 1 0 31096 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1318_
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1319_
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1320_
timestamp 1688980957
transform 1 0 22632 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1321_
timestamp 1688980957
transform 1 0 22356 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1322_
timestamp 1688980957
transform 1 0 22540 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1323_
timestamp 1688980957
transform 1 0 23184 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1324_
timestamp 1688980957
transform 1 0 25300 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1325_
timestamp 1688980957
transform 1 0 27600 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1326_
timestamp 1688980957
transform 1 0 28980 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1688980957
transform 1 0 27508 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1688980957
transform 1 0 27232 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1688980957
transform 1 0 29440 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1330_
timestamp 1688980957
transform 1 0 32752 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1331_
timestamp 1688980957
transform 1 0 37444 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1332_
timestamp 1688980957
transform 1 0 35052 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1333_
timestamp 1688980957
transform 1 0 34132 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1334_
timestamp 1688980957
transform 1 0 33856 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1335_
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1336_
timestamp 1688980957
transform 1 0 40020 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 1688980957
transform 1 0 39652 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1338_
timestamp 1688980957
transform 1 0 41124 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1339_
timestamp 1688980957
transform 1 0 41676 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1340_
timestamp 1688980957
transform 1 0 38180 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1688980957
transform 1 0 36340 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1343_
timestamp 1688980957
transform 1 0 32752 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1688980957
transform 1 0 25208 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1688980957
transform 1 0 23736 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1688980957
transform 1 0 38824 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1688980957
transform 1 0 38824 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1688980957
transform 1 0 40204 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1350_
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1351_
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1352_
timestamp 1688980957
transform 1 0 42964 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1353_
timestamp 1688980957
transform 1 0 43424 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1354_
timestamp 1688980957
transform 1 0 47104 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1355_
timestamp 1688980957
transform 1 0 45540 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1356_
timestamp 1688980957
transform 1 0 42964 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1357_
timestamp 1688980957
transform 1 0 48024 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1358_
timestamp 1688980957
transform 1 0 49496 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1359_
timestamp 1688980957
transform 1 0 46368 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1360_
timestamp 1688980957
transform 1 0 49220 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1361_
timestamp 1688980957
transform 1 0 43056 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1688980957
transform 1 0 41768 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1688980957
transform 1 0 41768 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1364_
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1688980957
transform 1 0 34408 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1688980957
transform 1 0 34868 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1367_
timestamp 1688980957
transform 1 0 42964 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1368_
timestamp 1688980957
transform 1 0 47564 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1369_
timestamp 1688980957
transform 1 0 46184 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1370_
timestamp 1688980957
transform 1 0 50508 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1371_
timestamp 1688980957
transform 1 0 49220 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1372_
timestamp 1688980957
transform 1 0 51980 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1373_
timestamp 1688980957
transform 1 0 48852 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1374_
timestamp 1688980957
transform 1 0 50140 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1375_
timestamp 1688980957
transform 1 0 52716 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1376_
timestamp 1688980957
transform 1 0 48208 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1688980957
transform 1 0 46736 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1378_
timestamp 1688980957
transform 1 0 43056 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1688980957
transform 1 0 40848 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1381_
timestamp 1688980957
transform 1 0 42964 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1382_
timestamp 1688980957
transform 1 0 49680 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1383_
timestamp 1688980957
transform 1 0 47564 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1384_
timestamp 1688980957
transform 1 0 50140 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1385_
timestamp 1688980957
transform 1 0 49036 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1386_
timestamp 1688980957
transform 1 0 47656 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1387_
timestamp 1688980957
transform 1 0 44068 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1388_
timestamp 1688980957
transform 1 0 43608 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1389_
timestamp 1688980957
transform 1 0 45540 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1390_
timestamp 1688980957
transform 1 0 42504 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1688980957
transform 1 0 40756 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1688980957
transform 1 0 42412 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1688980957
transform 1 0 45080 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 67712 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37444 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform 1 0 27508 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform 1 0 33120 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 33580 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform 1 0 28428 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform 1 0 28428 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform 1 0 34040 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform 1 0 40848 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 40756 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform 1 0 46368 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 47012 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 41308 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform 1 0 41308 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform 1 0 47656 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 47380 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_7 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_8
timestamp 1688980957
transform 1 0 20056 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_9
timestamp 1688980957
transform 1 0 22632 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_10
timestamp 1688980957
transform 1 0 58696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_11
timestamp 1688980957
transform 1 0 27784 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_12
timestamp 1688980957
transform 1 0 68264 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_13
timestamp 1688980957
transform 1 0 68264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_14
timestamp 1688980957
transform 1 0 32936 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_15
timestamp 1688980957
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_16
timestamp 1688980957
transform 1 0 68264 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_17
timestamp 1688980957
transform 1 0 68264 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_18
timestamp 1688980957
transform 1 0 68264 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_19
timestamp 1688980957
transform 1 0 58696 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_20
timestamp 1688980957
transform 1 0 68264 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_21
timestamp 1688980957
transform 1 0 68264 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_22
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_23
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_24
timestamp 1688980957
transform 1 0 68264 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_25
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_26
timestamp 1688980957
transform 1 0 1380 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_27
timestamp 1688980957
transform 1 0 38088 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_28
timestamp 1688980957
transform 1 0 63848 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_29
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_30
timestamp 1688980957
transform 1 0 68264 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_31
timestamp 1688980957
transform 1 0 1380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_32
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_33
timestamp 1688980957
transform 1 0 68264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_34
timestamp 1688980957
transform 1 0 53544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_35
timestamp 1688980957
transform 1 0 68264 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_36
timestamp 1688980957
transform 1 0 68264 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_37
timestamp 1688980957
transform 1 0 25208 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_38
timestamp 1688980957
transform 1 0 68264 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_39
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_40
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_41
timestamp 1688980957
transform 1 0 68264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_42
timestamp 1688980957
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_43
timestamp 1688980957
transform 1 0 68264 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_44
timestamp 1688980957
transform 1 0 1380 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_45
timestamp 1688980957
transform 1 0 68264 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_46
timestamp 1688980957
transform 1 0 68264 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_47
timestamp 1688980957
transform 1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_48
timestamp 1688980957
transform 1 0 61272 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_49
timestamp 1688980957
transform 1 0 45816 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_50
timestamp 1688980957
transform 1 0 30544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_51
timestamp 1688980957
transform 1 0 68264 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_52
timestamp 1688980957
transform 1 0 68264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_53
timestamp 1688980957
transform 1 0 2024 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_54
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_55
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_56
timestamp 1688980957
transform 1 0 40664 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_57
timestamp 1688980957
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_58
timestamp 1688980957
transform 1 0 17480 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_59
timestamp 1688980957
transform 1 0 1380 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_60
timestamp 1688980957
transform 1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_61
timestamp 1688980957
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_62
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_63
timestamp 1688980957
transform 1 0 66424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_64
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_65
timestamp 1688980957
transform 1 0 50968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_66
timestamp 1688980957
transform 1 0 1380 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_67
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_68
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_69
timestamp 1688980957
transform 1 0 68264 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_70
timestamp 1688980957
transform 1 0 68264 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_71
timestamp 1688980957
transform 1 0 56120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_72
timestamp 1688980957
transform 1 0 68264 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_73
timestamp 1688980957
transform 1 0 7176 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_74
timestamp 1688980957
transform 1 0 9752 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_75
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_76
timestamp 1688980957
transform 1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_77
timestamp 1688980957
transform 1 0 12328 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_78
timestamp 1688980957
transform 1 0 30360 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_79
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_80
timestamp 1688980957
transform 1 0 1380 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_81
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_82
timestamp 1688980957
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_83
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_84
timestamp 1688980957
transform 1 0 68264 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_85
timestamp 1688980957
transform 1 0 38456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_86
timestamp 1688980957
transform 1 0 53544 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_87
timestamp 1688980957
transform 1 0 4600 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_88
timestamp 1688980957
transform 1 0 14904 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_89
timestamp 1688980957
transform 1 0 56120 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_128
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_261
timestamp 1688980957
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_293 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_300
timestamp 1688980957
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_323
timestamp 1688980957
transform 1 0 30820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_373 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_384
timestamp 1688980957
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_401
timestamp 1688980957
transform 1 0 37996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_409
timestamp 1688980957
transform 1 0 38732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_432
timestamp 1688980957
transform 1 0 40848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_444
timestamp 1688980957
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_457
timestamp 1688980957
transform 1 0 43148 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 1688980957
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_477
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_485
timestamp 1688980957
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_489
timestamp 1688980957
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 1688980957
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_505
timestamp 1688980957
transform 1 0 47564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_513
timestamp 1688980957
transform 1 0 48300 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_520
timestamp 1688980957
transform 1 0 48944 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_533
timestamp 1688980957
transform 1 0 50140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_541
timestamp 1688980957
transform 1 0 50876 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_545
timestamp 1688980957
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 1688980957
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_561
timestamp 1688980957
transform 1 0 52716 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_569
timestamp 1688980957
transform 1 0 53452 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_573
timestamp 1688980957
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 1688980957
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_589
timestamp 1688980957
transform 1 0 55292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_597
timestamp 1688980957
transform 1 0 56028 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_601
timestamp 1688980957
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 1688980957
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_617
timestamp 1688980957
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_625
timestamp 1688980957
transform 1 0 58604 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_629
timestamp 1688980957
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_641
timestamp 1688980957
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_645
timestamp 1688980957
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_657
timestamp 1688980957
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_669
timestamp 1688980957
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_673
timestamp 1688980957
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_685
timestamp 1688980957
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_697
timestamp 1688980957
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_701
timestamp 1688980957
transform 1 0 65596 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_709
timestamp 1688980957
transform 1 0 66332 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_713
timestamp 1688980957
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_729
timestamp 1688980957
transform 1 0 68172 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_285
timestamp 1688980957
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_340
timestamp 1688980957
transform 1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_346
timestamp 1688980957
transform 1 0 32936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_358
timestamp 1688980957
transform 1 0 34040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_366
timestamp 1688980957
transform 1 0 34776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_416
timestamp 1688980957
transform 1 0 39376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_439
timestamp 1688980957
transform 1 0 41492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_485
timestamp 1688980957
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_497
timestamp 1688980957
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 1688980957
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_508
timestamp 1688980957
transform 1 0 47840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_520
timestamp 1688980957
transform 1 0 48944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_532
timestamp 1688980957
transform 1 0 50048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_544
timestamp 1688980957
transform 1 0 51152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_556
timestamp 1688980957
transform 1 0 52256 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_561
timestamp 1688980957
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_573
timestamp 1688980957
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_585
timestamp 1688980957
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_597
timestamp 1688980957
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_609
timestamp 1688980957
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_615
timestamp 1688980957
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_617
timestamp 1688980957
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_629
timestamp 1688980957
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_641
timestamp 1688980957
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_653
timestamp 1688980957
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_665
timestamp 1688980957
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_671
timestamp 1688980957
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_673
timestamp 1688980957
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_685
timestamp 1688980957
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_697
timestamp 1688980957
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_709
timestamp 1688980957
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_721
timestamp 1688980957
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_727
timestamp 1688980957
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_729
timestamp 1688980957
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_306
timestamp 1688980957
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_313
timestamp 1688980957
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_348
timestamp 1688980957
transform 1 0 33120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_360
timestamp 1688980957
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_368
timestamp 1688980957
transform 1 0 34960 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_376
timestamp 1688980957
transform 1 0 35696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_387
timestamp 1688980957
transform 1 0 36708 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_395
timestamp 1688980957
transform 1 0 37444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_411
timestamp 1688980957
transform 1 0 38916 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_444
timestamp 1688980957
transform 1 0 41952 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_456
timestamp 1688980957
transform 1 0 43056 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_468
timestamp 1688980957
transform 1 0 44160 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 1688980957
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 1688980957
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 1688980957
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 1688980957
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 1688980957
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1688980957
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1688980957
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 1688980957
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_569
timestamp 1688980957
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_581
timestamp 1688980957
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 1688980957
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_589
timestamp 1688980957
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_601
timestamp 1688980957
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_613
timestamp 1688980957
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_625
timestamp 1688980957
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_637
timestamp 1688980957
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_643
timestamp 1688980957
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_645
timestamp 1688980957
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_657
timestamp 1688980957
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_669
timestamp 1688980957
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_681
timestamp 1688980957
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_693
timestamp 1688980957
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_699
timestamp 1688980957
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_701
timestamp 1688980957
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_713
timestamp 1688980957
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_725
timestamp 1688980957
transform 1 0 67804 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_729
timestamp 1688980957
transform 1 0 68172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_284
timestamp 1688980957
transform 1 0 27232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_296
timestamp 1688980957
transform 1 0 28336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_302
timestamp 1688980957
transform 1 0 28888 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_310
timestamp 1688980957
transform 1 0 29624 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_320
timestamp 1688980957
transform 1 0 30544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_330
timestamp 1688980957
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_345
timestamp 1688980957
transform 1 0 32844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_355
timestamp 1688980957
transform 1 0 33764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_377
timestamp 1688980957
transform 1 0 35788 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_386
timestamp 1688980957
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_404
timestamp 1688980957
transform 1 0 38272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_419
timestamp 1688980957
transform 1 0 39652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_437
timestamp 1688980957
transform 1 0 41308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_445
timestamp 1688980957
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 1688980957
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 1688980957
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 1688980957
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_505
timestamp 1688980957
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_517
timestamp 1688980957
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 1688980957
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 1688980957
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 1688980957
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 1688980957
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 1688980957
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 1688980957
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 1688980957
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_597
timestamp 1688980957
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_609
timestamp 1688980957
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1688980957
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_617
timestamp 1688980957
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_629
timestamp 1688980957
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_641
timestamp 1688980957
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_653
timestamp 1688980957
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_665
timestamp 1688980957
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_671
timestamp 1688980957
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_673
timestamp 1688980957
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_685
timestamp 1688980957
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_697
timestamp 1688980957
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_709
timestamp 1688980957
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_721
timestamp 1688980957
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_727
timestamp 1688980957
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_729
timestamp 1688980957
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_297
timestamp 1688980957
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_305
timestamp 1688980957
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_317
timestamp 1688980957
transform 1 0 30268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_326
timestamp 1688980957
transform 1 0 31096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_354
timestamp 1688980957
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_362
timestamp 1688980957
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_371
timestamp 1688980957
transform 1 0 35236 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_404
timestamp 1688980957
transform 1 0 38272 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_412
timestamp 1688980957
transform 1 0 39008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_428
timestamp 1688980957
transform 1 0 40480 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_434
timestamp 1688980957
transform 1 0 41032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_458
timestamp 1688980957
transform 1 0 43240 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_473
timestamp 1688980957
transform 1 0 44620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_509
timestamp 1688980957
transform 1 0 47932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_521
timestamp 1688980957
transform 1 0 49036 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_529
timestamp 1688980957
transform 1 0 49772 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 1688980957
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 1688980957
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 1688980957
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 1688980957
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 1688980957
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 1688980957
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1688980957
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1688980957
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1688980957
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_625
timestamp 1688980957
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_637
timestamp 1688980957
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_643
timestamp 1688980957
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_645
timestamp 1688980957
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_657
timestamp 1688980957
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_669
timestamp 1688980957
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_681
timestamp 1688980957
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_693
timestamp 1688980957
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_699
timestamp 1688980957
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_701
timestamp 1688980957
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_713
timestamp 1688980957
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_725
timestamp 1688980957
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_269
timestamp 1688980957
transform 1 0 25852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1688980957
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_310
timestamp 1688980957
transform 1 0 29624 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_318
timestamp 1688980957
transform 1 0 30360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_324
timestamp 1688980957
transform 1 0 30912 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_330
timestamp 1688980957
transform 1 0 31464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_348
timestamp 1688980957
transform 1 0 33120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_357
timestamp 1688980957
transform 1 0 33948 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_387
timestamp 1688980957
transform 1 0 36708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_413
timestamp 1688980957
transform 1 0 39100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_421
timestamp 1688980957
transform 1 0 39836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_427
timestamp 1688980957
transform 1 0 40388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_440
timestamp 1688980957
transform 1 0 41584 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_457
timestamp 1688980957
transform 1 0 43148 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_502
timestamp 1688980957
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_516
timestamp 1688980957
transform 1 0 48576 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_528
timestamp 1688980957
transform 1 0 49680 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_540
timestamp 1688980957
transform 1 0 50784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_552
timestamp 1688980957
transform 1 0 51888 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 1688980957
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 1688980957
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 1688980957
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 1688980957
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 1688980957
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 1688980957
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_617
timestamp 1688980957
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_629
timestamp 1688980957
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_641
timestamp 1688980957
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_653
timestamp 1688980957
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_665
timestamp 1688980957
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_671
timestamp 1688980957
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_673
timestamp 1688980957
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_685
timestamp 1688980957
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_697
timestamp 1688980957
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_709
timestamp 1688980957
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_721
timestamp 1688980957
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_727
timestamp 1688980957
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_729
timestamp 1688980957
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_261
timestamp 1688980957
transform 1 0 25116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_299
timestamp 1688980957
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_315
timestamp 1688980957
transform 1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_336
timestamp 1688980957
transform 1 0 32016 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_356
timestamp 1688980957
transform 1 0 33856 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_386
timestamp 1688980957
transform 1 0 36616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_395
timestamp 1688980957
transform 1 0 37444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_405
timestamp 1688980957
transform 1 0 38364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_434
timestamp 1688980957
transform 1 0 41032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_440
timestamp 1688980957
transform 1 0 41584 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_464
timestamp 1688980957
transform 1 0 43792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_490
timestamp 1688980957
transform 1 0 46184 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_498
timestamp 1688980957
transform 1 0 46920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_523
timestamp 1688980957
transform 1 0 49220 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 1688980957
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1688980957
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 1688980957
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 1688980957
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 1688980957
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 1688980957
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 1688980957
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1688980957
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1688980957
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1688980957
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_625
timestamp 1688980957
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_637
timestamp 1688980957
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_643
timestamp 1688980957
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_645
timestamp 1688980957
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_657
timestamp 1688980957
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_669
timestamp 1688980957
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_681
timestamp 1688980957
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_693
timestamp 1688980957
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_699
timestamp 1688980957
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_701
timestamp 1688980957
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_713
timestamp 1688980957
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_725
timestamp 1688980957
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_322
timestamp 1688980957
transform 1 0 30728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_327
timestamp 1688980957
transform 1 0 31188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_334
timestamp 1688980957
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_343
timestamp 1688980957
transform 1 0 32660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_365
timestamp 1688980957
transform 1 0 34684 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_381
timestamp 1688980957
transform 1 0 36156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_400
timestamp 1688980957
transform 1 0 37904 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_415
timestamp 1688980957
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_430
timestamp 1688980957
transform 1 0 40664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_440
timestamp 1688980957
transform 1 0 41584 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_467
timestamp 1688980957
transform 1 0 44068 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_471
timestamp 1688980957
transform 1 0 44436 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_501
timestamp 1688980957
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_505
timestamp 1688980957
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_520
timestamp 1688980957
transform 1 0 48944 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_532
timestamp 1688980957
transform 1 0 50048 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_544
timestamp 1688980957
transform 1 0 51152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_556
timestamp 1688980957
transform 1 0 52256 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_561
timestamp 1688980957
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_573
timestamp 1688980957
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_585
timestamp 1688980957
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_597
timestamp 1688980957
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 1688980957
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 1688980957
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_617
timestamp 1688980957
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_629
timestamp 1688980957
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_641
timestamp 1688980957
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_653
timestamp 1688980957
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_665
timestamp 1688980957
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_671
timestamp 1688980957
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_673
timestamp 1688980957
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_685
timestamp 1688980957
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_697
timestamp 1688980957
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_709
timestamp 1688980957
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_721
timestamp 1688980957
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_727
timestamp 1688980957
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_729
timestamp 1688980957
transform 1 0 68172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_290
timestamp 1688980957
transform 1 0 27784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_306
timestamp 1688980957
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_316
timestamp 1688980957
transform 1 0 30176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_328
timestamp 1688980957
transform 1 0 31280 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_337
timestamp 1688980957
transform 1 0 32108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_349
timestamp 1688980957
transform 1 0 33212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_358
timestamp 1688980957
transform 1 0 34040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_374
timestamp 1688980957
transform 1 0 35512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_382
timestamp 1688980957
transform 1 0 36248 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_386
timestamp 1688980957
transform 1 0 36616 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_392
timestamp 1688980957
transform 1 0 37168 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_399
timestamp 1688980957
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_403
timestamp 1688980957
transform 1 0 38180 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_412
timestamp 1688980957
transform 1 0 39008 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_430
timestamp 1688980957
transform 1 0 40664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_442
timestamp 1688980957
transform 1 0 41768 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_447
timestamp 1688980957
transform 1 0 42228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_500
timestamp 1688980957
transform 1 0 47104 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_508
timestamp 1688980957
transform 1 0 47840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_530
timestamp 1688980957
transform 1 0 49864 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_533
timestamp 1688980957
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_545
timestamp 1688980957
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_557
timestamp 1688980957
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 1688980957
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 1688980957
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 1688980957
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 1688980957
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 1688980957
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 1688980957
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_625
timestamp 1688980957
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_637
timestamp 1688980957
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_643
timestamp 1688980957
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_645
timestamp 1688980957
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_657
timestamp 1688980957
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_669
timestamp 1688980957
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_681
timestamp 1688980957
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_693
timestamp 1688980957
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_699
timestamp 1688980957
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_701
timestamp 1688980957
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_713
timestamp 1688980957
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_725
timestamp 1688980957
transform 1 0 67804 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_276
timestamp 1688980957
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_324
timestamp 1688980957
transform 1 0 30912 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_346
timestamp 1688980957
transform 1 0 32936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_356
timestamp 1688980957
transform 1 0 33856 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_364
timestamp 1688980957
transform 1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_401
timestamp 1688980957
transform 1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_426
timestamp 1688980957
transform 1 0 40296 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_465
timestamp 1688980957
transform 1 0 43884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_469
timestamp 1688980957
transform 1 0 44252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_479
timestamp 1688980957
transform 1 0 45172 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_498
timestamp 1688980957
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_505
timestamp 1688980957
transform 1 0 47564 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_530
timestamp 1688980957
transform 1 0 49864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_542
timestamp 1688980957
transform 1 0 50968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_554
timestamp 1688980957
transform 1 0 52072 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_561
timestamp 1688980957
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 1688980957
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 1688980957
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 1688980957
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 1688980957
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 1688980957
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_617
timestamp 1688980957
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_629
timestamp 1688980957
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_641
timestamp 1688980957
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_653
timestamp 1688980957
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_665
timestamp 1688980957
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_671
timestamp 1688980957
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_673
timestamp 1688980957
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_685
timestamp 1688980957
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_697
timestamp 1688980957
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_709
timestamp 1688980957
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_721
timestamp 1688980957
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_727
timestamp 1688980957
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_729
timestamp 1688980957
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 1688980957
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 1688980957
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1688980957
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_256
timestamp 1688980957
transform 1 0 24656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_262
timestamp 1688980957
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_283
timestamp 1688980957
transform 1 0 27140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_287
timestamp 1688980957
transform 1 0 27508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_313
timestamp 1688980957
transform 1 0 29900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_317
timestamp 1688980957
transform 1 0 30268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_359
timestamp 1688980957
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_380
timestamp 1688980957
transform 1 0 36064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_468
timestamp 1688980957
transform 1 0 44160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_485
timestamp 1688980957
transform 1 0 45724 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_499
timestamp 1688980957
transform 1 0 47012 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_503
timestamp 1688980957
transform 1 0 47380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_517
timestamp 1688980957
transform 1 0 48668 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_530
timestamp 1688980957
transform 1 0 49864 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 1688980957
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 1688980957
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 1688980957
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 1688980957
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 1688980957
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 1688980957
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 1688980957
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 1688980957
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_613
timestamp 1688980957
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_625
timestamp 1688980957
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_637
timestamp 1688980957
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_643
timestamp 1688980957
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_645
timestamp 1688980957
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_657
timestamp 1688980957
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_669
timestamp 1688980957
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_681
timestamp 1688980957
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_693
timestamp 1688980957
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_699
timestamp 1688980957
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_701
timestamp 1688980957
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_713
timestamp 1688980957
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_725
timestamp 1688980957
transform 1 0 67804 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_260
timestamp 1688980957
transform 1 0 25024 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_272
timestamp 1688980957
transform 1 0 26128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_294
timestamp 1688980957
transform 1 0 28152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_306
timestamp 1688980957
transform 1 0 29256 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_318
timestamp 1688980957
transform 1 0 30360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_322
timestamp 1688980957
transform 1 0 30728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_326
timestamp 1688980957
transform 1 0 31096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 1688980957
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_346
timestamp 1688980957
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_352
timestamp 1688980957
transform 1 0 33488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_359
timestamp 1688980957
transform 1 0 34132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_389
timestamp 1688980957
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_402
timestamp 1688980957
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_408
timestamp 1688980957
transform 1 0 38640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_420
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_428
timestamp 1688980957
transform 1 0 40480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_446
timestamp 1688980957
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_455
timestamp 1688980957
transform 1 0 42964 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_479
timestamp 1688980957
transform 1 0 45172 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_485
timestamp 1688980957
transform 1 0 45724 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 1688980957
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_505
timestamp 1688980957
transform 1 0 47564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_511
timestamp 1688980957
transform 1 0 48116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_520
timestamp 1688980957
transform 1 0 48944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_550
timestamp 1688980957
transform 1 0 51704 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_558
timestamp 1688980957
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 1688980957
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 1688980957
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 1688980957
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 1688980957
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 1688980957
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1688980957
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_617
timestamp 1688980957
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_629
timestamp 1688980957
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_641
timestamp 1688980957
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_653
timestamp 1688980957
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_665
timestamp 1688980957
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_671
timestamp 1688980957
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_673
timestamp 1688980957
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_685
timestamp 1688980957
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_697
timestamp 1688980957
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_709
timestamp 1688980957
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_721
timestamp 1688980957
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_727
timestamp 1688980957
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_729
timestamp 1688980957
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_241
timestamp 1688980957
transform 1 0 23276 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_247
timestamp 1688980957
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_257
timestamp 1688980957
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_266
timestamp 1688980957
transform 1 0 25576 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_312
timestamp 1688980957
transform 1 0 29808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_316
timestamp 1688980957
transform 1 0 30176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_359
timestamp 1688980957
transform 1 0 34132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_371
timestamp 1688980957
transform 1 0 35236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_388
timestamp 1688980957
transform 1 0 36800 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_394
timestamp 1688980957
transform 1 0 37352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_416
timestamp 1688980957
transform 1 0 39376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_489
timestamp 1688980957
transform 1 0 46092 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_512
timestamp 1688980957
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 1688980957
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 1688980957
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 1688980957
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 1688980957
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 1688980957
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 1688980957
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 1688980957
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 1688980957
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 1688980957
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 1688980957
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_625
timestamp 1688980957
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_637
timestamp 1688980957
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_643
timestamp 1688980957
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_645
timestamp 1688980957
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_657
timestamp 1688980957
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_669
timestamp 1688980957
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_681
timestamp 1688980957
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_693
timestamp 1688980957
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_699
timestamp 1688980957
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_701
timestamp 1688980957
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_713
timestamp 1688980957
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_725
timestamp 1688980957
transform 1 0 67804 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_729
timestamp 1688980957
transform 1 0 68172 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_275
timestamp 1688980957
transform 1 0 26404 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_287
timestamp 1688980957
transform 1 0 27508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_292
timestamp 1688980957
transform 1 0 27968 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_300
timestamp 1688980957
transform 1 0 28704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_340
timestamp 1688980957
transform 1 0 32384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_371
timestamp 1688980957
transform 1 0 35236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_378
timestamp 1688980957
transform 1 0 35880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_388
timestamp 1688980957
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_407
timestamp 1688980957
transform 1 0 38548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_423
timestamp 1688980957
transform 1 0 40020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_445
timestamp 1688980957
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_457
timestamp 1688980957
transform 1 0 43148 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_461
timestamp 1688980957
transform 1 0 43516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_481
timestamp 1688980957
transform 1 0 45356 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_485
timestamp 1688980957
transform 1 0 45724 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_490
timestamp 1688980957
transform 1 0 46184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_497
timestamp 1688980957
transform 1 0 46828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_505
timestamp 1688980957
transform 1 0 47564 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_522
timestamp 1688980957
transform 1 0 49128 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_546
timestamp 1688980957
transform 1 0 51336 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_558
timestamp 1688980957
transform 1 0 52440 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_561
timestamp 1688980957
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_573
timestamp 1688980957
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_585
timestamp 1688980957
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_597
timestamp 1688980957
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_609
timestamp 1688980957
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 1688980957
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_617
timestamp 1688980957
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_629
timestamp 1688980957
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_641
timestamp 1688980957
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_653
timestamp 1688980957
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_665
timestamp 1688980957
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_671
timestamp 1688980957
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_673
timestamp 1688980957
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_685
timestamp 1688980957
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_697
timestamp 1688980957
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_709
timestamp 1688980957
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_721
timestamp 1688980957
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_727
timestamp 1688980957
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_729
timestamp 1688980957
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_263
timestamp 1688980957
transform 1 0 25300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_273
timestamp 1688980957
transform 1 0 26220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_317
timestamp 1688980957
transform 1 0 30268 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_374
timestamp 1688980957
transform 1 0 35512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_396
timestamp 1688980957
transform 1 0 37536 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_417
timestamp 1688980957
transform 1 0 39468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_421
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_436
timestamp 1688980957
transform 1 0 41216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_453
timestamp 1688980957
transform 1 0 42780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_492
timestamp 1688980957
transform 1 0 46368 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_498
timestamp 1688980957
transform 1 0 46920 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_515
timestamp 1688980957
transform 1 0 48484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_527
timestamp 1688980957
transform 1 0 49588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 1688980957
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_541
timestamp 1688980957
transform 1 0 50876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_553
timestamp 1688980957
transform 1 0 51980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_565
timestamp 1688980957
transform 1 0 53084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_577
timestamp 1688980957
transform 1 0 54188 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_585
timestamp 1688980957
transform 1 0 54924 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_589
timestamp 1688980957
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_601
timestamp 1688980957
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_613
timestamp 1688980957
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_625
timestamp 1688980957
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_637
timestamp 1688980957
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_643
timestamp 1688980957
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_645
timestamp 1688980957
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_657
timestamp 1688980957
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_669
timestamp 1688980957
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_681
timestamp 1688980957
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_693
timestamp 1688980957
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_699
timestamp 1688980957
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_701
timestamp 1688980957
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_713
timestamp 1688980957
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_725
timestamp 1688980957
transform 1 0 67804 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_6
timestamp 1688980957
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_18
timestamp 1688980957
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_30
timestamp 1688980957
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_42
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1688980957
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_246
timestamp 1688980957
transform 1 0 23736 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_252
timestamp 1688980957
transform 1 0 24288 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_271
timestamp 1688980957
transform 1 0 26036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_298
timestamp 1688980957
transform 1 0 28520 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_312
timestamp 1688980957
transform 1 0 29808 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_324
timestamp 1688980957
transform 1 0 30912 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_362
timestamp 1688980957
transform 1 0 34408 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_370
timestamp 1688980957
transform 1 0 35144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_401
timestamp 1688980957
transform 1 0 37996 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_413
timestamp 1688980957
transform 1 0 39100 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_421
timestamp 1688980957
transform 1 0 39836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_447
timestamp 1688980957
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_457
timestamp 1688980957
transform 1 0 43148 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_463
timestamp 1688980957
transform 1 0 43700 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_482
timestamp 1688980957
transform 1 0 45448 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_494
timestamp 1688980957
transform 1 0 46552 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_502
timestamp 1688980957
transform 1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_505
timestamp 1688980957
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_517
timestamp 1688980957
transform 1 0 48668 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_549
timestamp 1688980957
transform 1 0 51612 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_557
timestamp 1688980957
transform 1 0 52348 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_561
timestamp 1688980957
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_573
timestamp 1688980957
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_585
timestamp 1688980957
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_597
timestamp 1688980957
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_609
timestamp 1688980957
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_615
timestamp 1688980957
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_617
timestamp 1688980957
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_629
timestamp 1688980957
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_641
timestamp 1688980957
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_653
timestamp 1688980957
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_665
timestamp 1688980957
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_671
timestamp 1688980957
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_673
timestamp 1688980957
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_685
timestamp 1688980957
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_697
timestamp 1688980957
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_709
timestamp 1688980957
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_721
timestamp 1688980957
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_727
timestamp 1688980957
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_729
timestamp 1688980957
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_229
timestamp 1688980957
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_279
timestamp 1688980957
transform 1 0 26772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_327
timestamp 1688980957
transform 1 0 31188 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_347
timestamp 1688980957
transform 1 0 33028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_359
timestamp 1688980957
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_410
timestamp 1688980957
transform 1 0 38824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_417
timestamp 1688980957
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_437
timestamp 1688980957
transform 1 0 41308 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_458
timestamp 1688980957
transform 1 0 43240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_470
timestamp 1688980957
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_477
timestamp 1688980957
transform 1 0 44988 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_485
timestamp 1688980957
transform 1 0 45724 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_495
timestamp 1688980957
transform 1 0 46644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_501
timestamp 1688980957
transform 1 0 47196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_505
timestamp 1688980957
transform 1 0 47564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_518
timestamp 1688980957
transform 1 0 48760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_531
timestamp 1688980957
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_533
timestamp 1688980957
transform 1 0 50140 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_560
timestamp 1688980957
transform 1 0 52624 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_572
timestamp 1688980957
transform 1 0 53728 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_584
timestamp 1688980957
transform 1 0 54832 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_589
timestamp 1688980957
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_601
timestamp 1688980957
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_613
timestamp 1688980957
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_625
timestamp 1688980957
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_637
timestamp 1688980957
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_643
timestamp 1688980957
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_645
timestamp 1688980957
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_657
timestamp 1688980957
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_669
timestamp 1688980957
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_681
timestamp 1688980957
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_693
timestamp 1688980957
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_699
timestamp 1688980957
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_701
timestamp 1688980957
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_713
timestamp 1688980957
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_725
timestamp 1688980957
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_260
timestamp 1688980957
transform 1 0 25024 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_268
timestamp 1688980957
transform 1 0 25760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 1688980957
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_286
timestamp 1688980957
transform 1 0 27416 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_292
timestamp 1688980957
transform 1 0 27968 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_297
timestamp 1688980957
transform 1 0 28428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_334
timestamp 1688980957
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_363
timestamp 1688980957
transform 1 0 34500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_372
timestamp 1688980957
transform 1 0 35328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_409
timestamp 1688980957
transform 1 0 38732 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 1688980957
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_457
timestamp 1688980957
transform 1 0 43148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_465
timestamp 1688980957
transform 1 0 43884 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_482
timestamp 1688980957
transform 1 0 45448 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_494
timestamp 1688980957
transform 1 0 46552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_498
timestamp 1688980957
transform 1 0 46920 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_502
timestamp 1688980957
transform 1 0 47288 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_534
timestamp 1688980957
transform 1 0 50232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_558
timestamp 1688980957
transform 1 0 52440 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_564
timestamp 1688980957
transform 1 0 52992 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_576
timestamp 1688980957
transform 1 0 54096 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_588
timestamp 1688980957
transform 1 0 55200 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_600
timestamp 1688980957
transform 1 0 56304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_612
timestamp 1688980957
transform 1 0 57408 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_617
timestamp 1688980957
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_629
timestamp 1688980957
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_641
timestamp 1688980957
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_653
timestamp 1688980957
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_665
timestamp 1688980957
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_671
timestamp 1688980957
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_673
timestamp 1688980957
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_685
timestamp 1688980957
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_697
timestamp 1688980957
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_709
timestamp 1688980957
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_721
timestamp 1688980957
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_727
timestamp 1688980957
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_729
timestamp 1688980957
transform 1 0 68172 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_241
timestamp 1688980957
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_247
timestamp 1688980957
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_262
timestamp 1688980957
transform 1 0 25208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_274
timestamp 1688980957
transform 1 0 26312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_279
timestamp 1688980957
transform 1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_287
timestamp 1688980957
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_299
timestamp 1688980957
transform 1 0 28612 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_350
timestamp 1688980957
transform 1 0 33304 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_356
timestamp 1688980957
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_381
timestamp 1688980957
transform 1 0 36156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_415
timestamp 1688980957
transform 1 0 39284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 1688980957
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_425
timestamp 1688980957
transform 1 0 40204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_449
timestamp 1688980957
transform 1 0 42412 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_480
timestamp 1688980957
transform 1 0 45264 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_488
timestamp 1688980957
transform 1 0 46000 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_511
timestamp 1688980957
transform 1 0 48116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_523
timestamp 1688980957
transform 1 0 49220 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_531
timestamp 1688980957
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_540
timestamp 1688980957
transform 1 0 50784 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_551
timestamp 1688980957
transform 1 0 51796 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_563
timestamp 1688980957
transform 1 0 52900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_575
timestamp 1688980957
transform 1 0 54004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_587
timestamp 1688980957
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_589
timestamp 1688980957
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_601
timestamp 1688980957
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_613
timestamp 1688980957
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_625
timestamp 1688980957
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_637
timestamp 1688980957
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_643
timestamp 1688980957
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_645
timestamp 1688980957
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_657
timestamp 1688980957
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_669
timestamp 1688980957
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_681
timestamp 1688980957
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_693
timestamp 1688980957
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_699
timestamp 1688980957
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_701
timestamp 1688980957
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_713
timestamp 1688980957
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_725
timestamp 1688980957
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_233
timestamp 1688980957
transform 1 0 22540 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_350
timestamp 1688980957
transform 1 0 33304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_367
timestamp 1688980957
transform 1 0 34868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_403
timestamp 1688980957
transform 1 0 38180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_414
timestamp 1688980957
transform 1 0 39192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_418
timestamp 1688980957
transform 1 0 39560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_435
timestamp 1688980957
transform 1 0 41124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_439
timestamp 1688980957
transform 1 0 41492 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 1688980957
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_474
timestamp 1688980957
transform 1 0 44712 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_482
timestamp 1688980957
transform 1 0 45448 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_489
timestamp 1688980957
transform 1 0 46092 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_501
timestamp 1688980957
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_505
timestamp 1688980957
transform 1 0 47564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_519
timestamp 1688980957
transform 1 0 48852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_537
timestamp 1688980957
transform 1 0 50508 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_543
timestamp 1688980957
transform 1 0 51060 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_557
timestamp 1688980957
transform 1 0 52348 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_572
timestamp 1688980957
transform 1 0 53728 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_584
timestamp 1688980957
transform 1 0 54832 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_596
timestamp 1688980957
transform 1 0 55936 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_608
timestamp 1688980957
transform 1 0 57040 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_617
timestamp 1688980957
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_629
timestamp 1688980957
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_641
timestamp 1688980957
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_653
timestamp 1688980957
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_665
timestamp 1688980957
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_671
timestamp 1688980957
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_673
timestamp 1688980957
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_685
timestamp 1688980957
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_697
timestamp 1688980957
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_709
timestamp 1688980957
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_721
timestamp 1688980957
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_727
timestamp 1688980957
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_729
timestamp 1688980957
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_6
timestamp 1688980957
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_18
timestamp 1688980957
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_241
timestamp 1688980957
transform 1 0 23276 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_245
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1688980957
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_257
timestamp 1688980957
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_262
timestamp 1688980957
transform 1 0 25208 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_288
timestamp 1688980957
transform 1 0 27600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_300
timestamp 1688980957
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_385
timestamp 1688980957
transform 1 0 36524 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_419
timestamp 1688980957
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_437
timestamp 1688980957
transform 1 0 41308 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_443
timestamp 1688980957
transform 1 0 41860 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_477
timestamp 1688980957
transform 1 0 44988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_481
timestamp 1688980957
transform 1 0 45356 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_502
timestamp 1688980957
transform 1 0 47288 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_523
timestamp 1688980957
transform 1 0 49220 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_530
timestamp 1688980957
transform 1 0 49864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_533
timestamp 1688980957
transform 1 0 50140 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_573
timestamp 1688980957
transform 1 0 53820 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_585
timestamp 1688980957
transform 1 0 54924 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_589
timestamp 1688980957
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_601
timestamp 1688980957
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_613
timestamp 1688980957
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_625
timestamp 1688980957
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_637
timestamp 1688980957
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_643
timestamp 1688980957
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_645
timestamp 1688980957
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_657
timestamp 1688980957
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_669
timestamp 1688980957
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_681
timestamp 1688980957
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_693
timestamp 1688980957
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_699
timestamp 1688980957
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_701
timestamp 1688980957
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_713
timestamp 1688980957
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_725
timestamp 1688980957
transform 1 0 67804 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_260
timestamp 1688980957
transform 1 0 25024 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_272
timestamp 1688980957
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_289
timestamp 1688980957
transform 1 0 27692 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_296
timestamp 1688980957
transform 1 0 28336 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_324
timestamp 1688980957
transform 1 0 30912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_334
timestamp 1688980957
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_359
timestamp 1688980957
transform 1 0 34132 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_363
timestamp 1688980957
transform 1 0 34500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_375
timestamp 1688980957
transform 1 0 35604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_390
timestamp 1688980957
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_426
timestamp 1688980957
transform 1 0 40296 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_466
timestamp 1688980957
transform 1 0 43976 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_496
timestamp 1688980957
transform 1 0 46736 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_505
timestamp 1688980957
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_526
timestamp 1688980957
transform 1 0 49496 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_536
timestamp 1688980957
transform 1 0 50416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_558
timestamp 1688980957
transform 1 0 52440 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_561
timestamp 1688980957
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_573
timestamp 1688980957
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_585
timestamp 1688980957
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_597
timestamp 1688980957
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_609
timestamp 1688980957
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_615
timestamp 1688980957
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_617
timestamp 1688980957
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_629
timestamp 1688980957
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_641
timestamp 1688980957
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_653
timestamp 1688980957
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_665
timestamp 1688980957
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_671
timestamp 1688980957
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_673
timestamp 1688980957
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_685
timestamp 1688980957
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_697
timestamp 1688980957
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_709
timestamp 1688980957
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_721
timestamp 1688980957
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_727
timestamp 1688980957
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_729
timestamp 1688980957
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_261
timestamp 1688980957
transform 1 0 25116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_276
timestamp 1688980957
transform 1 0 26496 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_317
timestamp 1688980957
transform 1 0 30268 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_332
timestamp 1688980957
transform 1 0 31648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_351
timestamp 1688980957
transform 1 0 33396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_355
timestamp 1688980957
transform 1 0 33764 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_373
timestamp 1688980957
transform 1 0 35420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_385
timestamp 1688980957
transform 1 0 36524 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_394
timestamp 1688980957
transform 1 0 37352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_415
timestamp 1688980957
transform 1 0 39284 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1688980957
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_437
timestamp 1688980957
transform 1 0 41308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_447
timestamp 1688980957
transform 1 0 42228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_459
timestamp 1688980957
transform 1 0 43332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_465
timestamp 1688980957
transform 1 0 43884 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_473
timestamp 1688980957
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_477
timestamp 1688980957
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_489
timestamp 1688980957
transform 1 0 46092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_509
timestamp 1688980957
transform 1 0 47932 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_517
timestamp 1688980957
transform 1 0 48668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_525
timestamp 1688980957
transform 1 0 49404 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_529
timestamp 1688980957
transform 1 0 49772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_533
timestamp 1688980957
transform 1 0 50140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_537
timestamp 1688980957
transform 1 0 50508 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_546
timestamp 1688980957
transform 1 0 51336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_551
timestamp 1688980957
transform 1 0 51796 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_559
timestamp 1688980957
transform 1 0 52532 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_564
timestamp 1688980957
transform 1 0 52992 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_576
timestamp 1688980957
transform 1 0 54096 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_589
timestamp 1688980957
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_601
timestamp 1688980957
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_613
timestamp 1688980957
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_625
timestamp 1688980957
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_637
timestamp 1688980957
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_643
timestamp 1688980957
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_645
timestamp 1688980957
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_657
timestamp 1688980957
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_669
timestamp 1688980957
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_681
timestamp 1688980957
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_693
timestamp 1688980957
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_699
timestamp 1688980957
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_701
timestamp 1688980957
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_713
timestamp 1688980957
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_725
timestamp 1688980957
transform 1 0 67804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_729
timestamp 1688980957
transform 1 0 68172 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1688980957
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_245
timestamp 1688980957
transform 1 0 23644 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1688980957
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_324
timestamp 1688980957
transform 1 0 30912 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_355
timestamp 1688980957
transform 1 0 33764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_359
timestamp 1688980957
transform 1 0 34132 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_371
timestamp 1688980957
transform 1 0 35236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1688980957
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_411
timestamp 1688980957
transform 1 0 38916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_432
timestamp 1688980957
transform 1 0 40848 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_439
timestamp 1688980957
transform 1 0 41492 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 1688980957
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_456
timestamp 1688980957
transform 1 0 43056 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_462
timestamp 1688980957
transform 1 0 43608 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_474
timestamp 1688980957
transform 1 0 44712 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_482
timestamp 1688980957
transform 1 0 45448 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_486
timestamp 1688980957
transform 1 0 45816 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_503
timestamp 1688980957
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_539
timestamp 1688980957
transform 1 0 50692 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_581
timestamp 1688980957
transform 1 0 54556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_593
timestamp 1688980957
transform 1 0 55660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_605
timestamp 1688980957
transform 1 0 56764 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_613
timestamp 1688980957
transform 1 0 57500 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_617
timestamp 1688980957
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_629
timestamp 1688980957
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_641
timestamp 1688980957
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_653
timestamp 1688980957
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_665
timestamp 1688980957
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_671
timestamp 1688980957
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_673
timestamp 1688980957
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_685
timestamp 1688980957
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_697
timestamp 1688980957
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_709
timestamp 1688980957
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_721
timestamp 1688980957
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_727
timestamp 1688980957
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_729
timestamp 1688980957
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_259
timestamp 1688980957
transform 1 0 24932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_268
timestamp 1688980957
transform 1 0 25760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_315
timestamp 1688980957
transform 1 0 30084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_338
timestamp 1688980957
transform 1 0 32200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_358
timestamp 1688980957
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_382
timestamp 1688980957
transform 1 0 36248 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_394
timestamp 1688980957
transform 1 0 37352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_404
timestamp 1688980957
transform 1 0 38272 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_408
timestamp 1688980957
transform 1 0 38640 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_418
timestamp 1688980957
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_446
timestamp 1688980957
transform 1 0 42136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_477
timestamp 1688980957
transform 1 0 44988 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_486
timestamp 1688980957
transform 1 0 45816 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_515
timestamp 1688980957
transform 1 0 48484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_527
timestamp 1688980957
transform 1 0 49588 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_533
timestamp 1688980957
transform 1 0 50140 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_563
timestamp 1688980957
transform 1 0 52900 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_575
timestamp 1688980957
transform 1 0 54004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_587
timestamp 1688980957
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_589
timestamp 1688980957
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_601
timestamp 1688980957
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_613
timestamp 1688980957
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_625
timestamp 1688980957
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_637
timestamp 1688980957
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_643
timestamp 1688980957
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_645
timestamp 1688980957
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_657
timestamp 1688980957
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_669
timestamp 1688980957
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_681
timestamp 1688980957
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_693
timestamp 1688980957
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_699
timestamp 1688980957
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_701
timestamp 1688980957
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_713
timestamp 1688980957
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_725
timestamp 1688980957
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_6
timestamp 1688980957
transform 1 0 1656 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_18
timestamp 1688980957
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_30
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_42
timestamp 1688980957
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_261
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_267
timestamp 1688980957
transform 1 0 25668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_272
timestamp 1688980957
transform 1 0 26128 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_278
timestamp 1688980957
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_303
timestamp 1688980957
transform 1 0 28980 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_307
timestamp 1688980957
transform 1 0 29348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_316
timestamp 1688980957
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_342
timestamp 1688980957
transform 1 0 32568 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_363
timestamp 1688980957
transform 1 0 34500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_375
timestamp 1688980957
transform 1 0 35604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_387
timestamp 1688980957
transform 1 0 36708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1688980957
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_429
timestamp 1688980957
transform 1 0 40572 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_434
timestamp 1688980957
transform 1 0 41032 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_446
timestamp 1688980957
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_468
timestamp 1688980957
transform 1 0 44160 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_497
timestamp 1688980957
transform 1 0 46828 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_502
timestamp 1688980957
transform 1 0 47288 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_505
timestamp 1688980957
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_517
timestamp 1688980957
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_529
timestamp 1688980957
transform 1 0 49772 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_553
timestamp 1688980957
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_559
timestamp 1688980957
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_561
timestamp 1688980957
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_573
timestamp 1688980957
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_585
timestamp 1688980957
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_597
timestamp 1688980957
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_609
timestamp 1688980957
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_615
timestamp 1688980957
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_617
timestamp 1688980957
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_629
timestamp 1688980957
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_641
timestamp 1688980957
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_653
timestamp 1688980957
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_665
timestamp 1688980957
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_671
timestamp 1688980957
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_673
timestamp 1688980957
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_685
timestamp 1688980957
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_697
timestamp 1688980957
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_709
timestamp 1688980957
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_721
timestamp 1688980957
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_727
timestamp 1688980957
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_729
timestamp 1688980957
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_295
timestamp 1688980957
transform 1 0 28244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_327
timestamp 1688980957
transform 1 0 31188 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_339
timestamp 1688980957
transform 1 0 32292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_351
timestamp 1688980957
transform 1 0 33396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1688980957
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_371
timestamp 1688980957
transform 1 0 35236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_388
timestamp 1688980957
transform 1 0 36800 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_400
timestamp 1688980957
transform 1 0 37904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_405
timestamp 1688980957
transform 1 0 38364 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_448
timestamp 1688980957
transform 1 0 42320 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_484
timestamp 1688980957
transform 1 0 45632 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_531
timestamp 1688980957
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_533
timestamp 1688980957
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_548
timestamp 1688980957
transform 1 0 51520 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_558
timestamp 1688980957
transform 1 0 52440 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_570
timestamp 1688980957
transform 1 0 53544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_582
timestamp 1688980957
transform 1 0 54648 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_589
timestamp 1688980957
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_601
timestamp 1688980957
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_613
timestamp 1688980957
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_625
timestamp 1688980957
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_637
timestamp 1688980957
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_643
timestamp 1688980957
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_645
timestamp 1688980957
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_657
timestamp 1688980957
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_669
timestamp 1688980957
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_681
timestamp 1688980957
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_693
timestamp 1688980957
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_699
timestamp 1688980957
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_701
timestamp 1688980957
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_713
timestamp 1688980957
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_725
timestamp 1688980957
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_269
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_289
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_310
timestamp 1688980957
transform 1 0 29624 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_316
timestamp 1688980957
transform 1 0 30176 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_320
timestamp 1688980957
transform 1 0 30544 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_328
timestamp 1688980957
transform 1 0 31280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_370
timestamp 1688980957
transform 1 0 35144 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_379
timestamp 1688980957
transform 1 0 35972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_384
timestamp 1688980957
transform 1 0 36432 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_405
timestamp 1688980957
transform 1 0 38364 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_416
timestamp 1688980957
transform 1 0 39376 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_441
timestamp 1688980957
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_447
timestamp 1688980957
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_449
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_477
timestamp 1688980957
transform 1 0 44988 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_489
timestamp 1688980957
transform 1 0 46092 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_499
timestamp 1688980957
transform 1 0 47012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_503
timestamp 1688980957
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_505
timestamp 1688980957
transform 1 0 47564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_511
timestamp 1688980957
transform 1 0 48116 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_535
timestamp 1688980957
transform 1 0 50324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_547
timestamp 1688980957
transform 1 0 51428 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_559
timestamp 1688980957
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_561
timestamp 1688980957
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_573
timestamp 1688980957
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_585
timestamp 1688980957
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_597
timestamp 1688980957
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_609
timestamp 1688980957
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_615
timestamp 1688980957
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_617
timestamp 1688980957
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_629
timestamp 1688980957
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_641
timestamp 1688980957
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_653
timestamp 1688980957
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_665
timestamp 1688980957
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_671
timestamp 1688980957
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_673
timestamp 1688980957
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_685
timestamp 1688980957
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_697
timestamp 1688980957
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_709
timestamp 1688980957
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_721
timestamp 1688980957
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_727
timestamp 1688980957
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_729
timestamp 1688980957
transform 1 0 68172 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_297
timestamp 1688980957
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_301
timestamp 1688980957
transform 1 0 28796 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_373
timestamp 1688980957
transform 1 0 35420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 1688980957
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 1688980957
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_445
timestamp 1688980957
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_457
timestamp 1688980957
transform 1 0 43148 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_472
timestamp 1688980957
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_477
timestamp 1688980957
transform 1 0 44988 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_494
timestamp 1688980957
transform 1 0 46552 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_526
timestamp 1688980957
transform 1 0 49496 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_533
timestamp 1688980957
transform 1 0 50140 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_540
timestamp 1688980957
transform 1 0 50784 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_552
timestamp 1688980957
transform 1 0 51888 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_564
timestamp 1688980957
transform 1 0 52992 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_576
timestamp 1688980957
transform 1 0 54096 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_589
timestamp 1688980957
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_601
timestamp 1688980957
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_613
timestamp 1688980957
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_625
timestamp 1688980957
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_637
timestamp 1688980957
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_643
timestamp 1688980957
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_645
timestamp 1688980957
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_657
timestamp 1688980957
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_669
timestamp 1688980957
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_681
timestamp 1688980957
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_693
timestamp 1688980957
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_699
timestamp 1688980957
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_701
timestamp 1688980957
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_713
timestamp 1688980957
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_725
timestamp 1688980957
transform 1 0 67804 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1688980957
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_287
timestamp 1688980957
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_296
timestamp 1688980957
transform 1 0 28336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_300
timestamp 1688980957
transform 1 0 28704 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_322
timestamp 1688980957
transform 1 0 30728 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_332
timestamp 1688980957
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_360
timestamp 1688980957
transform 1 0 34224 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_368
timestamp 1688980957
transform 1 0 34960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_387
timestamp 1688980957
transform 1 0 36708 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_409
timestamp 1688980957
transform 1 0 38732 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_426
timestamp 1688980957
transform 1 0 40296 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_465
timestamp 1688980957
transform 1 0 43884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_551
timestamp 1688980957
transform 1 0 51796 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_559
timestamp 1688980957
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_561
timestamp 1688980957
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_573
timestamp 1688980957
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_585
timestamp 1688980957
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_597
timestamp 1688980957
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_609
timestamp 1688980957
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_615
timestamp 1688980957
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_617
timestamp 1688980957
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_629
timestamp 1688980957
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_641
timestamp 1688980957
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_653
timestamp 1688980957
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_665
timestamp 1688980957
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_671
timestamp 1688980957
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_673
timestamp 1688980957
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_685
timestamp 1688980957
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_697
timestamp 1688980957
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_709
timestamp 1688980957
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_721
timestamp 1688980957
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_727
timestamp 1688980957
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_729
timestamp 1688980957
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_6
timestamp 1688980957
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 1688980957
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1688980957
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_325
timestamp 1688980957
transform 1 0 31004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_334
timestamp 1688980957
transform 1 0 31832 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_342
timestamp 1688980957
transform 1 0 32568 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_362
timestamp 1688980957
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_376
timestamp 1688980957
transform 1 0 35696 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_387
timestamp 1688980957
transform 1 0 36708 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_408
timestamp 1688980957
transform 1 0 38640 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_418
timestamp 1688980957
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_447
timestamp 1688980957
transform 1 0 42228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_462
timestamp 1688980957
transform 1 0 43608 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_466
timestamp 1688980957
transform 1 0 43976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_471
timestamp 1688980957
transform 1 0 44436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_490
timestamp 1688980957
transform 1 0 46184 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_495
timestamp 1688980957
transform 1 0 46644 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_505
timestamp 1688980957
transform 1 0 47564 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_523
timestamp 1688980957
transform 1 0 49220 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_531
timestamp 1688980957
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_545
timestamp 1688980957
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_557
timestamp 1688980957
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_569
timestamp 1688980957
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_581
timestamp 1688980957
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_587
timestamp 1688980957
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 1688980957
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_601
timestamp 1688980957
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_613
timestamp 1688980957
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_625
timestamp 1688980957
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_637
timestamp 1688980957
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_643
timestamp 1688980957
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_645
timestamp 1688980957
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_657
timestamp 1688980957
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_669
timestamp 1688980957
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_681
timestamp 1688980957
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_693
timestamp 1688980957
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_699
timestamp 1688980957
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_701
timestamp 1688980957
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_713
timestamp 1688980957
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_725
timestamp 1688980957
transform 1 0 67804 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_269
timestamp 1688980957
transform 1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_275
timestamp 1688980957
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_302
timestamp 1688980957
transform 1 0 28888 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_306
timestamp 1688980957
transform 1 0 29256 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_318
timestamp 1688980957
transform 1 0 30360 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_330
timestamp 1688980957
transform 1 0 31464 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_376
timestamp 1688980957
transform 1 0 35696 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_387
timestamp 1688980957
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_401
timestamp 1688980957
transform 1 0 37996 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_413
timestamp 1688980957
transform 1 0 39100 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_422
timestamp 1688980957
transform 1 0 39928 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_434
timestamp 1688980957
transform 1 0 41032 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_453
timestamp 1688980957
transform 1 0 42780 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_467
timestamp 1688980957
transform 1 0 44068 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_479
timestamp 1688980957
transform 1 0 45172 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_495
timestamp 1688980957
transform 1 0 46644 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_503
timestamp 1688980957
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_510
timestamp 1688980957
transform 1 0 48024 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_522
timestamp 1688980957
transform 1 0 49128 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_530
timestamp 1688980957
transform 1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_539
timestamp 1688980957
transform 1 0 50692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_551
timestamp 1688980957
transform 1 0 51796 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_559
timestamp 1688980957
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_561
timestamp 1688980957
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_573
timestamp 1688980957
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_585
timestamp 1688980957
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_597
timestamp 1688980957
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_609
timestamp 1688980957
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_615
timestamp 1688980957
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_617
timestamp 1688980957
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_629
timestamp 1688980957
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_641
timestamp 1688980957
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_653
timestamp 1688980957
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_665
timestamp 1688980957
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_671
timestamp 1688980957
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_673
timestamp 1688980957
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_685
timestamp 1688980957
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_697
timestamp 1688980957
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_709
timestamp 1688980957
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_721
timestamp 1688980957
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_727
timestamp 1688980957
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_729
timestamp 1688980957
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_273
timestamp 1688980957
transform 1 0 26220 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_278
timestamp 1688980957
transform 1 0 26680 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_288
timestamp 1688980957
transform 1 0 27600 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_314
timestamp 1688980957
transform 1 0 29992 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_320
timestamp 1688980957
transform 1 0 30544 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_327
timestamp 1688980957
transform 1 0 31188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_337
timestamp 1688980957
transform 1 0 32108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_358
timestamp 1688980957
transform 1 0 34040 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_369
timestamp 1688980957
transform 1 0 35052 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_411
timestamp 1688980957
transform 1 0 38916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_417
timestamp 1688980957
transform 1 0 39468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_440
timestamp 1688980957
transform 1 0 41584 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_448
timestamp 1688980957
transform 1 0 42320 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_452
timestamp 1688980957
transform 1 0 42688 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_463
timestamp 1688980957
transform 1 0 43700 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_469
timestamp 1688980957
transform 1 0 44252 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_501
timestamp 1688980957
transform 1 0 47196 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_507
timestamp 1688980957
transform 1 0 47748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_514
timestamp 1688980957
transform 1 0 48392 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_522
timestamp 1688980957
transform 1 0 49128 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_556
timestamp 1688980957
transform 1 0 52256 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_568
timestamp 1688980957
transform 1 0 53360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_580
timestamp 1688980957
transform 1 0 54464 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_589
timestamp 1688980957
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_601
timestamp 1688980957
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_613
timestamp 1688980957
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_625
timestamp 1688980957
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_637
timestamp 1688980957
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_643
timestamp 1688980957
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_645
timestamp 1688980957
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_657
timestamp 1688980957
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_669
timestamp 1688980957
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_681
timestamp 1688980957
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_693
timestamp 1688980957
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_699
timestamp 1688980957
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_701
timestamp 1688980957
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_713
timestamp 1688980957
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_725
timestamp 1688980957
transform 1 0 67804 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_729
timestamp 1688980957
transform 1 0 68172 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_257
timestamp 1688980957
transform 1 0 24748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_296
timestamp 1688980957
transform 1 0 28336 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_333
timestamp 1688980957
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_377
timestamp 1688980957
transform 1 0 35788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_381
timestamp 1688980957
transform 1 0 36156 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1688980957
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_441
timestamp 1688980957
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 1688980957
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_449
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_482
timestamp 1688980957
transform 1 0 45448 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_494
timestamp 1688980957
transform 1 0 46552 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_505
timestamp 1688980957
transform 1 0 47564 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_522
timestamp 1688980957
transform 1 0 49128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_530
timestamp 1688980957
transform 1 0 49864 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_536
timestamp 1688980957
transform 1 0 50416 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_548
timestamp 1688980957
transform 1 0 51520 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_561
timestamp 1688980957
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_573
timestamp 1688980957
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_585
timestamp 1688980957
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_597
timestamp 1688980957
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_609
timestamp 1688980957
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_615
timestamp 1688980957
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_617
timestamp 1688980957
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_629
timestamp 1688980957
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_641
timestamp 1688980957
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_653
timestamp 1688980957
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_665
timestamp 1688980957
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_671
timestamp 1688980957
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_673
timestamp 1688980957
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_685
timestamp 1688980957
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_697
timestamp 1688980957
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_709
timestamp 1688980957
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_721
timestamp 1688980957
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_727
timestamp 1688980957
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_729
timestamp 1688980957
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_261
timestamp 1688980957
transform 1 0 25116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_275
timestamp 1688980957
transform 1 0 26404 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_284
timestamp 1688980957
transform 1 0 27232 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_296
timestamp 1688980957
transform 1 0 28336 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_316
timestamp 1688980957
transform 1 0 30176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_328
timestamp 1688980957
transform 1 0 31280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_360
timestamp 1688980957
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_381
timestamp 1688980957
transform 1 0 36156 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_387
timestamp 1688980957
transform 1 0 36708 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_391
timestamp 1688980957
transform 1 0 37076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_399
timestamp 1688980957
transform 1 0 37812 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_408
timestamp 1688980957
transform 1 0 38640 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_413
timestamp 1688980957
transform 1 0 39100 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_468
timestamp 1688980957
transform 1 0 44160 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_474
timestamp 1688980957
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_477
timestamp 1688980957
transform 1 0 44988 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_485
timestamp 1688980957
transform 1 0 45724 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_509
timestamp 1688980957
transform 1 0 47932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_515
timestamp 1688980957
transform 1 0 48484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_531
timestamp 1688980957
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_540
timestamp 1688980957
transform 1 0 50784 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_552
timestamp 1688980957
transform 1 0 51888 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_564
timestamp 1688980957
transform 1 0 52992 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_576
timestamp 1688980957
transform 1 0 54096 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_589
timestamp 1688980957
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_601
timestamp 1688980957
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_613
timestamp 1688980957
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_625
timestamp 1688980957
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_637
timestamp 1688980957
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_643
timestamp 1688980957
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_645
timestamp 1688980957
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_657
timestamp 1688980957
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_669
timestamp 1688980957
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_681
timestamp 1688980957
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_693
timestamp 1688980957
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_699
timestamp 1688980957
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_701
timestamp 1688980957
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_713
timestamp 1688980957
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_725
timestamp 1688980957
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_9
timestamp 1688980957
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_21
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_33
timestamp 1688980957
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_45
timestamp 1688980957
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_316
timestamp 1688980957
transform 1 0 30176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_320
timestamp 1688980957
transform 1 0 30544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_326
timestamp 1688980957
transform 1 0 31096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_334
timestamp 1688980957
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_371
timestamp 1688980957
transform 1 0 35236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1688980957
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_412
timestamp 1688980957
transform 1 0 39008 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_424
timestamp 1688980957
transform 1 0 40112 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_436
timestamp 1688980957
transform 1 0 41216 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_452
timestamp 1688980957
transform 1 0 42688 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_460
timestamp 1688980957
transform 1 0 43424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_505
timestamp 1688980957
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_510
timestamp 1688980957
transform 1 0 48024 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_549
timestamp 1688980957
transform 1 0 51612 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_557
timestamp 1688980957
transform 1 0 52348 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_561
timestamp 1688980957
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_573
timestamp 1688980957
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_585
timestamp 1688980957
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_597
timestamp 1688980957
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_609
timestamp 1688980957
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_615
timestamp 1688980957
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_617
timestamp 1688980957
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_629
timestamp 1688980957
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_641
timestamp 1688980957
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_653
timestamp 1688980957
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_665
timestamp 1688980957
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_671
timestamp 1688980957
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_673
timestamp 1688980957
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_685
timestamp 1688980957
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_697
timestamp 1688980957
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_709
timestamp 1688980957
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_721
timestamp 1688980957
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_727
timestamp 1688980957
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_729
timestamp 1688980957
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_283
timestamp 1688980957
transform 1 0 27140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_292
timestamp 1688980957
transform 1 0 27968 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 1688980957
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_315
timestamp 1688980957
transform 1 0 30084 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_332
timestamp 1688980957
transform 1 0 31648 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_344
timestamp 1688980957
transform 1 0 32752 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_356
timestamp 1688980957
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_377
timestamp 1688980957
transform 1 0 35788 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_394
timestamp 1688980957
transform 1 0 37352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_415
timestamp 1688980957
transform 1 0 39284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1688980957
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_433
timestamp 1688980957
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_445
timestamp 1688980957
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_457
timestamp 1688980957
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_469
timestamp 1688980957
transform 1 0 44252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_477
timestamp 1688980957
transform 1 0 44988 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_500
timestamp 1688980957
transform 1 0 47104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_524
timestamp 1688980957
transform 1 0 49312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_530
timestamp 1688980957
transform 1 0 49864 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_533
timestamp 1688980957
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_545
timestamp 1688980957
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_557
timestamp 1688980957
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_569
timestamp 1688980957
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_581
timestamp 1688980957
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_587
timestamp 1688980957
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_589
timestamp 1688980957
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_601
timestamp 1688980957
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_613
timestamp 1688980957
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_625
timestamp 1688980957
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_637
timestamp 1688980957
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_643
timestamp 1688980957
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_645
timestamp 1688980957
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_657
timestamp 1688980957
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_669
timestamp 1688980957
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_681
timestamp 1688980957
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_693
timestamp 1688980957
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_699
timestamp 1688980957
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_701
timestamp 1688980957
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_713
timestamp 1688980957
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_725
timestamp 1688980957
transform 1 0 67804 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_286
timestamp 1688980957
transform 1 0 27416 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_298
timestamp 1688980957
transform 1 0 28520 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_310
timestamp 1688980957
transform 1 0 29624 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_314
timestamp 1688980957
transform 1 0 29992 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_318
timestamp 1688980957
transform 1 0 30360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_351
timestamp 1688980957
transform 1 0 33396 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_357
timestamp 1688980957
transform 1 0 33948 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_374
timestamp 1688980957
transform 1 0 35512 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_386
timestamp 1688980957
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_411
timestamp 1688980957
transform 1 0 38916 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_423
timestamp 1688980957
transform 1 0 40020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_435
timestamp 1688980957
transform 1 0 41124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_447
timestamp 1688980957
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 1688980957
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_461
timestamp 1688980957
transform 1 0 43516 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_487
timestamp 1688980957
transform 1 0 45908 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_500
timestamp 1688980957
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_513
timestamp 1688980957
transform 1 0 48300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_517
timestamp 1688980957
transform 1 0 48668 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_526
timestamp 1688980957
transform 1 0 49496 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_538
timestamp 1688980957
transform 1 0 50600 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_550
timestamp 1688980957
transform 1 0 51704 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_558
timestamp 1688980957
transform 1 0 52440 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_561
timestamp 1688980957
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_573
timestamp 1688980957
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_585
timestamp 1688980957
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_597
timestamp 1688980957
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_609
timestamp 1688980957
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_615
timestamp 1688980957
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_617
timestamp 1688980957
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_629
timestamp 1688980957
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_641
timestamp 1688980957
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_653
timestamp 1688980957
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_665
timestamp 1688980957
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_671
timestamp 1688980957
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_673
timestamp 1688980957
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_685
timestamp 1688980957
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_697
timestamp 1688980957
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_709
timestamp 1688980957
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_721
timestamp 1688980957
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_727
timestamp 1688980957
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_729
timestamp 1688980957
transform 1 0 68172 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_293
timestamp 1688980957
transform 1 0 28060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_297
timestamp 1688980957
transform 1 0 28428 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_319
timestamp 1688980957
transform 1 0 30452 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_356
timestamp 1688980957
transform 1 0 33856 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_360
timestamp 1688980957
transform 1 0 34224 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_371
timestamp 1688980957
transform 1 0 35236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_385
timestamp 1688980957
transform 1 0 36524 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_396
timestamp 1688980957
transform 1 0 37536 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_402
timestamp 1688980957
transform 1 0 38088 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 1688980957
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_421
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_433
timestamp 1688980957
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_445
timestamp 1688980957
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_457
timestamp 1688980957
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_469
timestamp 1688980957
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_475
timestamp 1688980957
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_480
timestamp 1688980957
transform 1 0 45264 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_503
timestamp 1688980957
transform 1 0 47380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_529
timestamp 1688980957
transform 1 0 49772 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_533
timestamp 1688980957
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_545
timestamp 1688980957
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_557
timestamp 1688980957
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_569
timestamp 1688980957
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_581
timestamp 1688980957
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_587
timestamp 1688980957
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_589
timestamp 1688980957
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_601
timestamp 1688980957
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_613
timestamp 1688980957
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_625
timestamp 1688980957
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_637
timestamp 1688980957
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_643
timestamp 1688980957
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_645
timestamp 1688980957
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_657
timestamp 1688980957
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_669
timestamp 1688980957
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_681
timestamp 1688980957
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_693
timestamp 1688980957
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_699
timestamp 1688980957
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_701
timestamp 1688980957
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_713
timestamp 1688980957
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_725
timestamp 1688980957
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_284
timestamp 1688980957
transform 1 0 27232 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_292
timestamp 1688980957
transform 1 0 27968 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_311
timestamp 1688980957
transform 1 0 29716 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_324
timestamp 1688980957
transform 1 0 30912 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_334
timestamp 1688980957
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_345
timestamp 1688980957
transform 1 0 32844 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_357
timestamp 1688980957
transform 1 0 33948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_383
timestamp 1688980957
transform 1 0 36340 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_406
timestamp 1688980957
transform 1 0 38456 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_423
timestamp 1688980957
transform 1 0 40020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_435
timestamp 1688980957
transform 1 0 41124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 1688980957
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_449
timestamp 1688980957
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_461
timestamp 1688980957
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_473
timestamp 1688980957
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_485
timestamp 1688980957
transform 1 0 45724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_498
timestamp 1688980957
transform 1 0 46920 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_505
timestamp 1688980957
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_517
timestamp 1688980957
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_529
timestamp 1688980957
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_541
timestamp 1688980957
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_553
timestamp 1688980957
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_559
timestamp 1688980957
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_561
timestamp 1688980957
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_573
timestamp 1688980957
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_585
timestamp 1688980957
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_597
timestamp 1688980957
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_609
timestamp 1688980957
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 1688980957
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_617
timestamp 1688980957
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_629
timestamp 1688980957
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_641
timestamp 1688980957
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_653
timestamp 1688980957
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_665
timestamp 1688980957
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_671
timestamp 1688980957
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_673
timestamp 1688980957
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_685
timestamp 1688980957
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_697
timestamp 1688980957
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_709
timestamp 1688980957
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_721
timestamp 1688980957
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_727
timestamp 1688980957
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_729
timestamp 1688980957
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_6
timestamp 1688980957
transform 1 0 1656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_18
timestamp 1688980957
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_26
timestamp 1688980957
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_305
timestamp 1688980957
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_324
timestamp 1688980957
transform 1 0 30912 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_350
timestamp 1688980957
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_362
timestamp 1688980957
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_371
timestamp 1688980957
transform 1 0 35236 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_384
timestamp 1688980957
transform 1 0 36432 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_410
timestamp 1688980957
transform 1 0 38824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_418
timestamp 1688980957
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_433
timestamp 1688980957
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_445
timestamp 1688980957
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_457
timestamp 1688980957
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_469
timestamp 1688980957
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_475
timestamp 1688980957
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_477
timestamp 1688980957
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_489
timestamp 1688980957
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_501
timestamp 1688980957
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_513
timestamp 1688980957
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_525
timestamp 1688980957
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_531
timestamp 1688980957
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_533
timestamp 1688980957
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_545
timestamp 1688980957
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_557
timestamp 1688980957
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_569
timestamp 1688980957
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_581
timestamp 1688980957
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_587
timestamp 1688980957
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_589
timestamp 1688980957
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_601
timestamp 1688980957
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_613
timestamp 1688980957
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_625
timestamp 1688980957
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_637
timestamp 1688980957
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_643
timestamp 1688980957
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_645
timestamp 1688980957
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_657
timestamp 1688980957
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_669
timestamp 1688980957
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_681
timestamp 1688980957
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_693
timestamp 1688980957
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_699
timestamp 1688980957
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_701
timestamp 1688980957
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_713
timestamp 1688980957
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_725
timestamp 1688980957
transform 1 0 67804 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_310
timestamp 1688980957
transform 1 0 29624 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_330
timestamp 1688980957
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_389
timestamp 1688980957
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_401
timestamp 1688980957
transform 1 0 37996 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_413
timestamp 1688980957
transform 1 0 39100 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_425
timestamp 1688980957
transform 1 0 40204 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_437
timestamp 1688980957
transform 1 0 41308 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_445
timestamp 1688980957
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_461
timestamp 1688980957
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_473
timestamp 1688980957
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_485
timestamp 1688980957
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_497
timestamp 1688980957
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 1688980957
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_505
timestamp 1688980957
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_517
timestamp 1688980957
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_529
timestamp 1688980957
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_541
timestamp 1688980957
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_553
timestamp 1688980957
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_559
timestamp 1688980957
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_561
timestamp 1688980957
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_573
timestamp 1688980957
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_585
timestamp 1688980957
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_597
timestamp 1688980957
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_609
timestamp 1688980957
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_615
timestamp 1688980957
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_617
timestamp 1688980957
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_629
timestamp 1688980957
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_641
timestamp 1688980957
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_653
timestamp 1688980957
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_665
timestamp 1688980957
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_671
timestamp 1688980957
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_673
timestamp 1688980957
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_685
timestamp 1688980957
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_697
timestamp 1688980957
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_709
timestamp 1688980957
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_721
timestamp 1688980957
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_727
timestamp 1688980957
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_729
timestamp 1688980957
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_297
timestamp 1688980957
transform 1 0 28428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_303
timestamp 1688980957
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_325
timestamp 1688980957
transform 1 0 31004 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_334
timestamp 1688980957
transform 1 0 31832 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_346
timestamp 1688980957
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_358
timestamp 1688980957
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 1688980957
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 1688980957
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1688980957
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 1688980957
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 1688980957
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_457
timestamp 1688980957
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_469
timestamp 1688980957
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_475
timestamp 1688980957
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_477
timestamp 1688980957
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_489
timestamp 1688980957
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_501
timestamp 1688980957
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_513
timestamp 1688980957
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 1688980957
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 1688980957
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 1688980957
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_545
timestamp 1688980957
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_557
timestamp 1688980957
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_569
timestamp 1688980957
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_581
timestamp 1688980957
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_587
timestamp 1688980957
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_589
timestamp 1688980957
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_601
timestamp 1688980957
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_613
timestamp 1688980957
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_625
timestamp 1688980957
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_637
timestamp 1688980957
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_643
timestamp 1688980957
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_645
timestamp 1688980957
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_657
timestamp 1688980957
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_669
timestamp 1688980957
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_681
timestamp 1688980957
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_693
timestamp 1688980957
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_699
timestamp 1688980957
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_701
timestamp 1688980957
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_713
timestamp 1688980957
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_725
timestamp 1688980957
transform 1 0 67804 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_729
timestamp 1688980957
transform 1 0 68172 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1688980957
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1688980957
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 1688980957
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 1688980957
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 1688980957
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 1688980957
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_461
timestamp 1688980957
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_473
timestamp 1688980957
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_485
timestamp 1688980957
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_497
timestamp 1688980957
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 1688980957
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_505
timestamp 1688980957
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_517
timestamp 1688980957
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_529
timestamp 1688980957
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_541
timestamp 1688980957
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_553
timestamp 1688980957
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_559
timestamp 1688980957
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_561
timestamp 1688980957
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_573
timestamp 1688980957
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_585
timestamp 1688980957
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_597
timestamp 1688980957
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_609
timestamp 1688980957
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_615
timestamp 1688980957
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_617
timestamp 1688980957
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_629
timestamp 1688980957
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_641
timestamp 1688980957
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_653
timestamp 1688980957
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_665
timestamp 1688980957
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_671
timestamp 1688980957
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_673
timestamp 1688980957
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_685
timestamp 1688980957
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_697
timestamp 1688980957
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_709
timestamp 1688980957
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_721
timestamp 1688980957
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_727
timestamp 1688980957
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_729
timestamp 1688980957
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1688980957
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1688980957
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 1688980957
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 1688980957
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 1688980957
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 1688980957
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_457
timestamp 1688980957
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_469
timestamp 1688980957
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_475
timestamp 1688980957
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_477
timestamp 1688980957
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_489
timestamp 1688980957
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_501
timestamp 1688980957
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_513
timestamp 1688980957
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_525
timestamp 1688980957
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_531
timestamp 1688980957
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_533
timestamp 1688980957
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_545
timestamp 1688980957
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_557
timestamp 1688980957
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_569
timestamp 1688980957
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_581
timestamp 1688980957
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_587
timestamp 1688980957
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 1688980957
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 1688980957
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_613
timestamp 1688980957
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_625
timestamp 1688980957
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_637
timestamp 1688980957
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_643
timestamp 1688980957
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_645
timestamp 1688980957
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_657
timestamp 1688980957
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_669
timestamp 1688980957
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_681
timestamp 1688980957
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_693
timestamp 1688980957
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_699
timestamp 1688980957
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_701
timestamp 1688980957
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_713
timestamp 1688980957
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_725
timestamp 1688980957
transform 1 0 67804 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_6
timestamp 1688980957
transform 1 0 1656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_18
timestamp 1688980957
transform 1 0 2760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_30
timestamp 1688980957
transform 1 0 3864 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_42
timestamp 1688980957
transform 1 0 4968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 1688980957
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1688980957
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1688980957
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1688980957
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1688980957
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 1688980957
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 1688980957
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 1688980957
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 1688980957
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_461
timestamp 1688980957
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_473
timestamp 1688980957
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_485
timestamp 1688980957
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_497
timestamp 1688980957
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 1688980957
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_505
timestamp 1688980957
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_517
timestamp 1688980957
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_529
timestamp 1688980957
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_541
timestamp 1688980957
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_553
timestamp 1688980957
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 1688980957
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_561
timestamp 1688980957
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_573
timestamp 1688980957
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_585
timestamp 1688980957
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_597
timestamp 1688980957
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_609
timestamp 1688980957
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_615
timestamp 1688980957
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_617
timestamp 1688980957
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_629
timestamp 1688980957
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_641
timestamp 1688980957
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_653
timestamp 1688980957
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_665
timestamp 1688980957
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_671
timestamp 1688980957
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_673
timestamp 1688980957
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_685
timestamp 1688980957
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_697
timestamp 1688980957
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_709
timestamp 1688980957
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_721
timestamp 1688980957
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_727
timestamp 1688980957
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_729
timestamp 1688980957
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1688980957
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1688980957
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1688980957
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1688980957
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 1688980957
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1688980957
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_401
timestamp 1688980957
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_413
timestamp 1688980957
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 1688980957
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 1688980957
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_445
timestamp 1688980957
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_457
timestamp 1688980957
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_469
timestamp 1688980957
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_475
timestamp 1688980957
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 1688980957
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 1688980957
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_501
timestamp 1688980957
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_513
timestamp 1688980957
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_525
timestamp 1688980957
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_531
timestamp 1688980957
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 1688980957
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_545
timestamp 1688980957
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_557
timestamp 1688980957
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_569
timestamp 1688980957
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_581
timestamp 1688980957
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_587
timestamp 1688980957
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 1688980957
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 1688980957
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_613
timestamp 1688980957
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_625
timestamp 1688980957
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_637
timestamp 1688980957
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_643
timestamp 1688980957
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_645
timestamp 1688980957
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_657
timestamp 1688980957
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_669
timestamp 1688980957
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_681
timestamp 1688980957
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_693
timestamp 1688980957
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_699
timestamp 1688980957
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_701
timestamp 1688980957
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_713
timestamp 1688980957
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_725
timestamp 1688980957
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 1688980957
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 1688980957
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1688980957
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 1688980957
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 1688980957
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_429
timestamp 1688980957
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_441
timestamp 1688980957
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_447
timestamp 1688980957
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_449
timestamp 1688980957
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_461
timestamp 1688980957
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_473
timestamp 1688980957
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_485
timestamp 1688980957
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_497
timestamp 1688980957
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_503
timestamp 1688980957
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_505
timestamp 1688980957
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_517
timestamp 1688980957
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_529
timestamp 1688980957
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_541
timestamp 1688980957
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_553
timestamp 1688980957
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_559
timestamp 1688980957
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_561
timestamp 1688980957
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_573
timestamp 1688980957
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_585
timestamp 1688980957
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_597
timestamp 1688980957
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_609
timestamp 1688980957
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_615
timestamp 1688980957
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_617
timestamp 1688980957
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_629
timestamp 1688980957
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_641
timestamp 1688980957
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_653
timestamp 1688980957
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_665
timestamp 1688980957
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_671
timestamp 1688980957
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_673
timestamp 1688980957
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_685
timestamp 1688980957
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_697
timestamp 1688980957
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_709
timestamp 1688980957
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_721
timestamp 1688980957
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_727
timestamp 1688980957
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_729
timestamp 1688980957
transform 1 0 68172 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1688980957
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1688980957
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 1688980957
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 1688980957
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_401
timestamp 1688980957
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_413
timestamp 1688980957
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 1688980957
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 1688980957
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_433
timestamp 1688980957
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_445
timestamp 1688980957
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_457
timestamp 1688980957
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_469
timestamp 1688980957
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_475
timestamp 1688980957
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_477
timestamp 1688980957
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_489
timestamp 1688980957
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_501
timestamp 1688980957
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_513
timestamp 1688980957
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_525
timestamp 1688980957
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_531
timestamp 1688980957
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_533
timestamp 1688980957
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_545
timestamp 1688980957
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_557
timestamp 1688980957
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_569
timestamp 1688980957
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_581
timestamp 1688980957
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_587
timestamp 1688980957
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_589
timestamp 1688980957
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_601
timestamp 1688980957
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_613
timestamp 1688980957
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_625
timestamp 1688980957
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_637
timestamp 1688980957
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_643
timestamp 1688980957
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_645
timestamp 1688980957
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_657
timestamp 1688980957
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_669
timestamp 1688980957
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_681
timestamp 1688980957
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_693
timestamp 1688980957
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_699
timestamp 1688980957
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_701
timestamp 1688980957
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_713
timestamp 1688980957
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_725
timestamp 1688980957
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1688980957
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 1688980957
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 1688980957
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1688980957
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_405
timestamp 1688980957
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_417
timestamp 1688980957
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_429
timestamp 1688980957
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_441
timestamp 1688980957
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_447
timestamp 1688980957
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_449
timestamp 1688980957
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_461
timestamp 1688980957
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_473
timestamp 1688980957
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_485
timestamp 1688980957
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_497
timestamp 1688980957
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_503
timestamp 1688980957
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_505
timestamp 1688980957
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_517
timestamp 1688980957
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_529
timestamp 1688980957
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_541
timestamp 1688980957
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_553
timestamp 1688980957
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_559
timestamp 1688980957
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_561
timestamp 1688980957
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_573
timestamp 1688980957
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_585
timestamp 1688980957
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_597
timestamp 1688980957
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_609
timestamp 1688980957
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_615
timestamp 1688980957
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_617
timestamp 1688980957
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_629
timestamp 1688980957
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_641
timestamp 1688980957
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_653
timestamp 1688980957
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_665
timestamp 1688980957
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_671
timestamp 1688980957
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_673
timestamp 1688980957
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_685
timestamp 1688980957
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_697
timestamp 1688980957
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_709
timestamp 1688980957
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_721
timestamp 1688980957
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_727
timestamp 1688980957
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_729
timestamp 1688980957
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_6
timestamp 1688980957
transform 1 0 1656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_18
timestamp 1688980957
transform 1 0 2760 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_26
timestamp 1688980957
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1688980957
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 1688980957
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 1688980957
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_401
timestamp 1688980957
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_413
timestamp 1688980957
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_419
timestamp 1688980957
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 1688980957
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 1688980957
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_445
timestamp 1688980957
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_457
timestamp 1688980957
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_469
timestamp 1688980957
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_475
timestamp 1688980957
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_477
timestamp 1688980957
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_489
timestamp 1688980957
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_501
timestamp 1688980957
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_513
timestamp 1688980957
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_525
timestamp 1688980957
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_531
timestamp 1688980957
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_533
timestamp 1688980957
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_545
timestamp 1688980957
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_557
timestamp 1688980957
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_569
timestamp 1688980957
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_581
timestamp 1688980957
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_587
timestamp 1688980957
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_589
timestamp 1688980957
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_601
timestamp 1688980957
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_613
timestamp 1688980957
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_625
timestamp 1688980957
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_637
timestamp 1688980957
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_643
timestamp 1688980957
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_645
timestamp 1688980957
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_657
timestamp 1688980957
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_669
timestamp 1688980957
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_681
timestamp 1688980957
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_693
timestamp 1688980957
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_699
timestamp 1688980957
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_701
timestamp 1688980957
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_713
timestamp 1688980957
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_725
timestamp 1688980957
transform 1 0 67804 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1688980957
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1688980957
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1688980957
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 1688980957
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_429
timestamp 1688980957
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_441
timestamp 1688980957
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_447
timestamp 1688980957
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_449
timestamp 1688980957
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_461
timestamp 1688980957
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_473
timestamp 1688980957
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_485
timestamp 1688980957
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_497
timestamp 1688980957
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_503
timestamp 1688980957
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_505
timestamp 1688980957
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_517
timestamp 1688980957
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_529
timestamp 1688980957
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_541
timestamp 1688980957
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_553
timestamp 1688980957
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_559
timestamp 1688980957
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_561
timestamp 1688980957
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_573
timestamp 1688980957
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_585
timestamp 1688980957
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_597
timestamp 1688980957
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_609
timestamp 1688980957
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_615
timestamp 1688980957
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_617
timestamp 1688980957
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_629
timestamp 1688980957
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_641
timestamp 1688980957
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_653
timestamp 1688980957
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_665
timestamp 1688980957
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_671
timestamp 1688980957
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_673
timestamp 1688980957
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_685
timestamp 1688980957
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_697
timestamp 1688980957
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_709
timestamp 1688980957
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_721
timestamp 1688980957
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_727
timestamp 1688980957
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_729
timestamp 1688980957
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1688980957
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1688980957
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_401
timestamp 1688980957
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_413
timestamp 1688980957
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 1688980957
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 1688980957
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_433
timestamp 1688980957
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_445
timestamp 1688980957
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_457
timestamp 1688980957
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_469
timestamp 1688980957
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_475
timestamp 1688980957
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_477
timestamp 1688980957
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_489
timestamp 1688980957
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_501
timestamp 1688980957
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_513
timestamp 1688980957
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_525
timestamp 1688980957
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_531
timestamp 1688980957
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_533
timestamp 1688980957
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_545
timestamp 1688980957
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_557
timestamp 1688980957
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_569
timestamp 1688980957
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_581
timestamp 1688980957
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_587
timestamp 1688980957
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_589
timestamp 1688980957
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_601
timestamp 1688980957
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_613
timestamp 1688980957
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_625
timestamp 1688980957
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_637
timestamp 1688980957
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_643
timestamp 1688980957
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_645
timestamp 1688980957
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_657
timestamp 1688980957
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_669
timestamp 1688980957
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_681
timestamp 1688980957
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_693
timestamp 1688980957
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_699
timestamp 1688980957
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_701
timestamp 1688980957
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_713
timestamp 1688980957
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_725
timestamp 1688980957
transform 1 0 67804 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_729
timestamp 1688980957
transform 1 0 68172 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1688980957
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 1688980957
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1688980957
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 1688980957
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 1688980957
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_429
timestamp 1688980957
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_441
timestamp 1688980957
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_447
timestamp 1688980957
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 1688980957
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_461
timestamp 1688980957
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_473
timestamp 1688980957
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_485
timestamp 1688980957
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_497
timestamp 1688980957
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_503
timestamp 1688980957
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_505
timestamp 1688980957
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_517
timestamp 1688980957
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_529
timestamp 1688980957
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_541
timestamp 1688980957
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_553
timestamp 1688980957
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_559
timestamp 1688980957
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_561
timestamp 1688980957
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_573
timestamp 1688980957
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_585
timestamp 1688980957
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_597
timestamp 1688980957
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_609
timestamp 1688980957
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_615
timestamp 1688980957
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_617
timestamp 1688980957
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_629
timestamp 1688980957
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_641
timestamp 1688980957
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_653
timestamp 1688980957
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_665
timestamp 1688980957
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_671
timestamp 1688980957
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_673
timestamp 1688980957
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_685
timestamp 1688980957
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_697
timestamp 1688980957
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_709
timestamp 1688980957
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_721
timestamp 1688980957
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_727
timestamp 1688980957
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_729
timestamp 1688980957
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 1688980957
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1688980957
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_401
timestamp 1688980957
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_413
timestamp 1688980957
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 1688980957
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1688980957
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 1688980957
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 1688980957
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_457
timestamp 1688980957
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_469
timestamp 1688980957
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_475
timestamp 1688980957
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_477
timestamp 1688980957
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_489
timestamp 1688980957
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_501
timestamp 1688980957
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_513
timestamp 1688980957
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_525
timestamp 1688980957
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_531
timestamp 1688980957
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_533
timestamp 1688980957
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_545
timestamp 1688980957
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_557
timestamp 1688980957
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_569
timestamp 1688980957
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_581
timestamp 1688980957
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_587
timestamp 1688980957
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_589
timestamp 1688980957
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_601
timestamp 1688980957
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_613
timestamp 1688980957
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_625
timestamp 1688980957
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_637
timestamp 1688980957
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_643
timestamp 1688980957
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_645
timestamp 1688980957
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_657
timestamp 1688980957
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_669
timestamp 1688980957
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_681
timestamp 1688980957
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_693
timestamp 1688980957
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_699
timestamp 1688980957
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_701
timestamp 1688980957
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_713
timestamp 1688980957
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_725
timestamp 1688980957
transform 1 0 67804 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_6
timestamp 1688980957
transform 1 0 1656 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_18
timestamp 1688980957
transform 1 0 2760 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_30
timestamp 1688980957
transform 1 0 3864 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_42
timestamp 1688980957
transform 1 0 4968 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_54
timestamp 1688980957
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1688980957
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 1688980957
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1688980957
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1688980957
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1688980957
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 1688980957
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_441
timestamp 1688980957
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_447
timestamp 1688980957
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 1688980957
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_461
timestamp 1688980957
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_473
timestamp 1688980957
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_485
timestamp 1688980957
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_497
timestamp 1688980957
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_503
timestamp 1688980957
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_505
timestamp 1688980957
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_517
timestamp 1688980957
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_529
timestamp 1688980957
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_541
timestamp 1688980957
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_553
timestamp 1688980957
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_559
timestamp 1688980957
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_561
timestamp 1688980957
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_573
timestamp 1688980957
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_585
timestamp 1688980957
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_597
timestamp 1688980957
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_609
timestamp 1688980957
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_615
timestamp 1688980957
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_617
timestamp 1688980957
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_629
timestamp 1688980957
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_641
timestamp 1688980957
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_653
timestamp 1688980957
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_665
timestamp 1688980957
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_671
timestamp 1688980957
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_673
timestamp 1688980957
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_685
timestamp 1688980957
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_697
timestamp 1688980957
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_709
timestamp 1688980957
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_721
timestamp 1688980957
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_727
timestamp 1688980957
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_729
timestamp 1688980957
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1688980957
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1688980957
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 1688980957
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 1688980957
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 1688980957
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_421
timestamp 1688980957
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_433
timestamp 1688980957
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_445
timestamp 1688980957
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_457
timestamp 1688980957
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_469
timestamp 1688980957
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_475
timestamp 1688980957
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_477
timestamp 1688980957
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_489
timestamp 1688980957
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_501
timestamp 1688980957
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_513
timestamp 1688980957
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_525
timestamp 1688980957
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_531
timestamp 1688980957
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_533
timestamp 1688980957
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_545
timestamp 1688980957
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_557
timestamp 1688980957
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_569
timestamp 1688980957
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_581
timestamp 1688980957
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_587
timestamp 1688980957
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_589
timestamp 1688980957
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_601
timestamp 1688980957
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_613
timestamp 1688980957
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_625
timestamp 1688980957
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_637
timestamp 1688980957
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_643
timestamp 1688980957
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_645
timestamp 1688980957
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_657
timestamp 1688980957
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_669
timestamp 1688980957
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_681
timestamp 1688980957
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_693
timestamp 1688980957
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_699
timestamp 1688980957
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_701
timestamp 1688980957
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_713
timestamp 1688980957
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_725
timestamp 1688980957
transform 1 0 67804 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1688980957
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1688980957
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1688980957
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1688980957
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1688980957
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_429
timestamp 1688980957
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_441
timestamp 1688980957
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 1688980957
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_449
timestamp 1688980957
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_461
timestamp 1688980957
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_473
timestamp 1688980957
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_485
timestamp 1688980957
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_497
timestamp 1688980957
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_503
timestamp 1688980957
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_505
timestamp 1688980957
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_517
timestamp 1688980957
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_529
timestamp 1688980957
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_541
timestamp 1688980957
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_553
timestamp 1688980957
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_559
timestamp 1688980957
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_561
timestamp 1688980957
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_573
timestamp 1688980957
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_585
timestamp 1688980957
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_597
timestamp 1688980957
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_609
timestamp 1688980957
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_615
timestamp 1688980957
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_617
timestamp 1688980957
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_629
timestamp 1688980957
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_641
timestamp 1688980957
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_653
timestamp 1688980957
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_665
timestamp 1688980957
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_671
timestamp 1688980957
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_673
timestamp 1688980957
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_685
timestamp 1688980957
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_697
timestamp 1688980957
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_709
timestamp 1688980957
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_721
timestamp 1688980957
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_727
timestamp 1688980957
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1688980957
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1688980957
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 1688980957
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1688980957
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1688980957
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_433
timestamp 1688980957
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_445
timestamp 1688980957
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_457
timestamp 1688980957
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_469
timestamp 1688980957
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_475
timestamp 1688980957
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_477
timestamp 1688980957
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_489
timestamp 1688980957
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_501
timestamp 1688980957
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_513
timestamp 1688980957
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_525
timestamp 1688980957
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_531
timestamp 1688980957
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_533
timestamp 1688980957
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_545
timestamp 1688980957
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_557
timestamp 1688980957
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_569
timestamp 1688980957
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_581
timestamp 1688980957
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_587
timestamp 1688980957
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_589
timestamp 1688980957
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_601
timestamp 1688980957
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_613
timestamp 1688980957
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_625
timestamp 1688980957
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_637
timestamp 1688980957
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_643
timestamp 1688980957
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_645
timestamp 1688980957
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_657
timestamp 1688980957
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_669
timestamp 1688980957
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_681
timestamp 1688980957
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_693
timestamp 1688980957
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_699
timestamp 1688980957
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_701
timestamp 1688980957
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_713
timestamp 1688980957
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_725
timestamp 1688980957
transform 1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1688980957
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1688980957
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1688980957
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 1688980957
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 1688980957
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 1688980957
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 1688980957
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_461
timestamp 1688980957
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_473
timestamp 1688980957
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_485
timestamp 1688980957
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_497
timestamp 1688980957
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_503
timestamp 1688980957
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_505
timestamp 1688980957
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_517
timestamp 1688980957
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_529
timestamp 1688980957
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_541
timestamp 1688980957
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_553
timestamp 1688980957
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_559
timestamp 1688980957
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_561
timestamp 1688980957
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_573
timestamp 1688980957
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_585
timestamp 1688980957
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_597
timestamp 1688980957
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_609
timestamp 1688980957
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_615
timestamp 1688980957
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_617
timestamp 1688980957
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_629
timestamp 1688980957
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_641
timestamp 1688980957
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_653
timestamp 1688980957
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_665
timestamp 1688980957
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_671
timestamp 1688980957
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_673
timestamp 1688980957
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_685
timestamp 1688980957
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_697
timestamp 1688980957
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_709
timestamp 1688980957
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_721
timestamp 1688980957
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_727
timestamp 1688980957
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_729
timestamp 1688980957
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_6
timestamp 1688980957
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_18
timestamp 1688980957
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_26
timestamp 1688980957
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1688980957
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 1688980957
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 1688980957
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1688980957
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 1688980957
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 1688980957
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_457
timestamp 1688980957
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_469
timestamp 1688980957
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_475
timestamp 1688980957
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_477
timestamp 1688980957
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_489
timestamp 1688980957
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_501
timestamp 1688980957
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_513
timestamp 1688980957
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_525
timestamp 1688980957
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_531
timestamp 1688980957
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_533
timestamp 1688980957
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_545
timestamp 1688980957
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_557
timestamp 1688980957
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_569
timestamp 1688980957
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_581
timestamp 1688980957
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_587
timestamp 1688980957
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_589
timestamp 1688980957
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_601
timestamp 1688980957
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_613
timestamp 1688980957
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_625
timestamp 1688980957
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_637
timestamp 1688980957
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_643
timestamp 1688980957
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_645
timestamp 1688980957
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_657
timestamp 1688980957
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_669
timestamp 1688980957
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_681
timestamp 1688980957
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_693
timestamp 1688980957
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_699
timestamp 1688980957
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_701
timestamp 1688980957
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_713
timestamp 1688980957
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_725
timestamp 1688980957
transform 1 0 67804 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1688980957
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1688980957
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1688980957
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 1688980957
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 1688980957
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 1688980957
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1688980957
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 1688980957
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_473
timestamp 1688980957
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_485
timestamp 1688980957
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_497
timestamp 1688980957
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_503
timestamp 1688980957
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_505
timestamp 1688980957
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_517
timestamp 1688980957
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_529
timestamp 1688980957
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_541
timestamp 1688980957
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_553
timestamp 1688980957
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_559
timestamp 1688980957
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_561
timestamp 1688980957
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_573
timestamp 1688980957
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_585
timestamp 1688980957
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_597
timestamp 1688980957
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_609
timestamp 1688980957
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_615
timestamp 1688980957
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_617
timestamp 1688980957
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_629
timestamp 1688980957
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_641
timestamp 1688980957
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_653
timestamp 1688980957
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_665
timestamp 1688980957
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_671
timestamp 1688980957
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_673
timestamp 1688980957
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_685
timestamp 1688980957
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_697
timestamp 1688980957
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_709
timestamp 1688980957
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_721
timestamp 1688980957
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_727
timestamp 1688980957
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_729
timestamp 1688980957
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1688980957
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1688980957
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1688980957
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1688980957
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1688980957
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1688980957
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1688980957
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1688980957
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1688980957
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 1688980957
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_445
timestamp 1688980957
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_457
timestamp 1688980957
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_469
timestamp 1688980957
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_475
timestamp 1688980957
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_477
timestamp 1688980957
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_489
timestamp 1688980957
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_501
timestamp 1688980957
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_513
timestamp 1688980957
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_525
timestamp 1688980957
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_531
timestamp 1688980957
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_533
timestamp 1688980957
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_545
timestamp 1688980957
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_557
timestamp 1688980957
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_569
timestamp 1688980957
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_581
timestamp 1688980957
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_587
timestamp 1688980957
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_589
timestamp 1688980957
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_601
timestamp 1688980957
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_613
timestamp 1688980957
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_625
timestamp 1688980957
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_637
timestamp 1688980957
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_643
timestamp 1688980957
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_645
timestamp 1688980957
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_657
timestamp 1688980957
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_669
timestamp 1688980957
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_681
timestamp 1688980957
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_693
timestamp 1688980957
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_699
timestamp 1688980957
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_701
timestamp 1688980957
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_713
timestamp 1688980957
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_725
timestamp 1688980957
transform 1 0 67804 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_729
timestamp 1688980957
transform 1 0 68172 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1688980957
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1688980957
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1688980957
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1688980957
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1688980957
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1688980957
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1688980957
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1688980957
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1688980957
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1688980957
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1688980957
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_429
timestamp 1688980957
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_441
timestamp 1688980957
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_447
timestamp 1688980957
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_449
timestamp 1688980957
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_461
timestamp 1688980957
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_473
timestamp 1688980957
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_485
timestamp 1688980957
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_497
timestamp 1688980957
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_503
timestamp 1688980957
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_505
timestamp 1688980957
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_517
timestamp 1688980957
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_529
timestamp 1688980957
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_541
timestamp 1688980957
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_553
timestamp 1688980957
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_559
timestamp 1688980957
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_561
timestamp 1688980957
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_573
timestamp 1688980957
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_585
timestamp 1688980957
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_597
timestamp 1688980957
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_609
timestamp 1688980957
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_615
timestamp 1688980957
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_617
timestamp 1688980957
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_629
timestamp 1688980957
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_641
timestamp 1688980957
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_653
timestamp 1688980957
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_665
timestamp 1688980957
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_671
timestamp 1688980957
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_673
timestamp 1688980957
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_685
timestamp 1688980957
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_697
timestamp 1688980957
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_709
timestamp 1688980957
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_721
timestamp 1688980957
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_727
timestamp 1688980957
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_729
timestamp 1688980957
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1688980957
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1688980957
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 1688980957
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 1688980957
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1688980957
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 1688980957
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 1688980957
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 1688980957
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1688980957
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1688980957
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 1688980957
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1688980957
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 1688980957
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 1688980957
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 1688980957
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 1688980957
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_445
timestamp 1688980957
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_457
timestamp 1688980957
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_469
timestamp 1688980957
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_475
timestamp 1688980957
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_477
timestamp 1688980957
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_489
timestamp 1688980957
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_501
timestamp 1688980957
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_513
timestamp 1688980957
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_525
timestamp 1688980957
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_531
timestamp 1688980957
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_533
timestamp 1688980957
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_545
timestamp 1688980957
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_557
timestamp 1688980957
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_569
timestamp 1688980957
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_581
timestamp 1688980957
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_587
timestamp 1688980957
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_589
timestamp 1688980957
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_601
timestamp 1688980957
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_613
timestamp 1688980957
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_625
timestamp 1688980957
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_637
timestamp 1688980957
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_643
timestamp 1688980957
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_645
timestamp 1688980957
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_657
timestamp 1688980957
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_669
timestamp 1688980957
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_681
timestamp 1688980957
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_693
timestamp 1688980957
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_699
timestamp 1688980957
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_701
timestamp 1688980957
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_713
timestamp 1688980957
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_725
timestamp 1688980957
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_6
timestamp 1688980957
transform 1 0 1656 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_18
timestamp 1688980957
transform 1 0 2760 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_30
timestamp 1688980957
transform 1 0 3864 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_42
timestamp 1688980957
transform 1 0 4968 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_54
timestamp 1688980957
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1688980957
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 1688980957
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 1688980957
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 1688980957
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_261
timestamp 1688980957
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_273
timestamp 1688980957
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 1688980957
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 1688980957
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 1688980957
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 1688980957
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 1688980957
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 1688980957
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1688980957
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1688980957
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1688980957
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1688980957
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 1688980957
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_429
timestamp 1688980957
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_441
timestamp 1688980957
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_447
timestamp 1688980957
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_449
timestamp 1688980957
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_461
timestamp 1688980957
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_473
timestamp 1688980957
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_485
timestamp 1688980957
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_497
timestamp 1688980957
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_503
timestamp 1688980957
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_505
timestamp 1688980957
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_517
timestamp 1688980957
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_529
timestamp 1688980957
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_541
timestamp 1688980957
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_553
timestamp 1688980957
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_559
timestamp 1688980957
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_561
timestamp 1688980957
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_573
timestamp 1688980957
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_585
timestamp 1688980957
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_597
timestamp 1688980957
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_609
timestamp 1688980957
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_615
timestamp 1688980957
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_617
timestamp 1688980957
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_629
timestamp 1688980957
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_641
timestamp 1688980957
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_653
timestamp 1688980957
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_665
timestamp 1688980957
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_671
timestamp 1688980957
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_673
timestamp 1688980957
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_685
timestamp 1688980957
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_697
timestamp 1688980957
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_709
timestamp 1688980957
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_721
timestamp 1688980957
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_727
timestamp 1688980957
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_729
timestamp 1688980957
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_209
timestamp 1688980957
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_221
timestamp 1688980957
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_233
timestamp 1688980957
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 1688980957
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 1688980957
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 1688980957
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 1688980957
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1688980957
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1688980957
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1688980957
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1688980957
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1688980957
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1688980957
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1688980957
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 1688980957
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 1688980957
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 1688980957
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_433
timestamp 1688980957
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_445
timestamp 1688980957
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_457
timestamp 1688980957
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_469
timestamp 1688980957
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_475
timestamp 1688980957
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_477
timestamp 1688980957
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_489
timestamp 1688980957
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_501
timestamp 1688980957
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_513
timestamp 1688980957
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_525
timestamp 1688980957
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_531
timestamp 1688980957
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_533
timestamp 1688980957
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_545
timestamp 1688980957
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_557
timestamp 1688980957
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_569
timestamp 1688980957
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_581
timestamp 1688980957
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_587
timestamp 1688980957
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_589
timestamp 1688980957
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_601
timestamp 1688980957
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_613
timestamp 1688980957
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_625
timestamp 1688980957
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_637
timestamp 1688980957
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_643
timestamp 1688980957
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_645
timestamp 1688980957
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_657
timestamp 1688980957
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_669
timestamp 1688980957
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_681
timestamp 1688980957
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_693
timestamp 1688980957
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_699
timestamp 1688980957
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_701
timestamp 1688980957
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_713
timestamp 1688980957
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_725
timestamp 1688980957
transform 1 0 67804 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1688980957
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 1688980957
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_237
timestamp 1688980957
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_249
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 1688980957
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 1688980957
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 1688980957
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 1688980957
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 1688980957
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1688980957
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 1688980957
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 1688980957
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 1688980957
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1688980957
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1688980957
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_429
timestamp 1688980957
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_441
timestamp 1688980957
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_447
timestamp 1688980957
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_449
timestamp 1688980957
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_461
timestamp 1688980957
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_473
timestamp 1688980957
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_485
timestamp 1688980957
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_497
timestamp 1688980957
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_503
timestamp 1688980957
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_505
timestamp 1688980957
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_517
timestamp 1688980957
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_529
timestamp 1688980957
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_541
timestamp 1688980957
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_553
timestamp 1688980957
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_559
timestamp 1688980957
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_561
timestamp 1688980957
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_573
timestamp 1688980957
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_585
timestamp 1688980957
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_597
timestamp 1688980957
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_609
timestamp 1688980957
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_615
timestamp 1688980957
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_617
timestamp 1688980957
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_629
timestamp 1688980957
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_641
timestamp 1688980957
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_653
timestamp 1688980957
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_665
timestamp 1688980957
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_671
timestamp 1688980957
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_673
timestamp 1688980957
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_685
timestamp 1688980957
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_697
timestamp 1688980957
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_709
timestamp 1688980957
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_721
timestamp 1688980957
transform 1 0 67436 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_727
timestamp 1688980957
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_729
timestamp 1688980957
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1688980957
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 1688980957
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 1688980957
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 1688980957
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_233
timestamp 1688980957
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_245
timestamp 1688980957
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 1688980957
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 1688980957
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_277
timestamp 1688980957
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 1688980957
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 1688980957
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 1688980957
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 1688980957
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_333
timestamp 1688980957
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 1688980957
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 1688980957
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 1688980957
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1688980957
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1688980957
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1688980957
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1688980957
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 1688980957
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 1688980957
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 1688980957
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_433
timestamp 1688980957
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_445
timestamp 1688980957
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_457
timestamp 1688980957
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_469
timestamp 1688980957
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_475
timestamp 1688980957
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_477
timestamp 1688980957
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_489
timestamp 1688980957
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_501
timestamp 1688980957
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_513
timestamp 1688980957
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_525
timestamp 1688980957
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_531
timestamp 1688980957
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_533
timestamp 1688980957
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_545
timestamp 1688980957
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_557
timestamp 1688980957
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_569
timestamp 1688980957
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_581
timestamp 1688980957
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_587
timestamp 1688980957
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_589
timestamp 1688980957
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_601
timestamp 1688980957
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_613
timestamp 1688980957
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_625
timestamp 1688980957
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_637
timestamp 1688980957
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_643
timestamp 1688980957
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_645
timestamp 1688980957
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_657
timestamp 1688980957
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_669
timestamp 1688980957
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_681
timestamp 1688980957
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_693
timestamp 1688980957
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_699
timestamp 1688980957
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_701
timestamp 1688980957
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_713
timestamp 1688980957
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_725
timestamp 1688980957
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1688980957
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1688980957
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 1688980957
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_205
timestamp 1688980957
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_217
timestamp 1688980957
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 1688980957
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 1688980957
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 1688980957
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 1688980957
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 1688980957
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1688980957
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 1688980957
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 1688980957
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 1688980957
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 1688980957
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 1688980957
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 1688980957
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1688980957
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 1688980957
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 1688980957
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 1688980957
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 1688980957
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 1688980957
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1688980957
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1688980957
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 1688980957
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_429
timestamp 1688980957
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_441
timestamp 1688980957
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_447
timestamp 1688980957
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_449
timestamp 1688980957
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_461
timestamp 1688980957
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_473
timestamp 1688980957
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_485
timestamp 1688980957
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_497
timestamp 1688980957
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_503
timestamp 1688980957
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_505
timestamp 1688980957
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_517
timestamp 1688980957
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_529
timestamp 1688980957
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_541
timestamp 1688980957
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_553
timestamp 1688980957
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_559
timestamp 1688980957
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_561
timestamp 1688980957
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_573
timestamp 1688980957
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_585
timestamp 1688980957
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_597
timestamp 1688980957
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_609
timestamp 1688980957
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_615
timestamp 1688980957
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_617
timestamp 1688980957
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_629
timestamp 1688980957
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_641
timestamp 1688980957
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_653
timestamp 1688980957
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_665
timestamp 1688980957
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_671
timestamp 1688980957
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_673
timestamp 1688980957
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_685
timestamp 1688980957
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_697
timestamp 1688980957
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_709
timestamp 1688980957
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_721
timestamp 1688980957
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_727
timestamp 1688980957
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_729
timestamp 1688980957
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1688980957
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 1688980957
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1688980957
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 1688980957
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 1688980957
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 1688980957
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 1688980957
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 1688980957
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 1688980957
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 1688980957
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 1688980957
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 1688980957
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 1688980957
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1688980957
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1688980957
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1688980957
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1688980957
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 1688980957
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 1688980957
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1688980957
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1688980957
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1688980957
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 1688980957
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 1688980957
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 1688980957
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 1688980957
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_433
timestamp 1688980957
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_445
timestamp 1688980957
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_457
timestamp 1688980957
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_469
timestamp 1688980957
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_475
timestamp 1688980957
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_477
timestamp 1688980957
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_489
timestamp 1688980957
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_501
timestamp 1688980957
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_513
timestamp 1688980957
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_525
timestamp 1688980957
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_531
timestamp 1688980957
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_533
timestamp 1688980957
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_545
timestamp 1688980957
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_557
timestamp 1688980957
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_569
timestamp 1688980957
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_581
timestamp 1688980957
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_587
timestamp 1688980957
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_589
timestamp 1688980957
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_601
timestamp 1688980957
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_613
timestamp 1688980957
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_625
timestamp 1688980957
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_637
timestamp 1688980957
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_643
timestamp 1688980957
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_645
timestamp 1688980957
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_657
timestamp 1688980957
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_669
timestamp 1688980957
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_681
timestamp 1688980957
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_693
timestamp 1688980957
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_699
timestamp 1688980957
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_701
timestamp 1688980957
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_713
timestamp 1688980957
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_725
timestamp 1688980957
transform 1 0 67804 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 1688980957
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 1688980957
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 1688980957
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 1688980957
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 1688980957
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_261
timestamp 1688980957
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 1688980957
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 1688980957
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1688980957
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 1688980957
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 1688980957
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 1688980957
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 1688980957
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 1688980957
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1688980957
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1688980957
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 1688980957
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 1688980957
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 1688980957
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 1688980957
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1688980957
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1688980957
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1688980957
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 1688980957
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_441
timestamp 1688980957
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 1688980957
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_449
timestamp 1688980957
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_461
timestamp 1688980957
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_473
timestamp 1688980957
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_485
timestamp 1688980957
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_497
timestamp 1688980957
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_503
timestamp 1688980957
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_505
timestamp 1688980957
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_517
timestamp 1688980957
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_529
timestamp 1688980957
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_541
timestamp 1688980957
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_553
timestamp 1688980957
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_559
timestamp 1688980957
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_561
timestamp 1688980957
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_573
timestamp 1688980957
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_585
timestamp 1688980957
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_597
timestamp 1688980957
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_609
timestamp 1688980957
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_615
timestamp 1688980957
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_617
timestamp 1688980957
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_629
timestamp 1688980957
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_641
timestamp 1688980957
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_653
timestamp 1688980957
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_665
timestamp 1688980957
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_671
timestamp 1688980957
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_673
timestamp 1688980957
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_685
timestamp 1688980957
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_697
timestamp 1688980957
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_709
timestamp 1688980957
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_721
timestamp 1688980957
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_727
timestamp 1688980957
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_729
timestamp 1688980957
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 1688980957
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1688980957
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 1688980957
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 1688980957
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 1688980957
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 1688980957
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 1688980957
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 1688980957
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 1688980957
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 1688980957
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_301
timestamp 1688980957
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 1688980957
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1688980957
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 1688980957
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 1688980957
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 1688980957
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 1688980957
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 1688980957
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1688980957
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 1688980957
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 1688980957
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 1688980957
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 1688980957
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 1688980957
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 1688980957
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_433
timestamp 1688980957
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_445
timestamp 1688980957
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_457
timestamp 1688980957
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_469
timestamp 1688980957
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_475
timestamp 1688980957
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_477
timestamp 1688980957
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_489
timestamp 1688980957
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_501
timestamp 1688980957
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_513
timestamp 1688980957
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_525
timestamp 1688980957
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_531
timestamp 1688980957
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_533
timestamp 1688980957
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_545
timestamp 1688980957
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_557
timestamp 1688980957
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_569
timestamp 1688980957
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_581
timestamp 1688980957
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_587
timestamp 1688980957
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_589
timestamp 1688980957
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_601
timestamp 1688980957
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_613
timestamp 1688980957
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_625
timestamp 1688980957
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_637
timestamp 1688980957
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_643
timestamp 1688980957
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_645
timestamp 1688980957
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_657
timestamp 1688980957
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_669
timestamp 1688980957
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_681
timestamp 1688980957
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_693
timestamp 1688980957
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_699
timestamp 1688980957
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_701
timestamp 1688980957
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_713
timestamp 1688980957
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_725
timestamp 1688980957
transform 1 0 67804 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_729
timestamp 1688980957
transform 1 0 68172 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1688980957
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_193
timestamp 1688980957
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_205
timestamp 1688980957
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_217
timestamp 1688980957
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1688980957
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 1688980957
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_249
timestamp 1688980957
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_261
timestamp 1688980957
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_273
timestamp 1688980957
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_279
timestamp 1688980957
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 1688980957
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 1688980957
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_305
timestamp 1688980957
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_317
timestamp 1688980957
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_329
timestamp 1688980957
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 1688980957
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_337
timestamp 1688980957
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_349
timestamp 1688980957
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_361
timestamp 1688980957
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_373
timestamp 1688980957
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_385
timestamp 1688980957
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 1688980957
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1688980957
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 1688980957
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 1688980957
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_429
timestamp 1688980957
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_441
timestamp 1688980957
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_447
timestamp 1688980957
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_449
timestamp 1688980957
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_461
timestamp 1688980957
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_473
timestamp 1688980957
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_485
timestamp 1688980957
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_497
timestamp 1688980957
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_503
timestamp 1688980957
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_505
timestamp 1688980957
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_517
timestamp 1688980957
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_529
timestamp 1688980957
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_541
timestamp 1688980957
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_553
timestamp 1688980957
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_559
timestamp 1688980957
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_561
timestamp 1688980957
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_573
timestamp 1688980957
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_585
timestamp 1688980957
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_597
timestamp 1688980957
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_609
timestamp 1688980957
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_615
timestamp 1688980957
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_617
timestamp 1688980957
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_629
timestamp 1688980957
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_641
timestamp 1688980957
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_653
timestamp 1688980957
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_665
timestamp 1688980957
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_671
timestamp 1688980957
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_673
timestamp 1688980957
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_685
timestamp 1688980957
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_697
timestamp 1688980957
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_709
timestamp 1688980957
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_721
timestamp 1688980957
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_727
timestamp 1688980957
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_729
timestamp 1688980957
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1688980957
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1688980957
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1688980957
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 1688980957
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 1688980957
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1688980957
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_197
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_209
timestamp 1688980957
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_221
timestamp 1688980957
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_233
timestamp 1688980957
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_245
timestamp 1688980957
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_251
timestamp 1688980957
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_253
timestamp 1688980957
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_265
timestamp 1688980957
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_277
timestamp 1688980957
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_289
timestamp 1688980957
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_301
timestamp 1688980957
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_307
timestamp 1688980957
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 1688980957
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 1688980957
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 1688980957
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 1688980957
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 1688980957
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 1688980957
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_365
timestamp 1688980957
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_377
timestamp 1688980957
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_389
timestamp 1688980957
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_401
timestamp 1688980957
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_413
timestamp 1688980957
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_419
timestamp 1688980957
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_421
timestamp 1688980957
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_433
timestamp 1688980957
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_445
timestamp 1688980957
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_457
timestamp 1688980957
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_469
timestamp 1688980957
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_475
timestamp 1688980957
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_477
timestamp 1688980957
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_489
timestamp 1688980957
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_501
timestamp 1688980957
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_513
timestamp 1688980957
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_525
timestamp 1688980957
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_531
timestamp 1688980957
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_533
timestamp 1688980957
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_545
timestamp 1688980957
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_557
timestamp 1688980957
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_569
timestamp 1688980957
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_581
timestamp 1688980957
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_587
timestamp 1688980957
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_589
timestamp 1688980957
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_601
timestamp 1688980957
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_613
timestamp 1688980957
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_625
timestamp 1688980957
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_637
timestamp 1688980957
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_643
timestamp 1688980957
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_645
timestamp 1688980957
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_657
timestamp 1688980957
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_669
timestamp 1688980957
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_681
timestamp 1688980957
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_693
timestamp 1688980957
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_699
timestamp 1688980957
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_701
timestamp 1688980957
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_713
timestamp 1688980957
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_725
timestamp 1688980957
transform 1 0 67804 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_6
timestamp 1688980957
transform 1 0 1656 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_18
timestamp 1688980957
transform 1 0 2760 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_30
timestamp 1688980957
transform 1 0 3864 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_42
timestamp 1688980957
transform 1 0 4968 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_54
timestamp 1688980957
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1688980957
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 1688980957
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1688980957
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 1688980957
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_181
timestamp 1688980957
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_193
timestamp 1688980957
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_205
timestamp 1688980957
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 1688980957
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 1688980957
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 1688980957
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 1688980957
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 1688980957
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 1688980957
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 1688980957
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 1688980957
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_293
timestamp 1688980957
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_305
timestamp 1688980957
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_317
timestamp 1688980957
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 1688980957
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 1688980957
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 1688980957
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_349
timestamp 1688980957
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_361
timestamp 1688980957
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_373
timestamp 1688980957
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_385
timestamp 1688980957
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_391
timestamp 1688980957
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 1688980957
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 1688980957
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 1688980957
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_429
timestamp 1688980957
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_441
timestamp 1688980957
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_447
timestamp 1688980957
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_449
timestamp 1688980957
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_461
timestamp 1688980957
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_473
timestamp 1688980957
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_485
timestamp 1688980957
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_497
timestamp 1688980957
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_503
timestamp 1688980957
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_505
timestamp 1688980957
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_517
timestamp 1688980957
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_529
timestamp 1688980957
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_541
timestamp 1688980957
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_553
timestamp 1688980957
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_559
timestamp 1688980957
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_561
timestamp 1688980957
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_573
timestamp 1688980957
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_585
timestamp 1688980957
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_597
timestamp 1688980957
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_609
timestamp 1688980957
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_615
timestamp 1688980957
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_617
timestamp 1688980957
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_629
timestamp 1688980957
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_641
timestamp 1688980957
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_653
timestamp 1688980957
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_665
timestamp 1688980957
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_671
timestamp 1688980957
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_673
timestamp 1688980957
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_685
timestamp 1688980957
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_697
timestamp 1688980957
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_709
timestamp 1688980957
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_721
timestamp 1688980957
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_727
timestamp 1688980957
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_729
timestamp 1688980957
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1688980957
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1688980957
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1688980957
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 1688980957
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1688980957
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1688980957
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1688980957
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1688980957
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 1688980957
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1688980957
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 1688980957
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 1688980957
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 1688980957
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_189
timestamp 1688980957
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 1688980957
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_197
timestamp 1688980957
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_209
timestamp 1688980957
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_221
timestamp 1688980957
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_233
timestamp 1688980957
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_245
timestamp 1688980957
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 1688980957
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_253
timestamp 1688980957
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_265
timestamp 1688980957
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_277
timestamp 1688980957
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_289
timestamp 1688980957
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_301
timestamp 1688980957
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_307
timestamp 1688980957
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 1688980957
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_321
timestamp 1688980957
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_333
timestamp 1688980957
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_345
timestamp 1688980957
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 1688980957
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 1688980957
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 1688980957
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 1688980957
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 1688980957
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 1688980957
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 1688980957
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 1688980957
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_421
timestamp 1688980957
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_433
timestamp 1688980957
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_445
timestamp 1688980957
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_457
timestamp 1688980957
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_469
timestamp 1688980957
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_475
timestamp 1688980957
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_477
timestamp 1688980957
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_489
timestamp 1688980957
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_501
timestamp 1688980957
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_513
timestamp 1688980957
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_525
timestamp 1688980957
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_531
timestamp 1688980957
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_533
timestamp 1688980957
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_545
timestamp 1688980957
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_557
timestamp 1688980957
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_569
timestamp 1688980957
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_581
timestamp 1688980957
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_587
timestamp 1688980957
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_589
timestamp 1688980957
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_601
timestamp 1688980957
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_613
timestamp 1688980957
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_625
timestamp 1688980957
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_637
timestamp 1688980957
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_643
timestamp 1688980957
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_645
timestamp 1688980957
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_657
timestamp 1688980957
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_669
timestamp 1688980957
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_681
timestamp 1688980957
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_693
timestamp 1688980957
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_699
timestamp 1688980957
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_701
timestamp 1688980957
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_713
timestamp 1688980957
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_725
timestamp 1688980957
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1688980957
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1688980957
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1688980957
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1688980957
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1688980957
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 1688980957
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 1688980957
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1688980957
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 1688980957
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 1688980957
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 1688980957
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 1688980957
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 1688980957
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 1688980957
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_181
timestamp 1688980957
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_193
timestamp 1688980957
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_205
timestamp 1688980957
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_217
timestamp 1688980957
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 1688980957
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 1688980957
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 1688980957
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 1688980957
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 1688980957
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 1688980957
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 1688980957
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 1688980957
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 1688980957
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 1688980957
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 1688980957
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 1688980957
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 1688980957
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 1688980957
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 1688980957
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 1688980957
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 1688980957
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 1688980957
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 1688980957
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 1688980957
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 1688980957
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 1688980957
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_429
timestamp 1688980957
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_441
timestamp 1688980957
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_447
timestamp 1688980957
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_449
timestamp 1688980957
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_461
timestamp 1688980957
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_473
timestamp 1688980957
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_485
timestamp 1688980957
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_497
timestamp 1688980957
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_503
timestamp 1688980957
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_505
timestamp 1688980957
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_517
timestamp 1688980957
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_529
timestamp 1688980957
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_541
timestamp 1688980957
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_553
timestamp 1688980957
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_559
timestamp 1688980957
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_561
timestamp 1688980957
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_573
timestamp 1688980957
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_585
timestamp 1688980957
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_597
timestamp 1688980957
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_609
timestamp 1688980957
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_615
timestamp 1688980957
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_617
timestamp 1688980957
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_629
timestamp 1688980957
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_641
timestamp 1688980957
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_653
timestamp 1688980957
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_665
timestamp 1688980957
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_671
timestamp 1688980957
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_673
timestamp 1688980957
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_685
timestamp 1688980957
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_697
timestamp 1688980957
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_709
timestamp 1688980957
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_721
timestamp 1688980957
transform 1 0 67436 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_727
timestamp 1688980957
transform 1 0 67988 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_729
timestamp 1688980957
transform 1 0 68172 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1688980957
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1688980957
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1688980957
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1688980957
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1688980957
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1688980957
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1688980957
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 1688980957
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1688980957
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1688980957
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 1688980957
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 1688980957
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 1688980957
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 1688980957
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 1688980957
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 1688980957
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 1688980957
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 1688980957
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 1688980957
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_189
timestamp 1688980957
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 1688980957
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_197
timestamp 1688980957
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_209
timestamp 1688980957
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_221
timestamp 1688980957
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_233
timestamp 1688980957
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_245
timestamp 1688980957
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_251
timestamp 1688980957
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 1688980957
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 1688980957
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 1688980957
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 1688980957
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 1688980957
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 1688980957
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1688980957
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 1688980957
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_333
timestamp 1688980957
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_345
timestamp 1688980957
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_357
timestamp 1688980957
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_363
timestamp 1688980957
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 1688980957
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 1688980957
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 1688980957
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 1688980957
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 1688980957
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 1688980957
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_421
timestamp 1688980957
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_433
timestamp 1688980957
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_445
timestamp 1688980957
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_457
timestamp 1688980957
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_469
timestamp 1688980957
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_475
timestamp 1688980957
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_477
timestamp 1688980957
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_489
timestamp 1688980957
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_501
timestamp 1688980957
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_513
timestamp 1688980957
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_525
timestamp 1688980957
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_531
timestamp 1688980957
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_533
timestamp 1688980957
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_545
timestamp 1688980957
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_557
timestamp 1688980957
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_569
timestamp 1688980957
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_581
timestamp 1688980957
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_587
timestamp 1688980957
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_589
timestamp 1688980957
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_601
timestamp 1688980957
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_613
timestamp 1688980957
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_625
timestamp 1688980957
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_637
timestamp 1688980957
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_643
timestamp 1688980957
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_645
timestamp 1688980957
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_657
timestamp 1688980957
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_669
timestamp 1688980957
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_681
timestamp 1688980957
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_693
timestamp 1688980957
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_699
timestamp 1688980957
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_701
timestamp 1688980957
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_713
timestamp 1688980957
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_725
timestamp 1688980957
transform 1 0 67804 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1688980957
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1688980957
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 1688980957
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 1688980957
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 1688980957
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 1688980957
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 1688980957
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 1688980957
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_81
timestamp 1688980957
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_93
timestamp 1688980957
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_105
timestamp 1688980957
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_111
timestamp 1688980957
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1688980957
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1688980957
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 1688980957
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 1688980957
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 1688980957
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 1688980957
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 1688980957
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 1688980957
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_193
timestamp 1688980957
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_205
timestamp 1688980957
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_217
timestamp 1688980957
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_223
timestamp 1688980957
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 1688980957
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_237
timestamp 1688980957
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_249
timestamp 1688980957
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_261
timestamp 1688980957
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_273
timestamp 1688980957
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 1688980957
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 1688980957
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 1688980957
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_305
timestamp 1688980957
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_317
timestamp 1688980957
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_329
timestamp 1688980957
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_335
timestamp 1688980957
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 1688980957
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 1688980957
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 1688980957
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 1688980957
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 1688980957
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 1688980957
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 1688980957
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 1688980957
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 1688980957
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_429
timestamp 1688980957
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_441
timestamp 1688980957
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_447
timestamp 1688980957
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_449
timestamp 1688980957
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_461
timestamp 1688980957
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_473
timestamp 1688980957
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_485
timestamp 1688980957
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_497
timestamp 1688980957
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_503
timestamp 1688980957
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_505
timestamp 1688980957
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_517
timestamp 1688980957
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_529
timestamp 1688980957
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_541
timestamp 1688980957
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_553
timestamp 1688980957
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_559
timestamp 1688980957
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_561
timestamp 1688980957
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_573
timestamp 1688980957
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_585
timestamp 1688980957
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_597
timestamp 1688980957
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_609
timestamp 1688980957
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_615
timestamp 1688980957
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_617
timestamp 1688980957
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_629
timestamp 1688980957
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_641
timestamp 1688980957
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_653
timestamp 1688980957
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_665
timestamp 1688980957
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_671
timestamp 1688980957
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_673
timestamp 1688980957
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_685
timestamp 1688980957
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_697
timestamp 1688980957
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_709
timestamp 1688980957
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_721
timestamp 1688980957
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_727
timestamp 1688980957
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_729
timestamp 1688980957
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_6
timestamp 1688980957
transform 1 0 1656 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_18
timestamp 1688980957
transform 1 0 2760 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80_26
timestamp 1688980957
transform 1 0 3496 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1688980957
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1688980957
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 1688980957
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 1688980957
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 1688980957
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 1688980957
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 1688980957
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1688980957
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 1688980957
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 1688980957
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 1688980957
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 1688980957
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_141
timestamp 1688980957
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 1688980957
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_165
timestamp 1688980957
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_177
timestamp 1688980957
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_189
timestamp 1688980957
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_195
timestamp 1688980957
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 1688980957
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 1688980957
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_221
timestamp 1688980957
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_233
timestamp 1688980957
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_245
timestamp 1688980957
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 1688980957
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 1688980957
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_265
timestamp 1688980957
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_277
timestamp 1688980957
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_289
timestamp 1688980957
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_301
timestamp 1688980957
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 1688980957
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 1688980957
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 1688980957
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_333
timestamp 1688980957
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_345
timestamp 1688980957
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_357
timestamp 1688980957
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_363
timestamp 1688980957
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 1688980957
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 1688980957
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_389
timestamp 1688980957
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_401
timestamp 1688980957
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_413
timestamp 1688980957
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_419
timestamp 1688980957
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_421
timestamp 1688980957
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_433
timestamp 1688980957
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_445
timestamp 1688980957
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_457
timestamp 1688980957
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_469
timestamp 1688980957
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_475
timestamp 1688980957
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_477
timestamp 1688980957
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_489
timestamp 1688980957
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_501
timestamp 1688980957
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_513
timestamp 1688980957
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_525
timestamp 1688980957
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_531
timestamp 1688980957
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_533
timestamp 1688980957
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_545
timestamp 1688980957
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_557
timestamp 1688980957
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_569
timestamp 1688980957
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_581
timestamp 1688980957
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_587
timestamp 1688980957
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_589
timestamp 1688980957
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_601
timestamp 1688980957
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_613
timestamp 1688980957
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_625
timestamp 1688980957
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_637
timestamp 1688980957
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_643
timestamp 1688980957
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_645
timestamp 1688980957
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_657
timestamp 1688980957
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_669
timestamp 1688980957
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_681
timestamp 1688980957
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_693
timestamp 1688980957
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_699
timestamp 1688980957
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_701
timestamp 1688980957
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_713
timestamp 1688980957
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_725
timestamp 1688980957
transform 1 0 67804 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_3
timestamp 1688980957
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_15
timestamp 1688980957
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_27
timestamp 1688980957
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_39
timestamp 1688980957
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_51
timestamp 1688980957
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 1688980957
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 1688980957
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 1688980957
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 1688980957
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 1688980957
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 1688980957
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 1688980957
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 1688980957
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 1688980957
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 1688980957
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 1688980957
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 1688980957
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 1688980957
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 1688980957
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_181
timestamp 1688980957
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_193
timestamp 1688980957
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_205
timestamp 1688980957
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_217
timestamp 1688980957
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_223
timestamp 1688980957
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_225
timestamp 1688980957
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_237
timestamp 1688980957
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_249
timestamp 1688980957
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_261
timestamp 1688980957
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_273
timestamp 1688980957
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_279
timestamp 1688980957
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_281
timestamp 1688980957
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_293
timestamp 1688980957
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_305
timestamp 1688980957
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_317
timestamp 1688980957
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_329
timestamp 1688980957
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_335
timestamp 1688980957
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_337
timestamp 1688980957
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_349
timestamp 1688980957
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_361
timestamp 1688980957
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_373
timestamp 1688980957
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_385
timestamp 1688980957
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_391
timestamp 1688980957
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_393
timestamp 1688980957
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_405
timestamp 1688980957
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_417
timestamp 1688980957
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_429
timestamp 1688980957
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_441
timestamp 1688980957
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_447
timestamp 1688980957
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_449
timestamp 1688980957
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_461
timestamp 1688980957
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_473
timestamp 1688980957
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_485
timestamp 1688980957
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_497
timestamp 1688980957
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_503
timestamp 1688980957
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_505
timestamp 1688980957
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_517
timestamp 1688980957
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_529
timestamp 1688980957
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_541
timestamp 1688980957
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_553
timestamp 1688980957
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_559
timestamp 1688980957
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_561
timestamp 1688980957
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_573
timestamp 1688980957
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_585
timestamp 1688980957
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_597
timestamp 1688980957
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_609
timestamp 1688980957
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_615
timestamp 1688980957
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_617
timestamp 1688980957
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_629
timestamp 1688980957
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_641
timestamp 1688980957
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_653
timestamp 1688980957
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_665
timestamp 1688980957
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_671
timestamp 1688980957
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_673
timestamp 1688980957
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_685
timestamp 1688980957
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_697
timestamp 1688980957
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_709
timestamp 1688980957
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_721
timestamp 1688980957
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_727
timestamp 1688980957
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_729
timestamp 1688980957
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 1688980957
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 1688980957
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 1688980957
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 1688980957
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 1688980957
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_53
timestamp 1688980957
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_65
timestamp 1688980957
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_77
timestamp 1688980957
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 1688980957
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_85
timestamp 1688980957
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_97
timestamp 1688980957
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_109
timestamp 1688980957
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_121
timestamp 1688980957
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_133
timestamp 1688980957
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_139
timestamp 1688980957
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 1688980957
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 1688980957
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_165
timestamp 1688980957
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_177
timestamp 1688980957
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_189
timestamp 1688980957
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_195
timestamp 1688980957
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_197
timestamp 1688980957
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_209
timestamp 1688980957
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_221
timestamp 1688980957
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_233
timestamp 1688980957
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_245
timestamp 1688980957
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_251
timestamp 1688980957
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_253
timestamp 1688980957
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_265
timestamp 1688980957
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_277
timestamp 1688980957
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_289
timestamp 1688980957
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_301
timestamp 1688980957
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_307
timestamp 1688980957
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_309
timestamp 1688980957
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_321
timestamp 1688980957
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_333
timestamp 1688980957
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_345
timestamp 1688980957
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_357
timestamp 1688980957
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_363
timestamp 1688980957
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_365
timestamp 1688980957
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_377
timestamp 1688980957
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_389
timestamp 1688980957
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_401
timestamp 1688980957
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_413
timestamp 1688980957
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_419
timestamp 1688980957
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_421
timestamp 1688980957
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_433
timestamp 1688980957
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_445
timestamp 1688980957
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_457
timestamp 1688980957
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_469
timestamp 1688980957
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_475
timestamp 1688980957
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_477
timestamp 1688980957
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_489
timestamp 1688980957
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_501
timestamp 1688980957
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_513
timestamp 1688980957
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_525
timestamp 1688980957
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_531
timestamp 1688980957
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_533
timestamp 1688980957
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_545
timestamp 1688980957
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_557
timestamp 1688980957
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_569
timestamp 1688980957
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_581
timestamp 1688980957
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_587
timestamp 1688980957
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_589
timestamp 1688980957
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_601
timestamp 1688980957
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_613
timestamp 1688980957
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_625
timestamp 1688980957
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_637
timestamp 1688980957
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_643
timestamp 1688980957
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_645
timestamp 1688980957
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_657
timestamp 1688980957
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_669
timestamp 1688980957
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_681
timestamp 1688980957
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_693
timestamp 1688980957
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_699
timestamp 1688980957
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_701
timestamp 1688980957
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_713
timestamp 1688980957
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82_725
timestamp 1688980957
transform 1 0 67804 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_729
timestamp 1688980957
transform 1 0 68172 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_3
timestamp 1688980957
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_15
timestamp 1688980957
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_27
timestamp 1688980957
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_39
timestamp 1688980957
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_51
timestamp 1688980957
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_55
timestamp 1688980957
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_57
timestamp 1688980957
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_69
timestamp 1688980957
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_81
timestamp 1688980957
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_93
timestamp 1688980957
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_105
timestamp 1688980957
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_111
timestamp 1688980957
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_113
timestamp 1688980957
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_125
timestamp 1688980957
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_137
timestamp 1688980957
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_149
timestamp 1688980957
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_161
timestamp 1688980957
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_167
timestamp 1688980957
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_169
timestamp 1688980957
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_181
timestamp 1688980957
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_193
timestamp 1688980957
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_205
timestamp 1688980957
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_217
timestamp 1688980957
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_223
timestamp 1688980957
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_225
timestamp 1688980957
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_237
timestamp 1688980957
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_249
timestamp 1688980957
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_261
timestamp 1688980957
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_273
timestamp 1688980957
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_279
timestamp 1688980957
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_281
timestamp 1688980957
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_293
timestamp 1688980957
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_305
timestamp 1688980957
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_317
timestamp 1688980957
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_329
timestamp 1688980957
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_335
timestamp 1688980957
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_337
timestamp 1688980957
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_349
timestamp 1688980957
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_361
timestamp 1688980957
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_373
timestamp 1688980957
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_385
timestamp 1688980957
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_391
timestamp 1688980957
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_393
timestamp 1688980957
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_405
timestamp 1688980957
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_417
timestamp 1688980957
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_429
timestamp 1688980957
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_441
timestamp 1688980957
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_447
timestamp 1688980957
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_449
timestamp 1688980957
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_461
timestamp 1688980957
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_473
timestamp 1688980957
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_485
timestamp 1688980957
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_497
timestamp 1688980957
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_503
timestamp 1688980957
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_505
timestamp 1688980957
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_517
timestamp 1688980957
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_529
timestamp 1688980957
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_541
timestamp 1688980957
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_553
timestamp 1688980957
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_559
timestamp 1688980957
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_561
timestamp 1688980957
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_573
timestamp 1688980957
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_585
timestamp 1688980957
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_597
timestamp 1688980957
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_609
timestamp 1688980957
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_615
timestamp 1688980957
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_617
timestamp 1688980957
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_629
timestamp 1688980957
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_641
timestamp 1688980957
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_653
timestamp 1688980957
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_665
timestamp 1688980957
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_671
timestamp 1688980957
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_673
timestamp 1688980957
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_685
timestamp 1688980957
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_697
timestamp 1688980957
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_709
timestamp 1688980957
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_721
timestamp 1688980957
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_727
timestamp 1688980957
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_729
timestamp 1688980957
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_3
timestamp 1688980957
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_15
timestamp 1688980957
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 1688980957
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_29
timestamp 1688980957
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_41
timestamp 1688980957
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_53
timestamp 1688980957
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_65
timestamp 1688980957
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 1688980957
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 1688980957
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_85
timestamp 1688980957
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_97
timestamp 1688980957
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_109
timestamp 1688980957
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_121
timestamp 1688980957
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_133
timestamp 1688980957
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_139
timestamp 1688980957
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_141
timestamp 1688980957
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_153
timestamp 1688980957
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_165
timestamp 1688980957
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_177
timestamp 1688980957
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_189
timestamp 1688980957
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_195
timestamp 1688980957
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_197
timestamp 1688980957
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_209
timestamp 1688980957
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_221
timestamp 1688980957
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_233
timestamp 1688980957
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_245
timestamp 1688980957
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_251
timestamp 1688980957
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_253
timestamp 1688980957
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_265
timestamp 1688980957
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_277
timestamp 1688980957
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_289
timestamp 1688980957
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_301
timestamp 1688980957
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_307
timestamp 1688980957
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_309
timestamp 1688980957
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_321
timestamp 1688980957
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_333
timestamp 1688980957
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_345
timestamp 1688980957
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_357
timestamp 1688980957
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_363
timestamp 1688980957
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_365
timestamp 1688980957
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_377
timestamp 1688980957
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_389
timestamp 1688980957
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_401
timestamp 1688980957
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_413
timestamp 1688980957
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_419
timestamp 1688980957
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_421
timestamp 1688980957
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_433
timestamp 1688980957
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_445
timestamp 1688980957
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_457
timestamp 1688980957
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_469
timestamp 1688980957
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_475
timestamp 1688980957
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_477
timestamp 1688980957
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_489
timestamp 1688980957
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_501
timestamp 1688980957
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_513
timestamp 1688980957
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_525
timestamp 1688980957
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_531
timestamp 1688980957
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_533
timestamp 1688980957
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_545
timestamp 1688980957
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_557
timestamp 1688980957
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_569
timestamp 1688980957
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_581
timestamp 1688980957
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_587
timestamp 1688980957
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_589
timestamp 1688980957
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_601
timestamp 1688980957
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_613
timestamp 1688980957
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_625
timestamp 1688980957
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_637
timestamp 1688980957
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_643
timestamp 1688980957
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_645
timestamp 1688980957
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_657
timestamp 1688980957
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_669
timestamp 1688980957
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_681
timestamp 1688980957
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_693
timestamp 1688980957
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_699
timestamp 1688980957
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_701
timestamp 1688980957
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_713
timestamp 1688980957
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_725
timestamp 1688980957
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_6
timestamp 1688980957
transform 1 0 1656 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_18
timestamp 1688980957
transform 1 0 2760 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_30
timestamp 1688980957
transform 1 0 3864 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_42
timestamp 1688980957
transform 1 0 4968 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85_54
timestamp 1688980957
transform 1 0 6072 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_57
timestamp 1688980957
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 1688980957
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 1688980957
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_93
timestamp 1688980957
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_105
timestamp 1688980957
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_111
timestamp 1688980957
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_113
timestamp 1688980957
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_125
timestamp 1688980957
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_137
timestamp 1688980957
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_149
timestamp 1688980957
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_161
timestamp 1688980957
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_167
timestamp 1688980957
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_169
timestamp 1688980957
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_181
timestamp 1688980957
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_193
timestamp 1688980957
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_205
timestamp 1688980957
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_217
timestamp 1688980957
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_223
timestamp 1688980957
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_225
timestamp 1688980957
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_237
timestamp 1688980957
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_249
timestamp 1688980957
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_261
timestamp 1688980957
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_273
timestamp 1688980957
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_279
timestamp 1688980957
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_281
timestamp 1688980957
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_293
timestamp 1688980957
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_305
timestamp 1688980957
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_317
timestamp 1688980957
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_329
timestamp 1688980957
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_335
timestamp 1688980957
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_337
timestamp 1688980957
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_349
timestamp 1688980957
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_361
timestamp 1688980957
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_373
timestamp 1688980957
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_385
timestamp 1688980957
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_391
timestamp 1688980957
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_393
timestamp 1688980957
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_405
timestamp 1688980957
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_417
timestamp 1688980957
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_429
timestamp 1688980957
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_441
timestamp 1688980957
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_447
timestamp 1688980957
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_449
timestamp 1688980957
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_461
timestamp 1688980957
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_473
timestamp 1688980957
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_485
timestamp 1688980957
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_497
timestamp 1688980957
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_503
timestamp 1688980957
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_505
timestamp 1688980957
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_517
timestamp 1688980957
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_529
timestamp 1688980957
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_541
timestamp 1688980957
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_553
timestamp 1688980957
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_559
timestamp 1688980957
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_561
timestamp 1688980957
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_573
timestamp 1688980957
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_585
timestamp 1688980957
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_597
timestamp 1688980957
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_609
timestamp 1688980957
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_615
timestamp 1688980957
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_617
timestamp 1688980957
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_629
timestamp 1688980957
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_641
timestamp 1688980957
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_653
timestamp 1688980957
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_665
timestamp 1688980957
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_671
timestamp 1688980957
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_673
timestamp 1688980957
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_685
timestamp 1688980957
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_697
timestamp 1688980957
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_709
timestamp 1688980957
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_721
timestamp 1688980957
transform 1 0 67436 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_727
timestamp 1688980957
transform 1 0 67988 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_729
timestamp 1688980957
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_3
timestamp 1688980957
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_15
timestamp 1688980957
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 1688980957
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 1688980957
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 1688980957
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_53
timestamp 1688980957
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_65
timestamp 1688980957
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_77
timestamp 1688980957
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_83
timestamp 1688980957
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_85
timestamp 1688980957
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_97
timestamp 1688980957
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_109
timestamp 1688980957
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_121
timestamp 1688980957
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_133
timestamp 1688980957
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_139
timestamp 1688980957
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_141
timestamp 1688980957
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_153
timestamp 1688980957
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_165
timestamp 1688980957
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_177
timestamp 1688980957
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_189
timestamp 1688980957
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_195
timestamp 1688980957
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_197
timestamp 1688980957
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_209
timestamp 1688980957
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_221
timestamp 1688980957
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_233
timestamp 1688980957
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_245
timestamp 1688980957
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_251
timestamp 1688980957
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_253
timestamp 1688980957
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_265
timestamp 1688980957
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_277
timestamp 1688980957
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_289
timestamp 1688980957
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_301
timestamp 1688980957
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_307
timestamp 1688980957
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_309
timestamp 1688980957
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_321
timestamp 1688980957
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_333
timestamp 1688980957
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_345
timestamp 1688980957
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_357
timestamp 1688980957
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_363
timestamp 1688980957
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_365
timestamp 1688980957
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_377
timestamp 1688980957
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_389
timestamp 1688980957
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_401
timestamp 1688980957
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_413
timestamp 1688980957
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_419
timestamp 1688980957
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_421
timestamp 1688980957
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_433
timestamp 1688980957
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_445
timestamp 1688980957
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_457
timestamp 1688980957
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_469
timestamp 1688980957
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_475
timestamp 1688980957
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_477
timestamp 1688980957
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_489
timestamp 1688980957
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_501
timestamp 1688980957
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_513
timestamp 1688980957
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_525
timestamp 1688980957
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_531
timestamp 1688980957
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_533
timestamp 1688980957
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_545
timestamp 1688980957
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_557
timestamp 1688980957
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_569
timestamp 1688980957
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_581
timestamp 1688980957
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_587
timestamp 1688980957
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_589
timestamp 1688980957
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_601
timestamp 1688980957
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_613
timestamp 1688980957
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_625
timestamp 1688980957
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_637
timestamp 1688980957
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_643
timestamp 1688980957
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_645
timestamp 1688980957
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_657
timestamp 1688980957
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_669
timestamp 1688980957
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_681
timestamp 1688980957
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_693
timestamp 1688980957
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_699
timestamp 1688980957
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_701
timestamp 1688980957
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_713
timestamp 1688980957
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_725
timestamp 1688980957
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_3
timestamp 1688980957
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_15
timestamp 1688980957
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_27
timestamp 1688980957
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_39
timestamp 1688980957
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_51
timestamp 1688980957
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_55
timestamp 1688980957
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_57
timestamp 1688980957
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_69
timestamp 1688980957
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_81
timestamp 1688980957
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_93
timestamp 1688980957
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_105
timestamp 1688980957
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_111
timestamp 1688980957
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_113
timestamp 1688980957
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_125
timestamp 1688980957
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_137
timestamp 1688980957
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_149
timestamp 1688980957
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_161
timestamp 1688980957
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_167
timestamp 1688980957
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_169
timestamp 1688980957
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_181
timestamp 1688980957
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_193
timestamp 1688980957
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_205
timestamp 1688980957
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_217
timestamp 1688980957
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_223
timestamp 1688980957
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_225
timestamp 1688980957
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_237
timestamp 1688980957
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_249
timestamp 1688980957
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_261
timestamp 1688980957
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_273
timestamp 1688980957
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_279
timestamp 1688980957
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_281
timestamp 1688980957
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_293
timestamp 1688980957
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_305
timestamp 1688980957
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_317
timestamp 1688980957
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_329
timestamp 1688980957
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_335
timestamp 1688980957
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_337
timestamp 1688980957
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_349
timestamp 1688980957
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_361
timestamp 1688980957
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_373
timestamp 1688980957
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_385
timestamp 1688980957
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_391
timestamp 1688980957
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_393
timestamp 1688980957
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_405
timestamp 1688980957
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_417
timestamp 1688980957
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_429
timestamp 1688980957
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_441
timestamp 1688980957
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_447
timestamp 1688980957
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_449
timestamp 1688980957
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_461
timestamp 1688980957
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_473
timestamp 1688980957
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_485
timestamp 1688980957
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_497
timestamp 1688980957
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_503
timestamp 1688980957
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_505
timestamp 1688980957
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_517
timestamp 1688980957
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_529
timestamp 1688980957
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_541
timestamp 1688980957
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_553
timestamp 1688980957
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_559
timestamp 1688980957
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_561
timestamp 1688980957
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_573
timestamp 1688980957
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_585
timestamp 1688980957
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_597
timestamp 1688980957
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_609
timestamp 1688980957
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_615
timestamp 1688980957
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_617
timestamp 1688980957
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_629
timestamp 1688980957
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_641
timestamp 1688980957
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_653
timestamp 1688980957
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_665
timestamp 1688980957
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_671
timestamp 1688980957
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_673
timestamp 1688980957
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_685
timestamp 1688980957
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_697
timestamp 1688980957
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_709
timestamp 1688980957
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_721
timestamp 1688980957
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_727
timestamp 1688980957
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_729
timestamp 1688980957
transform 1 0 68172 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_3
timestamp 1688980957
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_15
timestamp 1688980957
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 1688980957
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 1688980957
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 1688980957
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_53
timestamp 1688980957
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_65
timestamp 1688980957
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_77
timestamp 1688980957
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 1688980957
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_85
timestamp 1688980957
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_97
timestamp 1688980957
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_109
timestamp 1688980957
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_121
timestamp 1688980957
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_133
timestamp 1688980957
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_139
timestamp 1688980957
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_141
timestamp 1688980957
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_153
timestamp 1688980957
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_165
timestamp 1688980957
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_177
timestamp 1688980957
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_189
timestamp 1688980957
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_195
timestamp 1688980957
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_197
timestamp 1688980957
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_209
timestamp 1688980957
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_221
timestamp 1688980957
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_233
timestamp 1688980957
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_245
timestamp 1688980957
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_251
timestamp 1688980957
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_253
timestamp 1688980957
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_265
timestamp 1688980957
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_277
timestamp 1688980957
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_289
timestamp 1688980957
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_301
timestamp 1688980957
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_307
timestamp 1688980957
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_309
timestamp 1688980957
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_321
timestamp 1688980957
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_333
timestamp 1688980957
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_345
timestamp 1688980957
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_357
timestamp 1688980957
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_363
timestamp 1688980957
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_365
timestamp 1688980957
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_377
timestamp 1688980957
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_389
timestamp 1688980957
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_401
timestamp 1688980957
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_413
timestamp 1688980957
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_419
timestamp 1688980957
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_421
timestamp 1688980957
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_433
timestamp 1688980957
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_445
timestamp 1688980957
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_457
timestamp 1688980957
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_469
timestamp 1688980957
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_475
timestamp 1688980957
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_477
timestamp 1688980957
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_489
timestamp 1688980957
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_501
timestamp 1688980957
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_513
timestamp 1688980957
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_525
timestamp 1688980957
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_531
timestamp 1688980957
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_533
timestamp 1688980957
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_545
timestamp 1688980957
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_557
timestamp 1688980957
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_569
timestamp 1688980957
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_581
timestamp 1688980957
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_587
timestamp 1688980957
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_589
timestamp 1688980957
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_601
timestamp 1688980957
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_613
timestamp 1688980957
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_625
timestamp 1688980957
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_637
timestamp 1688980957
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_643
timestamp 1688980957
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_645
timestamp 1688980957
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_657
timestamp 1688980957
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_669
timestamp 1688980957
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_681
timestamp 1688980957
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_693
timestamp 1688980957
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_699
timestamp 1688980957
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_701
timestamp 1688980957
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_713
timestamp 1688980957
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_725
timestamp 1688980957
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_3
timestamp 1688980957
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_15
timestamp 1688980957
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_27
timestamp 1688980957
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_39
timestamp 1688980957
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_51
timestamp 1688980957
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 1688980957
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_57
timestamp 1688980957
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_69
timestamp 1688980957
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_81
timestamp 1688980957
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_93
timestamp 1688980957
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_105
timestamp 1688980957
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_111
timestamp 1688980957
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_113
timestamp 1688980957
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_125
timestamp 1688980957
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_137
timestamp 1688980957
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_149
timestamp 1688980957
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_161
timestamp 1688980957
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_167
timestamp 1688980957
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_169
timestamp 1688980957
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_181
timestamp 1688980957
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_193
timestamp 1688980957
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_205
timestamp 1688980957
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_217
timestamp 1688980957
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_223
timestamp 1688980957
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_225
timestamp 1688980957
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_237
timestamp 1688980957
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_249
timestamp 1688980957
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_261
timestamp 1688980957
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_273
timestamp 1688980957
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_279
timestamp 1688980957
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_281
timestamp 1688980957
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_293
timestamp 1688980957
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_305
timestamp 1688980957
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_317
timestamp 1688980957
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_329
timestamp 1688980957
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_335
timestamp 1688980957
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_337
timestamp 1688980957
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_349
timestamp 1688980957
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_361
timestamp 1688980957
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_373
timestamp 1688980957
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_385
timestamp 1688980957
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_391
timestamp 1688980957
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_393
timestamp 1688980957
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_405
timestamp 1688980957
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_417
timestamp 1688980957
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_429
timestamp 1688980957
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_441
timestamp 1688980957
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_447
timestamp 1688980957
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_449
timestamp 1688980957
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_461
timestamp 1688980957
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_473
timestamp 1688980957
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_485
timestamp 1688980957
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_497
timestamp 1688980957
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_503
timestamp 1688980957
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_505
timestamp 1688980957
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_517
timestamp 1688980957
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_529
timestamp 1688980957
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_541
timestamp 1688980957
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_553
timestamp 1688980957
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_559
timestamp 1688980957
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_561
timestamp 1688980957
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_573
timestamp 1688980957
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_585
timestamp 1688980957
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_597
timestamp 1688980957
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_609
timestamp 1688980957
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_615
timestamp 1688980957
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_617
timestamp 1688980957
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_629
timestamp 1688980957
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_641
timestamp 1688980957
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_653
timestamp 1688980957
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_665
timestamp 1688980957
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_671
timestamp 1688980957
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_673
timestamp 1688980957
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_685
timestamp 1688980957
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_697
timestamp 1688980957
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_709
timestamp 1688980957
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_721
timestamp 1688980957
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_727
timestamp 1688980957
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_729
timestamp 1688980957
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_6
timestamp 1688980957
transform 1 0 1656 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_18
timestamp 1688980957
transform 1 0 2760 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90_26
timestamp 1688980957
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 1688980957
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 1688980957
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 1688980957
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 1688980957
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 1688980957
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 1688980957
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_85
timestamp 1688980957
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_97
timestamp 1688980957
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_109
timestamp 1688980957
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_121
timestamp 1688980957
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_133
timestamp 1688980957
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_139
timestamp 1688980957
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_141
timestamp 1688980957
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_153
timestamp 1688980957
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_165
timestamp 1688980957
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_177
timestamp 1688980957
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_189
timestamp 1688980957
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_195
timestamp 1688980957
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_197
timestamp 1688980957
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_209
timestamp 1688980957
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_221
timestamp 1688980957
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_233
timestamp 1688980957
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_245
timestamp 1688980957
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_251
timestamp 1688980957
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_253
timestamp 1688980957
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_265
timestamp 1688980957
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_277
timestamp 1688980957
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_289
timestamp 1688980957
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_301
timestamp 1688980957
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_307
timestamp 1688980957
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_309
timestamp 1688980957
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_321
timestamp 1688980957
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_333
timestamp 1688980957
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_345
timestamp 1688980957
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_357
timestamp 1688980957
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_363
timestamp 1688980957
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_365
timestamp 1688980957
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_377
timestamp 1688980957
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_389
timestamp 1688980957
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_401
timestamp 1688980957
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_413
timestamp 1688980957
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_419
timestamp 1688980957
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_421
timestamp 1688980957
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_433
timestamp 1688980957
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_445
timestamp 1688980957
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_457
timestamp 1688980957
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_469
timestamp 1688980957
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_475
timestamp 1688980957
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_477
timestamp 1688980957
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_489
timestamp 1688980957
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_501
timestamp 1688980957
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_513
timestamp 1688980957
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_525
timestamp 1688980957
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_531
timestamp 1688980957
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_533
timestamp 1688980957
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_545
timestamp 1688980957
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_557
timestamp 1688980957
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_569
timestamp 1688980957
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_581
timestamp 1688980957
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_587
timestamp 1688980957
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_589
timestamp 1688980957
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_601
timestamp 1688980957
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_613
timestamp 1688980957
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_625
timestamp 1688980957
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_637
timestamp 1688980957
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_643
timestamp 1688980957
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_645
timestamp 1688980957
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_657
timestamp 1688980957
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_669
timestamp 1688980957
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_681
timestamp 1688980957
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_693
timestamp 1688980957
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_699
timestamp 1688980957
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_701
timestamp 1688980957
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_713
timestamp 1688980957
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_725
timestamp 1688980957
transform 1 0 67804 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 1688980957
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 1688980957
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_27
timestamp 1688980957
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_39
timestamp 1688980957
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_51
timestamp 1688980957
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_55
timestamp 1688980957
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_57
timestamp 1688980957
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_69
timestamp 1688980957
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_81
timestamp 1688980957
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_93
timestamp 1688980957
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_105
timestamp 1688980957
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_111
timestamp 1688980957
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_113
timestamp 1688980957
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_125
timestamp 1688980957
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_137
timestamp 1688980957
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_149
timestamp 1688980957
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_161
timestamp 1688980957
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_167
timestamp 1688980957
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_169
timestamp 1688980957
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_181
timestamp 1688980957
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_193
timestamp 1688980957
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_205
timestamp 1688980957
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_217
timestamp 1688980957
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_223
timestamp 1688980957
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_225
timestamp 1688980957
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_237
timestamp 1688980957
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_249
timestamp 1688980957
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_261
timestamp 1688980957
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_273
timestamp 1688980957
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_279
timestamp 1688980957
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_281
timestamp 1688980957
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_293
timestamp 1688980957
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_305
timestamp 1688980957
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_317
timestamp 1688980957
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_329
timestamp 1688980957
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_335
timestamp 1688980957
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_337
timestamp 1688980957
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_349
timestamp 1688980957
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_361
timestamp 1688980957
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_373
timestamp 1688980957
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_385
timestamp 1688980957
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_391
timestamp 1688980957
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_393
timestamp 1688980957
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_405
timestamp 1688980957
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_417
timestamp 1688980957
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_429
timestamp 1688980957
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_441
timestamp 1688980957
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_447
timestamp 1688980957
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_449
timestamp 1688980957
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_461
timestamp 1688980957
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_473
timestamp 1688980957
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_485
timestamp 1688980957
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_497
timestamp 1688980957
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_503
timestamp 1688980957
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_505
timestamp 1688980957
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_517
timestamp 1688980957
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_529
timestamp 1688980957
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_541
timestamp 1688980957
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_553
timestamp 1688980957
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_559
timestamp 1688980957
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_561
timestamp 1688980957
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_573
timestamp 1688980957
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_585
timestamp 1688980957
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_597
timestamp 1688980957
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_609
timestamp 1688980957
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_615
timestamp 1688980957
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_617
timestamp 1688980957
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_629
timestamp 1688980957
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_641
timestamp 1688980957
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_653
timestamp 1688980957
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_665
timestamp 1688980957
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_671
timestamp 1688980957
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_673
timestamp 1688980957
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_685
timestamp 1688980957
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_697
timestamp 1688980957
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_709
timestamp 1688980957
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_721
timestamp 1688980957
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_727
timestamp 1688980957
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_729
timestamp 1688980957
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_3
timestamp 1688980957
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_15
timestamp 1688980957
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 1688980957
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_29
timestamp 1688980957
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_41
timestamp 1688980957
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_53
timestamp 1688980957
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_65
timestamp 1688980957
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_77
timestamp 1688980957
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_83
timestamp 1688980957
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_85
timestamp 1688980957
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_97
timestamp 1688980957
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_109
timestamp 1688980957
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_121
timestamp 1688980957
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_133
timestamp 1688980957
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_139
timestamp 1688980957
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_141
timestamp 1688980957
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_153
timestamp 1688980957
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_165
timestamp 1688980957
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_177
timestamp 1688980957
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_189
timestamp 1688980957
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_195
timestamp 1688980957
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_197
timestamp 1688980957
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_209
timestamp 1688980957
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_221
timestamp 1688980957
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_233
timestamp 1688980957
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_245
timestamp 1688980957
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_251
timestamp 1688980957
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_253
timestamp 1688980957
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_265
timestamp 1688980957
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_277
timestamp 1688980957
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_289
timestamp 1688980957
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_301
timestamp 1688980957
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_307
timestamp 1688980957
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_309
timestamp 1688980957
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_321
timestamp 1688980957
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_333
timestamp 1688980957
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_345
timestamp 1688980957
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_357
timestamp 1688980957
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_363
timestamp 1688980957
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_365
timestamp 1688980957
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_377
timestamp 1688980957
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_389
timestamp 1688980957
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_401
timestamp 1688980957
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_413
timestamp 1688980957
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_419
timestamp 1688980957
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_421
timestamp 1688980957
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_433
timestamp 1688980957
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_445
timestamp 1688980957
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_457
timestamp 1688980957
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_469
timestamp 1688980957
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_475
timestamp 1688980957
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_477
timestamp 1688980957
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_489
timestamp 1688980957
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_501
timestamp 1688980957
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_513
timestamp 1688980957
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_525
timestamp 1688980957
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_531
timestamp 1688980957
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_533
timestamp 1688980957
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_545
timestamp 1688980957
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_557
timestamp 1688980957
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_569
timestamp 1688980957
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_581
timestamp 1688980957
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_587
timestamp 1688980957
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_589
timestamp 1688980957
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_601
timestamp 1688980957
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_613
timestamp 1688980957
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_625
timestamp 1688980957
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_637
timestamp 1688980957
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_643
timestamp 1688980957
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_645
timestamp 1688980957
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_657
timestamp 1688980957
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_669
timestamp 1688980957
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_681
timestamp 1688980957
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_693
timestamp 1688980957
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_699
timestamp 1688980957
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_701
timestamp 1688980957
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_713
timestamp 1688980957
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92_725
timestamp 1688980957
transform 1 0 67804 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_729
timestamp 1688980957
transform 1 0 68172 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 1688980957
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 1688980957
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_27
timestamp 1688980957
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_39
timestamp 1688980957
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_51
timestamp 1688980957
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_55
timestamp 1688980957
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_57
timestamp 1688980957
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_69
timestamp 1688980957
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_81
timestamp 1688980957
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_93
timestamp 1688980957
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_105
timestamp 1688980957
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_111
timestamp 1688980957
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_113
timestamp 1688980957
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_125
timestamp 1688980957
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_137
timestamp 1688980957
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_149
timestamp 1688980957
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_161
timestamp 1688980957
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_167
timestamp 1688980957
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_169
timestamp 1688980957
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_181
timestamp 1688980957
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_193
timestamp 1688980957
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_205
timestamp 1688980957
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_217
timestamp 1688980957
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_223
timestamp 1688980957
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_225
timestamp 1688980957
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_237
timestamp 1688980957
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_249
timestamp 1688980957
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_261
timestamp 1688980957
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_273
timestamp 1688980957
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_279
timestamp 1688980957
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_281
timestamp 1688980957
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_293
timestamp 1688980957
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_305
timestamp 1688980957
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_317
timestamp 1688980957
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_329
timestamp 1688980957
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_335
timestamp 1688980957
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_337
timestamp 1688980957
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_349
timestamp 1688980957
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_361
timestamp 1688980957
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_373
timestamp 1688980957
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_385
timestamp 1688980957
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_391
timestamp 1688980957
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_393
timestamp 1688980957
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_405
timestamp 1688980957
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_417
timestamp 1688980957
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_429
timestamp 1688980957
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_441
timestamp 1688980957
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_447
timestamp 1688980957
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_449
timestamp 1688980957
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_461
timestamp 1688980957
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_473
timestamp 1688980957
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_485
timestamp 1688980957
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_497
timestamp 1688980957
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_503
timestamp 1688980957
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_505
timestamp 1688980957
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_517
timestamp 1688980957
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_529
timestamp 1688980957
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_541
timestamp 1688980957
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_553
timestamp 1688980957
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_559
timestamp 1688980957
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_561
timestamp 1688980957
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_573
timestamp 1688980957
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_585
timestamp 1688980957
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_597
timestamp 1688980957
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_609
timestamp 1688980957
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_615
timestamp 1688980957
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_617
timestamp 1688980957
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_629
timestamp 1688980957
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_641
timestamp 1688980957
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_653
timestamp 1688980957
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_665
timestamp 1688980957
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_671
timestamp 1688980957
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_673
timestamp 1688980957
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_685
timestamp 1688980957
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_697
timestamp 1688980957
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_709
timestamp 1688980957
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_721
timestamp 1688980957
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_727
timestamp 1688980957
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_729
timestamp 1688980957
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_3
timestamp 1688980957
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_15
timestamp 1688980957
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 1688980957
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_29
timestamp 1688980957
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_41
timestamp 1688980957
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_53
timestamp 1688980957
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_65
timestamp 1688980957
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_77
timestamp 1688980957
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_83
timestamp 1688980957
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_85
timestamp 1688980957
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_97
timestamp 1688980957
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_109
timestamp 1688980957
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_121
timestamp 1688980957
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_133
timestamp 1688980957
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_139
timestamp 1688980957
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_141
timestamp 1688980957
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_153
timestamp 1688980957
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_165
timestamp 1688980957
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_177
timestamp 1688980957
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_189
timestamp 1688980957
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_195
timestamp 1688980957
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_197
timestamp 1688980957
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_209
timestamp 1688980957
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_221
timestamp 1688980957
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_233
timestamp 1688980957
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_245
timestamp 1688980957
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_251
timestamp 1688980957
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_253
timestamp 1688980957
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_265
timestamp 1688980957
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_277
timestamp 1688980957
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_289
timestamp 1688980957
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_301
timestamp 1688980957
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_307
timestamp 1688980957
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_309
timestamp 1688980957
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_321
timestamp 1688980957
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_333
timestamp 1688980957
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_345
timestamp 1688980957
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_357
timestamp 1688980957
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_363
timestamp 1688980957
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_365
timestamp 1688980957
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_377
timestamp 1688980957
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_389
timestamp 1688980957
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_401
timestamp 1688980957
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_413
timestamp 1688980957
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_419
timestamp 1688980957
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_421
timestamp 1688980957
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_433
timestamp 1688980957
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_445
timestamp 1688980957
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_457
timestamp 1688980957
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_469
timestamp 1688980957
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_475
timestamp 1688980957
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_477
timestamp 1688980957
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_489
timestamp 1688980957
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_501
timestamp 1688980957
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_513
timestamp 1688980957
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_525
timestamp 1688980957
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_531
timestamp 1688980957
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_533
timestamp 1688980957
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_545
timestamp 1688980957
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_557
timestamp 1688980957
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_569
timestamp 1688980957
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_581
timestamp 1688980957
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_587
timestamp 1688980957
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_589
timestamp 1688980957
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_601
timestamp 1688980957
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_613
timestamp 1688980957
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_625
timestamp 1688980957
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_637
timestamp 1688980957
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_643
timestamp 1688980957
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_645
timestamp 1688980957
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_657
timestamp 1688980957
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_669
timestamp 1688980957
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_681
timestamp 1688980957
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_693
timestamp 1688980957
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_699
timestamp 1688980957
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_701
timestamp 1688980957
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_713
timestamp 1688980957
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_725
timestamp 1688980957
transform 1 0 67804 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_3
timestamp 1688980957
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_15
timestamp 1688980957
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_27
timestamp 1688980957
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_39
timestamp 1688980957
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_51
timestamp 1688980957
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_55
timestamp 1688980957
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_57
timestamp 1688980957
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_69
timestamp 1688980957
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_81
timestamp 1688980957
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_93
timestamp 1688980957
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_105
timestamp 1688980957
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_111
timestamp 1688980957
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_113
timestamp 1688980957
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_125
timestamp 1688980957
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_137
timestamp 1688980957
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_149
timestamp 1688980957
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_161
timestamp 1688980957
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_167
timestamp 1688980957
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_169
timestamp 1688980957
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_181
timestamp 1688980957
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_193
timestamp 1688980957
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_205
timestamp 1688980957
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_217
timestamp 1688980957
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_223
timestamp 1688980957
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_225
timestamp 1688980957
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_237
timestamp 1688980957
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_249
timestamp 1688980957
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_261
timestamp 1688980957
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_273
timestamp 1688980957
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_279
timestamp 1688980957
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_281
timestamp 1688980957
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_293
timestamp 1688980957
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_305
timestamp 1688980957
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_317
timestamp 1688980957
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_329
timestamp 1688980957
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_335
timestamp 1688980957
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_337
timestamp 1688980957
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_349
timestamp 1688980957
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_361
timestamp 1688980957
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_373
timestamp 1688980957
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_385
timestamp 1688980957
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_391
timestamp 1688980957
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_393
timestamp 1688980957
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_405
timestamp 1688980957
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_417
timestamp 1688980957
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_429
timestamp 1688980957
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_441
timestamp 1688980957
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_447
timestamp 1688980957
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_449
timestamp 1688980957
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_461
timestamp 1688980957
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_473
timestamp 1688980957
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_485
timestamp 1688980957
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_497
timestamp 1688980957
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_503
timestamp 1688980957
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_505
timestamp 1688980957
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_517
timestamp 1688980957
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_529
timestamp 1688980957
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_541
timestamp 1688980957
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_553
timestamp 1688980957
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_559
timestamp 1688980957
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_561
timestamp 1688980957
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_573
timestamp 1688980957
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_585
timestamp 1688980957
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_597
timestamp 1688980957
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_609
timestamp 1688980957
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_615
timestamp 1688980957
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_617
timestamp 1688980957
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_629
timestamp 1688980957
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_641
timestamp 1688980957
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_653
timestamp 1688980957
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_665
timestamp 1688980957
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_671
timestamp 1688980957
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_673
timestamp 1688980957
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_685
timestamp 1688980957
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_697
timestamp 1688980957
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_709
timestamp 1688980957
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_721
timestamp 1688980957
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_727
timestamp 1688980957
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_729
timestamp 1688980957
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 1688980957
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 1688980957
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 1688980957
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_29
timestamp 1688980957
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_41
timestamp 1688980957
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_53
timestamp 1688980957
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_65
timestamp 1688980957
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_77
timestamp 1688980957
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 1688980957
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_85
timestamp 1688980957
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_97
timestamp 1688980957
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_109
timestamp 1688980957
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_121
timestamp 1688980957
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_133
timestamp 1688980957
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_139
timestamp 1688980957
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_141
timestamp 1688980957
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_153
timestamp 1688980957
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_165
timestamp 1688980957
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_177
timestamp 1688980957
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_189
timestamp 1688980957
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_195
timestamp 1688980957
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_197
timestamp 1688980957
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_209
timestamp 1688980957
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_221
timestamp 1688980957
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_233
timestamp 1688980957
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_245
timestamp 1688980957
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_251
timestamp 1688980957
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_253
timestamp 1688980957
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_265
timestamp 1688980957
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_277
timestamp 1688980957
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_289
timestamp 1688980957
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_301
timestamp 1688980957
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_307
timestamp 1688980957
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_309
timestamp 1688980957
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_321
timestamp 1688980957
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_333
timestamp 1688980957
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_345
timestamp 1688980957
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_357
timestamp 1688980957
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_363
timestamp 1688980957
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_365
timestamp 1688980957
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_377
timestamp 1688980957
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_389
timestamp 1688980957
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_401
timestamp 1688980957
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_413
timestamp 1688980957
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_419
timestamp 1688980957
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_421
timestamp 1688980957
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_433
timestamp 1688980957
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_445
timestamp 1688980957
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_457
timestamp 1688980957
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_469
timestamp 1688980957
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_475
timestamp 1688980957
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_477
timestamp 1688980957
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_489
timestamp 1688980957
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_501
timestamp 1688980957
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_513
timestamp 1688980957
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_525
timestamp 1688980957
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_531
timestamp 1688980957
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_533
timestamp 1688980957
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_545
timestamp 1688980957
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_557
timestamp 1688980957
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_569
timestamp 1688980957
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_581
timestamp 1688980957
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_587
timestamp 1688980957
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_589
timestamp 1688980957
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_601
timestamp 1688980957
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_613
timestamp 1688980957
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_625
timestamp 1688980957
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_637
timestamp 1688980957
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_643
timestamp 1688980957
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_645
timestamp 1688980957
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_657
timestamp 1688980957
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_669
timestamp 1688980957
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_681
timestamp 1688980957
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_693
timestamp 1688980957
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_699
timestamp 1688980957
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_701
timestamp 1688980957
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_713
timestamp 1688980957
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_725
timestamp 1688980957
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_3
timestamp 1688980957
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_15
timestamp 1688980957
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_27
timestamp 1688980957
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_39
timestamp 1688980957
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_51
timestamp 1688980957
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_55
timestamp 1688980957
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_57
timestamp 1688980957
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_69
timestamp 1688980957
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_81
timestamp 1688980957
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_93
timestamp 1688980957
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_105
timestamp 1688980957
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_111
timestamp 1688980957
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_113
timestamp 1688980957
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_125
timestamp 1688980957
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_137
timestamp 1688980957
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_149
timestamp 1688980957
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_161
timestamp 1688980957
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_167
timestamp 1688980957
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_169
timestamp 1688980957
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_181
timestamp 1688980957
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_193
timestamp 1688980957
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_205
timestamp 1688980957
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_217
timestamp 1688980957
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_223
timestamp 1688980957
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_225
timestamp 1688980957
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_237
timestamp 1688980957
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_249
timestamp 1688980957
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_261
timestamp 1688980957
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_273
timestamp 1688980957
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_279
timestamp 1688980957
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_281
timestamp 1688980957
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_293
timestamp 1688980957
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_305
timestamp 1688980957
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_317
timestamp 1688980957
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_329
timestamp 1688980957
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_335
timestamp 1688980957
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_337
timestamp 1688980957
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_349
timestamp 1688980957
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_361
timestamp 1688980957
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_373
timestamp 1688980957
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_385
timestamp 1688980957
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_391
timestamp 1688980957
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_393
timestamp 1688980957
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_405
timestamp 1688980957
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_417
timestamp 1688980957
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_429
timestamp 1688980957
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_441
timestamp 1688980957
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_447
timestamp 1688980957
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_449
timestamp 1688980957
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_461
timestamp 1688980957
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_473
timestamp 1688980957
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_485
timestamp 1688980957
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_497
timestamp 1688980957
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_503
timestamp 1688980957
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_505
timestamp 1688980957
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_517
timestamp 1688980957
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_529
timestamp 1688980957
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_541
timestamp 1688980957
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_553
timestamp 1688980957
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_559
timestamp 1688980957
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_561
timestamp 1688980957
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_573
timestamp 1688980957
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_585
timestamp 1688980957
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_597
timestamp 1688980957
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_609
timestamp 1688980957
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_615
timestamp 1688980957
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_617
timestamp 1688980957
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_629
timestamp 1688980957
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_641
timestamp 1688980957
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_653
timestamp 1688980957
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_665
timestamp 1688980957
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_671
timestamp 1688980957
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_673
timestamp 1688980957
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_685
timestamp 1688980957
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_697
timestamp 1688980957
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_709
timestamp 1688980957
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_721
timestamp 1688980957
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_727
timestamp 1688980957
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_729
timestamp 1688980957
transform 1 0 68172 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_3
timestamp 1688980957
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_15
timestamp 1688980957
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 1688980957
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_29
timestamp 1688980957
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_41
timestamp 1688980957
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_53
timestamp 1688980957
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_65
timestamp 1688980957
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_77
timestamp 1688980957
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_83
timestamp 1688980957
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_85
timestamp 1688980957
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_97
timestamp 1688980957
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_109
timestamp 1688980957
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_121
timestamp 1688980957
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_133
timestamp 1688980957
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_139
timestamp 1688980957
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_141
timestamp 1688980957
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_153
timestamp 1688980957
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_165
timestamp 1688980957
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_177
timestamp 1688980957
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_189
timestamp 1688980957
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_195
timestamp 1688980957
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_197
timestamp 1688980957
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_209
timestamp 1688980957
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_221
timestamp 1688980957
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_233
timestamp 1688980957
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_245
timestamp 1688980957
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_251
timestamp 1688980957
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_253
timestamp 1688980957
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_265
timestamp 1688980957
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_277
timestamp 1688980957
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_289
timestamp 1688980957
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_301
timestamp 1688980957
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_307
timestamp 1688980957
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_309
timestamp 1688980957
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_321
timestamp 1688980957
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_333
timestamp 1688980957
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_345
timestamp 1688980957
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_357
timestamp 1688980957
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_363
timestamp 1688980957
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_365
timestamp 1688980957
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_377
timestamp 1688980957
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_389
timestamp 1688980957
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_401
timestamp 1688980957
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_413
timestamp 1688980957
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_419
timestamp 1688980957
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_421
timestamp 1688980957
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_433
timestamp 1688980957
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_445
timestamp 1688980957
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_457
timestamp 1688980957
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_469
timestamp 1688980957
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_475
timestamp 1688980957
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_477
timestamp 1688980957
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_489
timestamp 1688980957
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_501
timestamp 1688980957
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_513
timestamp 1688980957
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_525
timestamp 1688980957
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_531
timestamp 1688980957
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_533
timestamp 1688980957
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_545
timestamp 1688980957
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_557
timestamp 1688980957
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_569
timestamp 1688980957
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_581
timestamp 1688980957
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_587
timestamp 1688980957
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_589
timestamp 1688980957
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_601
timestamp 1688980957
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_613
timestamp 1688980957
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_625
timestamp 1688980957
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_637
timestamp 1688980957
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_643
timestamp 1688980957
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_645
timestamp 1688980957
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_657
timestamp 1688980957
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_669
timestamp 1688980957
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_681
timestamp 1688980957
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_693
timestamp 1688980957
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_699
timestamp 1688980957
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_701
timestamp 1688980957
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_713
timestamp 1688980957
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_725
timestamp 1688980957
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_3
timestamp 1688980957
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_15
timestamp 1688980957
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_27
timestamp 1688980957
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_39
timestamp 1688980957
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_51
timestamp 1688980957
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_55
timestamp 1688980957
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 1688980957
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 1688980957
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 1688980957
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_93
timestamp 1688980957
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_105
timestamp 1688980957
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_111
timestamp 1688980957
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_113
timestamp 1688980957
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_125
timestamp 1688980957
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_137
timestamp 1688980957
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_149
timestamp 1688980957
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_161
timestamp 1688980957
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_167
timestamp 1688980957
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_169
timestamp 1688980957
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_181
timestamp 1688980957
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_193
timestamp 1688980957
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_205
timestamp 1688980957
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_217
timestamp 1688980957
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_223
timestamp 1688980957
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_225
timestamp 1688980957
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_237
timestamp 1688980957
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_249
timestamp 1688980957
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_261
timestamp 1688980957
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_273
timestamp 1688980957
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_279
timestamp 1688980957
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_281
timestamp 1688980957
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_293
timestamp 1688980957
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_305
timestamp 1688980957
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_317
timestamp 1688980957
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_329
timestamp 1688980957
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_335
timestamp 1688980957
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_337
timestamp 1688980957
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_349
timestamp 1688980957
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_361
timestamp 1688980957
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_373
timestamp 1688980957
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_385
timestamp 1688980957
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_391
timestamp 1688980957
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_393
timestamp 1688980957
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_405
timestamp 1688980957
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_417
timestamp 1688980957
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_429
timestamp 1688980957
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_441
timestamp 1688980957
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_447
timestamp 1688980957
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_449
timestamp 1688980957
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_461
timestamp 1688980957
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_473
timestamp 1688980957
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_485
timestamp 1688980957
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_497
timestamp 1688980957
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_503
timestamp 1688980957
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_505
timestamp 1688980957
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_517
timestamp 1688980957
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_529
timestamp 1688980957
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_541
timestamp 1688980957
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_553
timestamp 1688980957
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_559
timestamp 1688980957
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_561
timestamp 1688980957
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_573
timestamp 1688980957
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_585
timestamp 1688980957
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_597
timestamp 1688980957
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_609
timestamp 1688980957
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_615
timestamp 1688980957
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_617
timestamp 1688980957
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_629
timestamp 1688980957
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_641
timestamp 1688980957
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_653
timestamp 1688980957
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_665
timestamp 1688980957
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_671
timestamp 1688980957
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_673
timestamp 1688980957
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_685
timestamp 1688980957
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_697
timestamp 1688980957
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_709
timestamp 1688980957
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_721
timestamp 1688980957
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_727
timestamp 1688980957
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_729
timestamp 1688980957
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_6
timestamp 1688980957
transform 1 0 1656 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_18
timestamp 1688980957
transform 1 0 2760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_26
timestamp 1688980957
transform 1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_29
timestamp 1688980957
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_41
timestamp 1688980957
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_53
timestamp 1688980957
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_65
timestamp 1688980957
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_77
timestamp 1688980957
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_83
timestamp 1688980957
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_85
timestamp 1688980957
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_97
timestamp 1688980957
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_109
timestamp 1688980957
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_121
timestamp 1688980957
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_133
timestamp 1688980957
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_139
timestamp 1688980957
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_141
timestamp 1688980957
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_153
timestamp 1688980957
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_165
timestamp 1688980957
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_177
timestamp 1688980957
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_189
timestamp 1688980957
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_195
timestamp 1688980957
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_197
timestamp 1688980957
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_209
timestamp 1688980957
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_221
timestamp 1688980957
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_233
timestamp 1688980957
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_245
timestamp 1688980957
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_251
timestamp 1688980957
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_253
timestamp 1688980957
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_265
timestamp 1688980957
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_277
timestamp 1688980957
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_289
timestamp 1688980957
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_301
timestamp 1688980957
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_307
timestamp 1688980957
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_309
timestamp 1688980957
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_321
timestamp 1688980957
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_333
timestamp 1688980957
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_345
timestamp 1688980957
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_357
timestamp 1688980957
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_363
timestamp 1688980957
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_365
timestamp 1688980957
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_377
timestamp 1688980957
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_389
timestamp 1688980957
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_401
timestamp 1688980957
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_413
timestamp 1688980957
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_419
timestamp 1688980957
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_421
timestamp 1688980957
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_433
timestamp 1688980957
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_445
timestamp 1688980957
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_457
timestamp 1688980957
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_469
timestamp 1688980957
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_475
timestamp 1688980957
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_477
timestamp 1688980957
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_489
timestamp 1688980957
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_501
timestamp 1688980957
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_513
timestamp 1688980957
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_525
timestamp 1688980957
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_531
timestamp 1688980957
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_533
timestamp 1688980957
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_545
timestamp 1688980957
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_557
timestamp 1688980957
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_569
timestamp 1688980957
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_581
timestamp 1688980957
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_587
timestamp 1688980957
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_589
timestamp 1688980957
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_601
timestamp 1688980957
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_613
timestamp 1688980957
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_625
timestamp 1688980957
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_637
timestamp 1688980957
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_643
timestamp 1688980957
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_645
timestamp 1688980957
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_657
timestamp 1688980957
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_669
timestamp 1688980957
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_681
timestamp 1688980957
transform 1 0 63756 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_693
timestamp 1688980957
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_699
timestamp 1688980957
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_701
timestamp 1688980957
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_713
timestamp 1688980957
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_725
timestamp 1688980957
transform 1 0 67804 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_3
timestamp 1688980957
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_15
timestamp 1688980957
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_27
timestamp 1688980957
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_39
timestamp 1688980957
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_51
timestamp 1688980957
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_55
timestamp 1688980957
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_57
timestamp 1688980957
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_69
timestamp 1688980957
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_81
timestamp 1688980957
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_93
timestamp 1688980957
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_105
timestamp 1688980957
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_111
timestamp 1688980957
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_113
timestamp 1688980957
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_125
timestamp 1688980957
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_137
timestamp 1688980957
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_149
timestamp 1688980957
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_161
timestamp 1688980957
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_167
timestamp 1688980957
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_169
timestamp 1688980957
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_181
timestamp 1688980957
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_193
timestamp 1688980957
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_205
timestamp 1688980957
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_217
timestamp 1688980957
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_223
timestamp 1688980957
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_225
timestamp 1688980957
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_237
timestamp 1688980957
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_249
timestamp 1688980957
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_261
timestamp 1688980957
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_273
timestamp 1688980957
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_279
timestamp 1688980957
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_281
timestamp 1688980957
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_293
timestamp 1688980957
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_305
timestamp 1688980957
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_317
timestamp 1688980957
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_329
timestamp 1688980957
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_335
timestamp 1688980957
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_337
timestamp 1688980957
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_349
timestamp 1688980957
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_361
timestamp 1688980957
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_373
timestamp 1688980957
transform 1 0 35420 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_385
timestamp 1688980957
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_391
timestamp 1688980957
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_393
timestamp 1688980957
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_405
timestamp 1688980957
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_417
timestamp 1688980957
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_429
timestamp 1688980957
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_441
timestamp 1688980957
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_447
timestamp 1688980957
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_449
timestamp 1688980957
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_461
timestamp 1688980957
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_473
timestamp 1688980957
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_485
timestamp 1688980957
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_497
timestamp 1688980957
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_503
timestamp 1688980957
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_505
timestamp 1688980957
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_517
timestamp 1688980957
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_529
timestamp 1688980957
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_541
timestamp 1688980957
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_553
timestamp 1688980957
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_559
timestamp 1688980957
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_561
timestamp 1688980957
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_573
timestamp 1688980957
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_585
timestamp 1688980957
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_597
timestamp 1688980957
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_609
timestamp 1688980957
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_615
timestamp 1688980957
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_617
timestamp 1688980957
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_629
timestamp 1688980957
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_641
timestamp 1688980957
transform 1 0 60076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_653
timestamp 1688980957
transform 1 0 61180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_665
timestamp 1688980957
transform 1 0 62284 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_671
timestamp 1688980957
transform 1 0 62836 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_673
timestamp 1688980957
transform 1 0 63020 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_685
timestamp 1688980957
transform 1 0 64124 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_697
timestamp 1688980957
transform 1 0 65228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_709
timestamp 1688980957
transform 1 0 66332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_721
timestamp 1688980957
transform 1 0 67436 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_727
timestamp 1688980957
transform 1 0 67988 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_729
timestamp 1688980957
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_3
timestamp 1688980957
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_15
timestamp 1688980957
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_27
timestamp 1688980957
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_29
timestamp 1688980957
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_41
timestamp 1688980957
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_53
timestamp 1688980957
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_65
timestamp 1688980957
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_77
timestamp 1688980957
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_83
timestamp 1688980957
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_85
timestamp 1688980957
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_97
timestamp 1688980957
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_109
timestamp 1688980957
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_121
timestamp 1688980957
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_133
timestamp 1688980957
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_139
timestamp 1688980957
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_141
timestamp 1688980957
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_153
timestamp 1688980957
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_165
timestamp 1688980957
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_177
timestamp 1688980957
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_189
timestamp 1688980957
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_195
timestamp 1688980957
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_197
timestamp 1688980957
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_209
timestamp 1688980957
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_221
timestamp 1688980957
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_233
timestamp 1688980957
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_245
timestamp 1688980957
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_251
timestamp 1688980957
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_253
timestamp 1688980957
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_265
timestamp 1688980957
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_277
timestamp 1688980957
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_289
timestamp 1688980957
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_301
timestamp 1688980957
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_307
timestamp 1688980957
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_309
timestamp 1688980957
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_321
timestamp 1688980957
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_333
timestamp 1688980957
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_345
timestamp 1688980957
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_357
timestamp 1688980957
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_363
timestamp 1688980957
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_365
timestamp 1688980957
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_377
timestamp 1688980957
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_389
timestamp 1688980957
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_401
timestamp 1688980957
transform 1 0 37996 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_413
timestamp 1688980957
transform 1 0 39100 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_419
timestamp 1688980957
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_421
timestamp 1688980957
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_433
timestamp 1688980957
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_445
timestamp 1688980957
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_457
timestamp 1688980957
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_469
timestamp 1688980957
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_475
timestamp 1688980957
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_477
timestamp 1688980957
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_489
timestamp 1688980957
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_501
timestamp 1688980957
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_513
timestamp 1688980957
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_525
timestamp 1688980957
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_531
timestamp 1688980957
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_533
timestamp 1688980957
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_545
timestamp 1688980957
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_557
timestamp 1688980957
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_569
timestamp 1688980957
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_581
timestamp 1688980957
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_587
timestamp 1688980957
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_589
timestamp 1688980957
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_601
timestamp 1688980957
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_613
timestamp 1688980957
transform 1 0 57500 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_625
timestamp 1688980957
transform 1 0 58604 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_637
timestamp 1688980957
transform 1 0 59708 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_643
timestamp 1688980957
transform 1 0 60260 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_645
timestamp 1688980957
transform 1 0 60444 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_657
timestamp 1688980957
transform 1 0 61548 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_669
timestamp 1688980957
transform 1 0 62652 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_681
timestamp 1688980957
transform 1 0 63756 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_693
timestamp 1688980957
transform 1 0 64860 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_699
timestamp 1688980957
transform 1 0 65412 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_701
timestamp 1688980957
transform 1 0 65596 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_713
timestamp 1688980957
transform 1 0 66700 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_725
timestamp 1688980957
transform 1 0 67804 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_729
timestamp 1688980957
transform 1 0 68172 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_3
timestamp 1688980957
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_15
timestamp 1688980957
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_27
timestamp 1688980957
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_39
timestamp 1688980957
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_51
timestamp 1688980957
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_55
timestamp 1688980957
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_57
timestamp 1688980957
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_69
timestamp 1688980957
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_81
timestamp 1688980957
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_93
timestamp 1688980957
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_105
timestamp 1688980957
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_111
timestamp 1688980957
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_113
timestamp 1688980957
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_125
timestamp 1688980957
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_137
timestamp 1688980957
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_149
timestamp 1688980957
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_161
timestamp 1688980957
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_167
timestamp 1688980957
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_169
timestamp 1688980957
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_181
timestamp 1688980957
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_193
timestamp 1688980957
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_205
timestamp 1688980957
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_217
timestamp 1688980957
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_223
timestamp 1688980957
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_225
timestamp 1688980957
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_237
timestamp 1688980957
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_249
timestamp 1688980957
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_261
timestamp 1688980957
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_273
timestamp 1688980957
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_279
timestamp 1688980957
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_281
timestamp 1688980957
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_293
timestamp 1688980957
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_305
timestamp 1688980957
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_317
timestamp 1688980957
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_329
timestamp 1688980957
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_335
timestamp 1688980957
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_337
timestamp 1688980957
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_349
timestamp 1688980957
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_361
timestamp 1688980957
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_373
timestamp 1688980957
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_385
timestamp 1688980957
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_391
timestamp 1688980957
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_393
timestamp 1688980957
transform 1 0 37260 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_405
timestamp 1688980957
transform 1 0 38364 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_417
timestamp 1688980957
transform 1 0 39468 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_429
timestamp 1688980957
transform 1 0 40572 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_441
timestamp 1688980957
transform 1 0 41676 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_447
timestamp 1688980957
transform 1 0 42228 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_449
timestamp 1688980957
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_461
timestamp 1688980957
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_473
timestamp 1688980957
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_485
timestamp 1688980957
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_497
timestamp 1688980957
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_503
timestamp 1688980957
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_505
timestamp 1688980957
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_517
timestamp 1688980957
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_529
timestamp 1688980957
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_541
timestamp 1688980957
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_553
timestamp 1688980957
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_559
timestamp 1688980957
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_561
timestamp 1688980957
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_573
timestamp 1688980957
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_585
timestamp 1688980957
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_597
timestamp 1688980957
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_609
timestamp 1688980957
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_615
timestamp 1688980957
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_617
timestamp 1688980957
transform 1 0 57868 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_629
timestamp 1688980957
transform 1 0 58972 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_641
timestamp 1688980957
transform 1 0 60076 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_653
timestamp 1688980957
transform 1 0 61180 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_665
timestamp 1688980957
transform 1 0 62284 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_671
timestamp 1688980957
transform 1 0 62836 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_673
timestamp 1688980957
transform 1 0 63020 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_685
timestamp 1688980957
transform 1 0 64124 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_697
timestamp 1688980957
transform 1 0 65228 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_709
timestamp 1688980957
transform 1 0 66332 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_721
timestamp 1688980957
transform 1 0 67436 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_727
timestamp 1688980957
transform 1 0 67988 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_729
timestamp 1688980957
transform 1 0 68172 0 -1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_3
timestamp 1688980957
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_15
timestamp 1688980957
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_27
timestamp 1688980957
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_29
timestamp 1688980957
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_41
timestamp 1688980957
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_53
timestamp 1688980957
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_65
timestamp 1688980957
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_77
timestamp 1688980957
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_83
timestamp 1688980957
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_85
timestamp 1688980957
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_97
timestamp 1688980957
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_109
timestamp 1688980957
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_121
timestamp 1688980957
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_133
timestamp 1688980957
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_139
timestamp 1688980957
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_141
timestamp 1688980957
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_153
timestamp 1688980957
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_165
timestamp 1688980957
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_177
timestamp 1688980957
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_189
timestamp 1688980957
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_195
timestamp 1688980957
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_197
timestamp 1688980957
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_209
timestamp 1688980957
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_221
timestamp 1688980957
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_233
timestamp 1688980957
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_245
timestamp 1688980957
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_251
timestamp 1688980957
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_253
timestamp 1688980957
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_265
timestamp 1688980957
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_277
timestamp 1688980957
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_289
timestamp 1688980957
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_301
timestamp 1688980957
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_307
timestamp 1688980957
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_309
timestamp 1688980957
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_321
timestamp 1688980957
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_333
timestamp 1688980957
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_345
timestamp 1688980957
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_357
timestamp 1688980957
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_363
timestamp 1688980957
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_365
timestamp 1688980957
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_377
timestamp 1688980957
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_389
timestamp 1688980957
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_401
timestamp 1688980957
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_413
timestamp 1688980957
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_419
timestamp 1688980957
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_421
timestamp 1688980957
transform 1 0 39836 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_433
timestamp 1688980957
transform 1 0 40940 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_445
timestamp 1688980957
transform 1 0 42044 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_457
timestamp 1688980957
transform 1 0 43148 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_469
timestamp 1688980957
transform 1 0 44252 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_475
timestamp 1688980957
transform 1 0 44804 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_477
timestamp 1688980957
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_489
timestamp 1688980957
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_501
timestamp 1688980957
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_513
timestamp 1688980957
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_525
timestamp 1688980957
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_531
timestamp 1688980957
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_533
timestamp 1688980957
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_545
timestamp 1688980957
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_557
timestamp 1688980957
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_569
timestamp 1688980957
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_581
timestamp 1688980957
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_587
timestamp 1688980957
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_589
timestamp 1688980957
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_601
timestamp 1688980957
transform 1 0 56396 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_613
timestamp 1688980957
transform 1 0 57500 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_625
timestamp 1688980957
transform 1 0 58604 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_637
timestamp 1688980957
transform 1 0 59708 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_643
timestamp 1688980957
transform 1 0 60260 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_645
timestamp 1688980957
transform 1 0 60444 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_657
timestamp 1688980957
transform 1 0 61548 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_669
timestamp 1688980957
transform 1 0 62652 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_681
timestamp 1688980957
transform 1 0 63756 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_693
timestamp 1688980957
transform 1 0 64860 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_699
timestamp 1688980957
transform 1 0 65412 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_701
timestamp 1688980957
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_713
timestamp 1688980957
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_725
timestamp 1688980957
transform 1 0 67804 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_6
timestamp 1688980957
transform 1 0 1656 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_18
timestamp 1688980957
transform 1 0 2760 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_30
timestamp 1688980957
transform 1 0 3864 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_42
timestamp 1688980957
transform 1 0 4968 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105_54
timestamp 1688980957
transform 1 0 6072 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_57
timestamp 1688980957
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_69
timestamp 1688980957
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_81
timestamp 1688980957
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_93
timestamp 1688980957
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_105
timestamp 1688980957
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_111
timestamp 1688980957
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_113
timestamp 1688980957
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_125
timestamp 1688980957
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_137
timestamp 1688980957
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_149
timestamp 1688980957
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_161
timestamp 1688980957
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_167
timestamp 1688980957
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_169
timestamp 1688980957
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_181
timestamp 1688980957
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_193
timestamp 1688980957
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_205
timestamp 1688980957
transform 1 0 19964 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_217
timestamp 1688980957
transform 1 0 21068 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_223
timestamp 1688980957
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_225
timestamp 1688980957
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_237
timestamp 1688980957
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_249
timestamp 1688980957
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_261
timestamp 1688980957
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_273
timestamp 1688980957
transform 1 0 26220 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_279
timestamp 1688980957
transform 1 0 26772 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_281
timestamp 1688980957
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_293
timestamp 1688980957
transform 1 0 28060 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_305
timestamp 1688980957
transform 1 0 29164 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_317
timestamp 1688980957
transform 1 0 30268 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_329
timestamp 1688980957
transform 1 0 31372 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_335
timestamp 1688980957
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_337
timestamp 1688980957
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_349
timestamp 1688980957
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_361
timestamp 1688980957
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_373
timestamp 1688980957
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_385
timestamp 1688980957
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_391
timestamp 1688980957
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_393
timestamp 1688980957
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_405
timestamp 1688980957
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_417
timestamp 1688980957
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_429
timestamp 1688980957
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_441
timestamp 1688980957
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_447
timestamp 1688980957
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_449
timestamp 1688980957
transform 1 0 42412 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_461
timestamp 1688980957
transform 1 0 43516 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_473
timestamp 1688980957
transform 1 0 44620 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_485
timestamp 1688980957
transform 1 0 45724 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_497
timestamp 1688980957
transform 1 0 46828 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_503
timestamp 1688980957
transform 1 0 47380 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_505
timestamp 1688980957
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_517
timestamp 1688980957
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_529
timestamp 1688980957
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_541
timestamp 1688980957
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_553
timestamp 1688980957
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_559
timestamp 1688980957
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_561
timestamp 1688980957
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_573
timestamp 1688980957
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_585
timestamp 1688980957
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_597
timestamp 1688980957
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_609
timestamp 1688980957
transform 1 0 57132 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_615
timestamp 1688980957
transform 1 0 57684 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_617
timestamp 1688980957
transform 1 0 57868 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_629
timestamp 1688980957
transform 1 0 58972 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_641
timestamp 1688980957
transform 1 0 60076 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_653
timestamp 1688980957
transform 1 0 61180 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_665
timestamp 1688980957
transform 1 0 62284 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_671
timestamp 1688980957
transform 1 0 62836 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_673
timestamp 1688980957
transform 1 0 63020 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_685
timestamp 1688980957
transform 1 0 64124 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_697
timestamp 1688980957
transform 1 0 65228 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_709
timestamp 1688980957
transform 1 0 66332 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_721
timestamp 1688980957
transform 1 0 67436 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_727
timestamp 1688980957
transform 1 0 67988 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105_729
timestamp 1688980957
transform 1 0 68172 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_3
timestamp 1688980957
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_15
timestamp 1688980957
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_27
timestamp 1688980957
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_29
timestamp 1688980957
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_41
timestamp 1688980957
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_53
timestamp 1688980957
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_65
timestamp 1688980957
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_77
timestamp 1688980957
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_83
timestamp 1688980957
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_85
timestamp 1688980957
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_97
timestamp 1688980957
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_109
timestamp 1688980957
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_121
timestamp 1688980957
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_133
timestamp 1688980957
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_139
timestamp 1688980957
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_141
timestamp 1688980957
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_153
timestamp 1688980957
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_165
timestamp 1688980957
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_177
timestamp 1688980957
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_189
timestamp 1688980957
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_195
timestamp 1688980957
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_197
timestamp 1688980957
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_209
timestamp 1688980957
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_221
timestamp 1688980957
transform 1 0 21436 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_233
timestamp 1688980957
transform 1 0 22540 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_245
timestamp 1688980957
transform 1 0 23644 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_251
timestamp 1688980957
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_253
timestamp 1688980957
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_265
timestamp 1688980957
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_277
timestamp 1688980957
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_289
timestamp 1688980957
transform 1 0 27692 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_301
timestamp 1688980957
transform 1 0 28796 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_307
timestamp 1688980957
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_309
timestamp 1688980957
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_321
timestamp 1688980957
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_333
timestamp 1688980957
transform 1 0 31740 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_345
timestamp 1688980957
transform 1 0 32844 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_357
timestamp 1688980957
transform 1 0 33948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_363
timestamp 1688980957
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_365
timestamp 1688980957
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_377
timestamp 1688980957
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_389
timestamp 1688980957
transform 1 0 36892 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_401
timestamp 1688980957
transform 1 0 37996 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_413
timestamp 1688980957
transform 1 0 39100 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_419
timestamp 1688980957
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_421
timestamp 1688980957
transform 1 0 39836 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_433
timestamp 1688980957
transform 1 0 40940 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_445
timestamp 1688980957
transform 1 0 42044 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_457
timestamp 1688980957
transform 1 0 43148 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_469
timestamp 1688980957
transform 1 0 44252 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_475
timestamp 1688980957
transform 1 0 44804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_477
timestamp 1688980957
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_489
timestamp 1688980957
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_501
timestamp 1688980957
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_513
timestamp 1688980957
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_525
timestamp 1688980957
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_531
timestamp 1688980957
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_533
timestamp 1688980957
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_545
timestamp 1688980957
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_557
timestamp 1688980957
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_569
timestamp 1688980957
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_581
timestamp 1688980957
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_587
timestamp 1688980957
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_589
timestamp 1688980957
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_601
timestamp 1688980957
transform 1 0 56396 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_613
timestamp 1688980957
transform 1 0 57500 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_625
timestamp 1688980957
transform 1 0 58604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_637
timestamp 1688980957
transform 1 0 59708 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_643
timestamp 1688980957
transform 1 0 60260 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_645
timestamp 1688980957
transform 1 0 60444 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_657
timestamp 1688980957
transform 1 0 61548 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_669
timestamp 1688980957
transform 1 0 62652 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_681
timestamp 1688980957
transform 1 0 63756 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_693
timestamp 1688980957
transform 1 0 64860 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_699
timestamp 1688980957
transform 1 0 65412 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_701
timestamp 1688980957
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_713
timestamp 1688980957
transform 1 0 66700 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_725
timestamp 1688980957
transform 1 0 67804 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_3
timestamp 1688980957
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_15
timestamp 1688980957
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_27
timestamp 1688980957
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_39
timestamp 1688980957
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_51
timestamp 1688980957
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_55
timestamp 1688980957
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_57
timestamp 1688980957
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_69
timestamp 1688980957
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_81
timestamp 1688980957
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_93
timestamp 1688980957
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_105
timestamp 1688980957
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_111
timestamp 1688980957
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_113
timestamp 1688980957
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_125
timestamp 1688980957
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_137
timestamp 1688980957
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_149
timestamp 1688980957
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_161
timestamp 1688980957
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_167
timestamp 1688980957
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_169
timestamp 1688980957
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_181
timestamp 1688980957
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_193
timestamp 1688980957
transform 1 0 18860 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_205
timestamp 1688980957
transform 1 0 19964 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_217
timestamp 1688980957
transform 1 0 21068 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_223
timestamp 1688980957
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_225
timestamp 1688980957
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_237
timestamp 1688980957
transform 1 0 22908 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_249
timestamp 1688980957
transform 1 0 24012 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_261
timestamp 1688980957
transform 1 0 25116 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_273
timestamp 1688980957
transform 1 0 26220 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_279
timestamp 1688980957
transform 1 0 26772 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_281
timestamp 1688980957
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_293
timestamp 1688980957
transform 1 0 28060 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_305
timestamp 1688980957
transform 1 0 29164 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_317
timestamp 1688980957
transform 1 0 30268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_329
timestamp 1688980957
transform 1 0 31372 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_335
timestamp 1688980957
transform 1 0 31924 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_337
timestamp 1688980957
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_349
timestamp 1688980957
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_361
timestamp 1688980957
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_373
timestamp 1688980957
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_385
timestamp 1688980957
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_391
timestamp 1688980957
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_393
timestamp 1688980957
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_405
timestamp 1688980957
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_417
timestamp 1688980957
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_429
timestamp 1688980957
transform 1 0 40572 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_441
timestamp 1688980957
transform 1 0 41676 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_447
timestamp 1688980957
transform 1 0 42228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_449
timestamp 1688980957
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_461
timestamp 1688980957
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_473
timestamp 1688980957
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_485
timestamp 1688980957
transform 1 0 45724 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_497
timestamp 1688980957
transform 1 0 46828 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_503
timestamp 1688980957
transform 1 0 47380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_505
timestamp 1688980957
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_517
timestamp 1688980957
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_529
timestamp 1688980957
transform 1 0 49772 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_541
timestamp 1688980957
transform 1 0 50876 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_553
timestamp 1688980957
transform 1 0 51980 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_559
timestamp 1688980957
transform 1 0 52532 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_561
timestamp 1688980957
transform 1 0 52716 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_573
timestamp 1688980957
transform 1 0 53820 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_585
timestamp 1688980957
transform 1 0 54924 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_597
timestamp 1688980957
transform 1 0 56028 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_609
timestamp 1688980957
transform 1 0 57132 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_615
timestamp 1688980957
transform 1 0 57684 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_617
timestamp 1688980957
transform 1 0 57868 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_629
timestamp 1688980957
transform 1 0 58972 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_641
timestamp 1688980957
transform 1 0 60076 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_653
timestamp 1688980957
transform 1 0 61180 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_665
timestamp 1688980957
transform 1 0 62284 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_671
timestamp 1688980957
transform 1 0 62836 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_673
timestamp 1688980957
transform 1 0 63020 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_685
timestamp 1688980957
transform 1 0 64124 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_697
timestamp 1688980957
transform 1 0 65228 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_709
timestamp 1688980957
transform 1 0 66332 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_107_721
timestamp 1688980957
transform 1 0 67436 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107_726
timestamp 1688980957
transform 1 0 67896 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_3
timestamp 1688980957
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_15
timestamp 1688980957
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_27
timestamp 1688980957
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_29
timestamp 1688980957
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_41
timestamp 1688980957
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_53
timestamp 1688980957
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_65
timestamp 1688980957
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_77
timestamp 1688980957
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_83
timestamp 1688980957
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_85
timestamp 1688980957
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_97
timestamp 1688980957
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_109
timestamp 1688980957
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_121
timestamp 1688980957
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_133
timestamp 1688980957
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_139
timestamp 1688980957
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_141
timestamp 1688980957
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_153
timestamp 1688980957
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_165
timestamp 1688980957
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_177
timestamp 1688980957
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_189
timestamp 1688980957
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_195
timestamp 1688980957
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_197
timestamp 1688980957
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_209
timestamp 1688980957
transform 1 0 20332 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_221
timestamp 1688980957
transform 1 0 21436 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_233
timestamp 1688980957
transform 1 0 22540 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_245
timestamp 1688980957
transform 1 0 23644 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_251
timestamp 1688980957
transform 1 0 24196 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_253
timestamp 1688980957
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_265
timestamp 1688980957
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_277
timestamp 1688980957
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_289
timestamp 1688980957
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_301
timestamp 1688980957
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_307
timestamp 1688980957
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_309
timestamp 1688980957
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_321
timestamp 1688980957
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_333
timestamp 1688980957
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_345
timestamp 1688980957
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_357
timestamp 1688980957
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_363
timestamp 1688980957
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_365
timestamp 1688980957
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_377
timestamp 1688980957
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_389
timestamp 1688980957
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_401
timestamp 1688980957
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_413
timestamp 1688980957
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_419
timestamp 1688980957
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_421
timestamp 1688980957
transform 1 0 39836 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_433
timestamp 1688980957
transform 1 0 40940 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_445
timestamp 1688980957
transform 1 0 42044 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_457
timestamp 1688980957
transform 1 0 43148 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_469
timestamp 1688980957
transform 1 0 44252 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_475
timestamp 1688980957
transform 1 0 44804 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_477
timestamp 1688980957
transform 1 0 44988 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_489
timestamp 1688980957
transform 1 0 46092 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_501
timestamp 1688980957
transform 1 0 47196 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_513
timestamp 1688980957
transform 1 0 48300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_525
timestamp 1688980957
transform 1 0 49404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_531
timestamp 1688980957
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_533
timestamp 1688980957
transform 1 0 50140 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_545
timestamp 1688980957
transform 1 0 51244 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_557
timestamp 1688980957
transform 1 0 52348 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_569
timestamp 1688980957
transform 1 0 53452 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_581
timestamp 1688980957
transform 1 0 54556 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_587
timestamp 1688980957
transform 1 0 55108 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_589
timestamp 1688980957
transform 1 0 55292 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_601
timestamp 1688980957
transform 1 0 56396 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_613
timestamp 1688980957
transform 1 0 57500 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_625
timestamp 1688980957
transform 1 0 58604 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_637
timestamp 1688980957
transform 1 0 59708 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_643
timestamp 1688980957
transform 1 0 60260 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_645
timestamp 1688980957
transform 1 0 60444 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_657
timestamp 1688980957
transform 1 0 61548 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_669
timestamp 1688980957
transform 1 0 62652 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_681
timestamp 1688980957
transform 1 0 63756 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_693
timestamp 1688980957
transform 1 0 64860 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_699
timestamp 1688980957
transform 1 0 65412 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_701
timestamp 1688980957
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_713
timestamp 1688980957
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_725
timestamp 1688980957
transform 1 0 67804 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_3
timestamp 1688980957
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_15
timestamp 1688980957
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_27
timestamp 1688980957
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_39
timestamp 1688980957
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_51
timestamp 1688980957
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_55
timestamp 1688980957
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_57
timestamp 1688980957
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_69
timestamp 1688980957
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_81
timestamp 1688980957
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_93
timestamp 1688980957
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_105
timestamp 1688980957
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_111
timestamp 1688980957
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_113
timestamp 1688980957
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_125
timestamp 1688980957
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_137
timestamp 1688980957
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_149
timestamp 1688980957
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_161
timestamp 1688980957
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_167
timestamp 1688980957
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_169
timestamp 1688980957
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_181
timestamp 1688980957
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_193
timestamp 1688980957
transform 1 0 18860 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_205
timestamp 1688980957
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_217
timestamp 1688980957
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_223
timestamp 1688980957
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_225
timestamp 1688980957
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_237
timestamp 1688980957
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_249
timestamp 1688980957
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_261
timestamp 1688980957
transform 1 0 25116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_273
timestamp 1688980957
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_279
timestamp 1688980957
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_281
timestamp 1688980957
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_293
timestamp 1688980957
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_305
timestamp 1688980957
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_317
timestamp 1688980957
transform 1 0 30268 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_329
timestamp 1688980957
transform 1 0 31372 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_335
timestamp 1688980957
transform 1 0 31924 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_337
timestamp 1688980957
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_349
timestamp 1688980957
transform 1 0 33212 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_361
timestamp 1688980957
transform 1 0 34316 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_373
timestamp 1688980957
transform 1 0 35420 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_385
timestamp 1688980957
transform 1 0 36524 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_391
timestamp 1688980957
transform 1 0 37076 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_393
timestamp 1688980957
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_405
timestamp 1688980957
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_417
timestamp 1688980957
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_429
timestamp 1688980957
transform 1 0 40572 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_441
timestamp 1688980957
transform 1 0 41676 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_447
timestamp 1688980957
transform 1 0 42228 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_449
timestamp 1688980957
transform 1 0 42412 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_461
timestamp 1688980957
transform 1 0 43516 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_473
timestamp 1688980957
transform 1 0 44620 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_485
timestamp 1688980957
transform 1 0 45724 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_497
timestamp 1688980957
transform 1 0 46828 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_503
timestamp 1688980957
transform 1 0 47380 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_505
timestamp 1688980957
transform 1 0 47564 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_517
timestamp 1688980957
transform 1 0 48668 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_529
timestamp 1688980957
transform 1 0 49772 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_541
timestamp 1688980957
transform 1 0 50876 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_553
timestamp 1688980957
transform 1 0 51980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_559
timestamp 1688980957
transform 1 0 52532 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_561
timestamp 1688980957
transform 1 0 52716 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_573
timestamp 1688980957
transform 1 0 53820 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_585
timestamp 1688980957
transform 1 0 54924 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_597
timestamp 1688980957
transform 1 0 56028 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_609
timestamp 1688980957
transform 1 0 57132 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_615
timestamp 1688980957
transform 1 0 57684 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_617
timestamp 1688980957
transform 1 0 57868 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_629
timestamp 1688980957
transform 1 0 58972 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_641
timestamp 1688980957
transform 1 0 60076 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_653
timestamp 1688980957
transform 1 0 61180 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_665
timestamp 1688980957
transform 1 0 62284 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_671
timestamp 1688980957
transform 1 0 62836 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_673
timestamp 1688980957
transform 1 0 63020 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_685
timestamp 1688980957
transform 1 0 64124 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_697
timestamp 1688980957
transform 1 0 65228 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_709
timestamp 1688980957
transform 1 0 66332 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_721
timestamp 1688980957
transform 1 0 67436 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_727
timestamp 1688980957
transform 1 0 67988 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_729
timestamp 1688980957
transform 1 0 68172 0 -1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_3
timestamp 1688980957
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_15
timestamp 1688980957
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_27
timestamp 1688980957
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_29
timestamp 1688980957
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_41
timestamp 1688980957
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_53
timestamp 1688980957
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_65
timestamp 1688980957
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_77
timestamp 1688980957
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_83
timestamp 1688980957
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_85
timestamp 1688980957
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_97
timestamp 1688980957
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_109
timestamp 1688980957
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_121
timestamp 1688980957
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_133
timestamp 1688980957
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_139
timestamp 1688980957
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_141
timestamp 1688980957
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_153
timestamp 1688980957
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_165
timestamp 1688980957
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_177
timestamp 1688980957
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_189
timestamp 1688980957
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_195
timestamp 1688980957
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_197
timestamp 1688980957
transform 1 0 19228 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_209
timestamp 1688980957
transform 1 0 20332 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_221
timestamp 1688980957
transform 1 0 21436 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_233
timestamp 1688980957
transform 1 0 22540 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_245
timestamp 1688980957
transform 1 0 23644 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_251
timestamp 1688980957
transform 1 0 24196 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_253
timestamp 1688980957
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_265
timestamp 1688980957
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_277
timestamp 1688980957
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_289
timestamp 1688980957
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_301
timestamp 1688980957
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_307
timestamp 1688980957
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_309
timestamp 1688980957
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_321
timestamp 1688980957
transform 1 0 30636 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_333
timestamp 1688980957
transform 1 0 31740 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_345
timestamp 1688980957
transform 1 0 32844 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_357
timestamp 1688980957
transform 1 0 33948 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_363
timestamp 1688980957
transform 1 0 34500 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_365
timestamp 1688980957
transform 1 0 34684 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_377
timestamp 1688980957
transform 1 0 35788 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_389
timestamp 1688980957
transform 1 0 36892 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_401
timestamp 1688980957
transform 1 0 37996 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_413
timestamp 1688980957
transform 1 0 39100 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_419
timestamp 1688980957
transform 1 0 39652 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_421
timestamp 1688980957
transform 1 0 39836 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_433
timestamp 1688980957
transform 1 0 40940 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_445
timestamp 1688980957
transform 1 0 42044 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_457
timestamp 1688980957
transform 1 0 43148 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_469
timestamp 1688980957
transform 1 0 44252 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_475
timestamp 1688980957
transform 1 0 44804 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_477
timestamp 1688980957
transform 1 0 44988 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_489
timestamp 1688980957
transform 1 0 46092 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_501
timestamp 1688980957
transform 1 0 47196 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_513
timestamp 1688980957
transform 1 0 48300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_525
timestamp 1688980957
transform 1 0 49404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_531
timestamp 1688980957
transform 1 0 49956 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_533
timestamp 1688980957
transform 1 0 50140 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_545
timestamp 1688980957
transform 1 0 51244 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_557
timestamp 1688980957
transform 1 0 52348 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_569
timestamp 1688980957
transform 1 0 53452 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_581
timestamp 1688980957
transform 1 0 54556 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_587
timestamp 1688980957
transform 1 0 55108 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_589
timestamp 1688980957
transform 1 0 55292 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_601
timestamp 1688980957
transform 1 0 56396 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_613
timestamp 1688980957
transform 1 0 57500 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_625
timestamp 1688980957
transform 1 0 58604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_637
timestamp 1688980957
transform 1 0 59708 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_643
timestamp 1688980957
transform 1 0 60260 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_645
timestamp 1688980957
transform 1 0 60444 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_657
timestamp 1688980957
transform 1 0 61548 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_669
timestamp 1688980957
transform 1 0 62652 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_681
timestamp 1688980957
transform 1 0 63756 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_693
timestamp 1688980957
transform 1 0 64860 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_699
timestamp 1688980957
transform 1 0 65412 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_701
timestamp 1688980957
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_713
timestamp 1688980957
transform 1 0 66700 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_725
timestamp 1688980957
transform 1 0 67804 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_3
timestamp 1688980957
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_15
timestamp 1688980957
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_27
timestamp 1688980957
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_39
timestamp 1688980957
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_51
timestamp 1688980957
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_55
timestamp 1688980957
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_57
timestamp 1688980957
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_69
timestamp 1688980957
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_81
timestamp 1688980957
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_93
timestamp 1688980957
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_105
timestamp 1688980957
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_111
timestamp 1688980957
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_113
timestamp 1688980957
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_125
timestamp 1688980957
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_137
timestamp 1688980957
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_149
timestamp 1688980957
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_161
timestamp 1688980957
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_167
timestamp 1688980957
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_169
timestamp 1688980957
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_181
timestamp 1688980957
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_193
timestamp 1688980957
transform 1 0 18860 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_205
timestamp 1688980957
transform 1 0 19964 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_217
timestamp 1688980957
transform 1 0 21068 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_223
timestamp 1688980957
transform 1 0 21620 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_225
timestamp 1688980957
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_237
timestamp 1688980957
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_249
timestamp 1688980957
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_261
timestamp 1688980957
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_273
timestamp 1688980957
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_279
timestamp 1688980957
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_281
timestamp 1688980957
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_293
timestamp 1688980957
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_305
timestamp 1688980957
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_317
timestamp 1688980957
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_329
timestamp 1688980957
transform 1 0 31372 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_335
timestamp 1688980957
transform 1 0 31924 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_337
timestamp 1688980957
transform 1 0 32108 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_349
timestamp 1688980957
transform 1 0 33212 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_361
timestamp 1688980957
transform 1 0 34316 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_373
timestamp 1688980957
transform 1 0 35420 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_385
timestamp 1688980957
transform 1 0 36524 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_391
timestamp 1688980957
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_393
timestamp 1688980957
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_405
timestamp 1688980957
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_417
timestamp 1688980957
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_429
timestamp 1688980957
transform 1 0 40572 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_441
timestamp 1688980957
transform 1 0 41676 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_447
timestamp 1688980957
transform 1 0 42228 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_449
timestamp 1688980957
transform 1 0 42412 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_461
timestamp 1688980957
transform 1 0 43516 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_473
timestamp 1688980957
transform 1 0 44620 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_485
timestamp 1688980957
transform 1 0 45724 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_497
timestamp 1688980957
transform 1 0 46828 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_503
timestamp 1688980957
transform 1 0 47380 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_505
timestamp 1688980957
transform 1 0 47564 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_517
timestamp 1688980957
transform 1 0 48668 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_529
timestamp 1688980957
transform 1 0 49772 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_541
timestamp 1688980957
transform 1 0 50876 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_553
timestamp 1688980957
transform 1 0 51980 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_559
timestamp 1688980957
transform 1 0 52532 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_561
timestamp 1688980957
transform 1 0 52716 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_573
timestamp 1688980957
transform 1 0 53820 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_585
timestamp 1688980957
transform 1 0 54924 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_597
timestamp 1688980957
transform 1 0 56028 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_609
timestamp 1688980957
transform 1 0 57132 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_615
timestamp 1688980957
transform 1 0 57684 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_617
timestamp 1688980957
transform 1 0 57868 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_629
timestamp 1688980957
transform 1 0 58972 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_641
timestamp 1688980957
transform 1 0 60076 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_653
timestamp 1688980957
transform 1 0 61180 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_665
timestamp 1688980957
transform 1 0 62284 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_671
timestamp 1688980957
transform 1 0 62836 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_673
timestamp 1688980957
transform 1 0 63020 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_685
timestamp 1688980957
transform 1 0 64124 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_697
timestamp 1688980957
transform 1 0 65228 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_709
timestamp 1688980957
transform 1 0 66332 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_721
timestamp 1688980957
transform 1 0 67436 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_727
timestamp 1688980957
transform 1 0 67988 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_729
timestamp 1688980957
transform 1 0 68172 0 -1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_3
timestamp 1688980957
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_15
timestamp 1688980957
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_27
timestamp 1688980957
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_29
timestamp 1688980957
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_41
timestamp 1688980957
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_53
timestamp 1688980957
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_65
timestamp 1688980957
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_77
timestamp 1688980957
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_83
timestamp 1688980957
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_85
timestamp 1688980957
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_97
timestamp 1688980957
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_109
timestamp 1688980957
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_121
timestamp 1688980957
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_133
timestamp 1688980957
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_139
timestamp 1688980957
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_141
timestamp 1688980957
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_153
timestamp 1688980957
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_165
timestamp 1688980957
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_177
timestamp 1688980957
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_189
timestamp 1688980957
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_195
timestamp 1688980957
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_197
timestamp 1688980957
transform 1 0 19228 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_209
timestamp 1688980957
transform 1 0 20332 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_221
timestamp 1688980957
transform 1 0 21436 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_233
timestamp 1688980957
transform 1 0 22540 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_245
timestamp 1688980957
transform 1 0 23644 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_251
timestamp 1688980957
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_253
timestamp 1688980957
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_265
timestamp 1688980957
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_277
timestamp 1688980957
transform 1 0 26588 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_289
timestamp 1688980957
transform 1 0 27692 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_301
timestamp 1688980957
transform 1 0 28796 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_307
timestamp 1688980957
transform 1 0 29348 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_309
timestamp 1688980957
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_321
timestamp 1688980957
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_333
timestamp 1688980957
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_345
timestamp 1688980957
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_357
timestamp 1688980957
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_363
timestamp 1688980957
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_365
timestamp 1688980957
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_377
timestamp 1688980957
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_389
timestamp 1688980957
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_401
timestamp 1688980957
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_413
timestamp 1688980957
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_419
timestamp 1688980957
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_421
timestamp 1688980957
transform 1 0 39836 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_433
timestamp 1688980957
transform 1 0 40940 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_445
timestamp 1688980957
transform 1 0 42044 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_457
timestamp 1688980957
transform 1 0 43148 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_469
timestamp 1688980957
transform 1 0 44252 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_475
timestamp 1688980957
transform 1 0 44804 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_477
timestamp 1688980957
transform 1 0 44988 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_489
timestamp 1688980957
transform 1 0 46092 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_501
timestamp 1688980957
transform 1 0 47196 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_513
timestamp 1688980957
transform 1 0 48300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_525
timestamp 1688980957
transform 1 0 49404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_531
timestamp 1688980957
transform 1 0 49956 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_533
timestamp 1688980957
transform 1 0 50140 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_545
timestamp 1688980957
transform 1 0 51244 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_557
timestamp 1688980957
transform 1 0 52348 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_569
timestamp 1688980957
transform 1 0 53452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_581
timestamp 1688980957
transform 1 0 54556 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_587
timestamp 1688980957
transform 1 0 55108 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_589
timestamp 1688980957
transform 1 0 55292 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_601
timestamp 1688980957
transform 1 0 56396 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_613
timestamp 1688980957
transform 1 0 57500 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_625
timestamp 1688980957
transform 1 0 58604 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_637
timestamp 1688980957
transform 1 0 59708 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_643
timestamp 1688980957
transform 1 0 60260 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_645
timestamp 1688980957
transform 1 0 60444 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_657
timestamp 1688980957
transform 1 0 61548 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_669
timestamp 1688980957
transform 1 0 62652 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_681
timestamp 1688980957
transform 1 0 63756 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_693
timestamp 1688980957
transform 1 0 64860 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_699
timestamp 1688980957
transform 1 0 65412 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_701
timestamp 1688980957
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_713
timestamp 1688980957
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112_725
timestamp 1688980957
transform 1 0 67804 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_729
timestamp 1688980957
transform 1 0 68172 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_3
timestamp 1688980957
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_15
timestamp 1688980957
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_27
timestamp 1688980957
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_39
timestamp 1688980957
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_51
timestamp 1688980957
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_55
timestamp 1688980957
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_57
timestamp 1688980957
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_69
timestamp 1688980957
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_81
timestamp 1688980957
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_93
timestamp 1688980957
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_105
timestamp 1688980957
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_111
timestamp 1688980957
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_113
timestamp 1688980957
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_125
timestamp 1688980957
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_137
timestamp 1688980957
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_149
timestamp 1688980957
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_161
timestamp 1688980957
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_167
timestamp 1688980957
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_169
timestamp 1688980957
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_181
timestamp 1688980957
transform 1 0 17756 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_193
timestamp 1688980957
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_205
timestamp 1688980957
transform 1 0 19964 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_217
timestamp 1688980957
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_223
timestamp 1688980957
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_225
timestamp 1688980957
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_237
timestamp 1688980957
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_249
timestamp 1688980957
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_261
timestamp 1688980957
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_273
timestamp 1688980957
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_279
timestamp 1688980957
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_281
timestamp 1688980957
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_293
timestamp 1688980957
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_305
timestamp 1688980957
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_317
timestamp 1688980957
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_329
timestamp 1688980957
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_335
timestamp 1688980957
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_337
timestamp 1688980957
transform 1 0 32108 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_349
timestamp 1688980957
transform 1 0 33212 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_361
timestamp 1688980957
transform 1 0 34316 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_373
timestamp 1688980957
transform 1 0 35420 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_385
timestamp 1688980957
transform 1 0 36524 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_391
timestamp 1688980957
transform 1 0 37076 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_393
timestamp 1688980957
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_405
timestamp 1688980957
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_417
timestamp 1688980957
transform 1 0 39468 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_429
timestamp 1688980957
transform 1 0 40572 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_441
timestamp 1688980957
transform 1 0 41676 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_447
timestamp 1688980957
transform 1 0 42228 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_449
timestamp 1688980957
transform 1 0 42412 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_461
timestamp 1688980957
transform 1 0 43516 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_473
timestamp 1688980957
transform 1 0 44620 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_485
timestamp 1688980957
transform 1 0 45724 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_497
timestamp 1688980957
transform 1 0 46828 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_503
timestamp 1688980957
transform 1 0 47380 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_505
timestamp 1688980957
transform 1 0 47564 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_517
timestamp 1688980957
transform 1 0 48668 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_529
timestamp 1688980957
transform 1 0 49772 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_541
timestamp 1688980957
transform 1 0 50876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_553
timestamp 1688980957
transform 1 0 51980 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_559
timestamp 1688980957
transform 1 0 52532 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_561
timestamp 1688980957
transform 1 0 52716 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_573
timestamp 1688980957
transform 1 0 53820 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_585
timestamp 1688980957
transform 1 0 54924 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_597
timestamp 1688980957
transform 1 0 56028 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_609
timestamp 1688980957
transform 1 0 57132 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_615
timestamp 1688980957
transform 1 0 57684 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_617
timestamp 1688980957
transform 1 0 57868 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_629
timestamp 1688980957
transform 1 0 58972 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_641
timestamp 1688980957
transform 1 0 60076 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_653
timestamp 1688980957
transform 1 0 61180 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_665
timestamp 1688980957
transform 1 0 62284 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_671
timestamp 1688980957
transform 1 0 62836 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_673
timestamp 1688980957
transform 1 0 63020 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_685
timestamp 1688980957
transform 1 0 64124 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_697
timestamp 1688980957
transform 1 0 65228 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_709
timestamp 1688980957
transform 1 0 66332 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_721
timestamp 1688980957
transform 1 0 67436 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_727
timestamp 1688980957
transform 1 0 67988 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_729
timestamp 1688980957
transform 1 0 68172 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_3
timestamp 1688980957
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_15
timestamp 1688980957
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_27
timestamp 1688980957
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_29
timestamp 1688980957
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_41
timestamp 1688980957
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_53
timestamp 1688980957
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_65
timestamp 1688980957
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_77
timestamp 1688980957
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_83
timestamp 1688980957
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_85
timestamp 1688980957
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_97
timestamp 1688980957
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_109
timestamp 1688980957
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_121
timestamp 1688980957
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_133
timestamp 1688980957
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_139
timestamp 1688980957
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_141
timestamp 1688980957
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_153
timestamp 1688980957
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_165
timestamp 1688980957
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_177
timestamp 1688980957
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_189
timestamp 1688980957
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_195
timestamp 1688980957
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_197
timestamp 1688980957
transform 1 0 19228 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_209
timestamp 1688980957
transform 1 0 20332 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_221
timestamp 1688980957
transform 1 0 21436 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_233
timestamp 1688980957
transform 1 0 22540 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_245
timestamp 1688980957
transform 1 0 23644 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_251
timestamp 1688980957
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_253
timestamp 1688980957
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_265
timestamp 1688980957
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_277
timestamp 1688980957
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_289
timestamp 1688980957
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_301
timestamp 1688980957
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_307
timestamp 1688980957
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_309
timestamp 1688980957
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_321
timestamp 1688980957
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_333
timestamp 1688980957
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_345
timestamp 1688980957
transform 1 0 32844 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_357
timestamp 1688980957
transform 1 0 33948 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_363
timestamp 1688980957
transform 1 0 34500 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_365
timestamp 1688980957
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_377
timestamp 1688980957
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_389
timestamp 1688980957
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_401
timestamp 1688980957
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_413
timestamp 1688980957
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_419
timestamp 1688980957
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_421
timestamp 1688980957
transform 1 0 39836 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_433
timestamp 1688980957
transform 1 0 40940 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_445
timestamp 1688980957
transform 1 0 42044 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_457
timestamp 1688980957
transform 1 0 43148 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_469
timestamp 1688980957
transform 1 0 44252 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_475
timestamp 1688980957
transform 1 0 44804 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_477
timestamp 1688980957
transform 1 0 44988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_489
timestamp 1688980957
transform 1 0 46092 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_501
timestamp 1688980957
transform 1 0 47196 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_513
timestamp 1688980957
transform 1 0 48300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_525
timestamp 1688980957
transform 1 0 49404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_531
timestamp 1688980957
transform 1 0 49956 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_533
timestamp 1688980957
transform 1 0 50140 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_545
timestamp 1688980957
transform 1 0 51244 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_557
timestamp 1688980957
transform 1 0 52348 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_569
timestamp 1688980957
transform 1 0 53452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_581
timestamp 1688980957
transform 1 0 54556 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_587
timestamp 1688980957
transform 1 0 55108 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_589
timestamp 1688980957
transform 1 0 55292 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_601
timestamp 1688980957
transform 1 0 56396 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_613
timestamp 1688980957
transform 1 0 57500 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_625
timestamp 1688980957
transform 1 0 58604 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_637
timestamp 1688980957
transform 1 0 59708 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_643
timestamp 1688980957
transform 1 0 60260 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_645
timestamp 1688980957
transform 1 0 60444 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_657
timestamp 1688980957
transform 1 0 61548 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_669
timestamp 1688980957
transform 1 0 62652 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_681
timestamp 1688980957
transform 1 0 63756 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_693
timestamp 1688980957
transform 1 0 64860 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_699
timestamp 1688980957
transform 1 0 65412 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_701
timestamp 1688980957
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_713
timestamp 1688980957
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_725
timestamp 1688980957
transform 1 0 67804 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_6
timestamp 1688980957
transform 1 0 1656 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_18
timestamp 1688980957
transform 1 0 2760 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_30
timestamp 1688980957
transform 1 0 3864 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_42
timestamp 1688980957
transform 1 0 4968 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115_54
timestamp 1688980957
transform 1 0 6072 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_57
timestamp 1688980957
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_69
timestamp 1688980957
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_81
timestamp 1688980957
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_93
timestamp 1688980957
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_105
timestamp 1688980957
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_111
timestamp 1688980957
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_113
timestamp 1688980957
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_125
timestamp 1688980957
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_137
timestamp 1688980957
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_149
timestamp 1688980957
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_161
timestamp 1688980957
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_167
timestamp 1688980957
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_169
timestamp 1688980957
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_181
timestamp 1688980957
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_193
timestamp 1688980957
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_205
timestamp 1688980957
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_217
timestamp 1688980957
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_223
timestamp 1688980957
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_225
timestamp 1688980957
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_237
timestamp 1688980957
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_249
timestamp 1688980957
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_261
timestamp 1688980957
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_273
timestamp 1688980957
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_279
timestamp 1688980957
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_281
timestamp 1688980957
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_293
timestamp 1688980957
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_305
timestamp 1688980957
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_317
timestamp 1688980957
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_329
timestamp 1688980957
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_335
timestamp 1688980957
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_337
timestamp 1688980957
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_349
timestamp 1688980957
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_361
timestamp 1688980957
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_373
timestamp 1688980957
transform 1 0 35420 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_385
timestamp 1688980957
transform 1 0 36524 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_391
timestamp 1688980957
transform 1 0 37076 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_393
timestamp 1688980957
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_405
timestamp 1688980957
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_417
timestamp 1688980957
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_429
timestamp 1688980957
transform 1 0 40572 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_441
timestamp 1688980957
transform 1 0 41676 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_447
timestamp 1688980957
transform 1 0 42228 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_449
timestamp 1688980957
transform 1 0 42412 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_461
timestamp 1688980957
transform 1 0 43516 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_473
timestamp 1688980957
transform 1 0 44620 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_485
timestamp 1688980957
transform 1 0 45724 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_497
timestamp 1688980957
transform 1 0 46828 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_503
timestamp 1688980957
transform 1 0 47380 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_505
timestamp 1688980957
transform 1 0 47564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_517
timestamp 1688980957
transform 1 0 48668 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_529
timestamp 1688980957
transform 1 0 49772 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_541
timestamp 1688980957
transform 1 0 50876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_553
timestamp 1688980957
transform 1 0 51980 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_559
timestamp 1688980957
transform 1 0 52532 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_561
timestamp 1688980957
transform 1 0 52716 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_573
timestamp 1688980957
transform 1 0 53820 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_585
timestamp 1688980957
transform 1 0 54924 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_597
timestamp 1688980957
transform 1 0 56028 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_609
timestamp 1688980957
transform 1 0 57132 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_615
timestamp 1688980957
transform 1 0 57684 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_617
timestamp 1688980957
transform 1 0 57868 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_629
timestamp 1688980957
transform 1 0 58972 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_641
timestamp 1688980957
transform 1 0 60076 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_653
timestamp 1688980957
transform 1 0 61180 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_665
timestamp 1688980957
transform 1 0 62284 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_671
timestamp 1688980957
transform 1 0 62836 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_673
timestamp 1688980957
transform 1 0 63020 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_685
timestamp 1688980957
transform 1 0 64124 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_697
timestamp 1688980957
transform 1 0 65228 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_709
timestamp 1688980957
transform 1 0 66332 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_721
timestamp 1688980957
transform 1 0 67436 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_727
timestamp 1688980957
transform 1 0 67988 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_729
timestamp 1688980957
transform 1 0 68172 0 -1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_3
timestamp 1688980957
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_15
timestamp 1688980957
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_27
timestamp 1688980957
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_29
timestamp 1688980957
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_41
timestamp 1688980957
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_53
timestamp 1688980957
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_65
timestamp 1688980957
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_77
timestamp 1688980957
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_83
timestamp 1688980957
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_85
timestamp 1688980957
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_97
timestamp 1688980957
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_109
timestamp 1688980957
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_121
timestamp 1688980957
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_133
timestamp 1688980957
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_139
timestamp 1688980957
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_141
timestamp 1688980957
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_153
timestamp 1688980957
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_165
timestamp 1688980957
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_177
timestamp 1688980957
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_189
timestamp 1688980957
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_195
timestamp 1688980957
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_197
timestamp 1688980957
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_209
timestamp 1688980957
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_221
timestamp 1688980957
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_233
timestamp 1688980957
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_245
timestamp 1688980957
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_251
timestamp 1688980957
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_253
timestamp 1688980957
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_265
timestamp 1688980957
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_277
timestamp 1688980957
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_289
timestamp 1688980957
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_301
timestamp 1688980957
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_307
timestamp 1688980957
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_309
timestamp 1688980957
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_321
timestamp 1688980957
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_333
timestamp 1688980957
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_345
timestamp 1688980957
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_357
timestamp 1688980957
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_363
timestamp 1688980957
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_365
timestamp 1688980957
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_377
timestamp 1688980957
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_389
timestamp 1688980957
transform 1 0 36892 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_401
timestamp 1688980957
transform 1 0 37996 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_413
timestamp 1688980957
transform 1 0 39100 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_419
timestamp 1688980957
transform 1 0 39652 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_421
timestamp 1688980957
transform 1 0 39836 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_433
timestamp 1688980957
transform 1 0 40940 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_445
timestamp 1688980957
transform 1 0 42044 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_457
timestamp 1688980957
transform 1 0 43148 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_469
timestamp 1688980957
transform 1 0 44252 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_475
timestamp 1688980957
transform 1 0 44804 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_477
timestamp 1688980957
transform 1 0 44988 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_489
timestamp 1688980957
transform 1 0 46092 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_501
timestamp 1688980957
transform 1 0 47196 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_513
timestamp 1688980957
transform 1 0 48300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_525
timestamp 1688980957
transform 1 0 49404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_531
timestamp 1688980957
transform 1 0 49956 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_533
timestamp 1688980957
transform 1 0 50140 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_545
timestamp 1688980957
transform 1 0 51244 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_557
timestamp 1688980957
transform 1 0 52348 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_569
timestamp 1688980957
transform 1 0 53452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_581
timestamp 1688980957
transform 1 0 54556 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_587
timestamp 1688980957
transform 1 0 55108 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_589
timestamp 1688980957
transform 1 0 55292 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_601
timestamp 1688980957
transform 1 0 56396 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_613
timestamp 1688980957
transform 1 0 57500 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_625
timestamp 1688980957
transform 1 0 58604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_637
timestamp 1688980957
transform 1 0 59708 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_643
timestamp 1688980957
transform 1 0 60260 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_645
timestamp 1688980957
transform 1 0 60444 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_657
timestamp 1688980957
transform 1 0 61548 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_669
timestamp 1688980957
transform 1 0 62652 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_681
timestamp 1688980957
transform 1 0 63756 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_693
timestamp 1688980957
transform 1 0 64860 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_699
timestamp 1688980957
transform 1 0 65412 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_701
timestamp 1688980957
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_713
timestamp 1688980957
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_725
timestamp 1688980957
transform 1 0 67804 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_3
timestamp 1688980957
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_15
timestamp 1688980957
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_27
timestamp 1688980957
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_39
timestamp 1688980957
transform 1 0 4692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_51
timestamp 1688980957
transform 1 0 5796 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_55
timestamp 1688980957
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_57
timestamp 1688980957
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_69
timestamp 1688980957
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_81
timestamp 1688980957
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_93
timestamp 1688980957
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_105
timestamp 1688980957
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_111
timestamp 1688980957
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_113
timestamp 1688980957
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_125
timestamp 1688980957
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_137
timestamp 1688980957
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_149
timestamp 1688980957
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_161
timestamp 1688980957
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_167
timestamp 1688980957
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_169
timestamp 1688980957
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_181
timestamp 1688980957
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_193
timestamp 1688980957
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_205
timestamp 1688980957
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_217
timestamp 1688980957
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_223
timestamp 1688980957
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_225
timestamp 1688980957
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_237
timestamp 1688980957
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_249
timestamp 1688980957
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_261
timestamp 1688980957
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_273
timestamp 1688980957
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_279
timestamp 1688980957
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_281
timestamp 1688980957
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_293
timestamp 1688980957
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_305
timestamp 1688980957
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_317
timestamp 1688980957
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_329
timestamp 1688980957
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_335
timestamp 1688980957
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_337
timestamp 1688980957
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_349
timestamp 1688980957
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_361
timestamp 1688980957
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_373
timestamp 1688980957
transform 1 0 35420 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_385
timestamp 1688980957
transform 1 0 36524 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_391
timestamp 1688980957
transform 1 0 37076 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_393
timestamp 1688980957
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_405
timestamp 1688980957
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_417
timestamp 1688980957
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_429
timestamp 1688980957
transform 1 0 40572 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_441
timestamp 1688980957
transform 1 0 41676 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_447
timestamp 1688980957
transform 1 0 42228 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_449
timestamp 1688980957
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_461
timestamp 1688980957
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_473
timestamp 1688980957
transform 1 0 44620 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_485
timestamp 1688980957
transform 1 0 45724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_497
timestamp 1688980957
transform 1 0 46828 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_503
timestamp 1688980957
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_505
timestamp 1688980957
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_517
timestamp 1688980957
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_529
timestamp 1688980957
transform 1 0 49772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_541
timestamp 1688980957
transform 1 0 50876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_553
timestamp 1688980957
transform 1 0 51980 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_559
timestamp 1688980957
transform 1 0 52532 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_561
timestamp 1688980957
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_573
timestamp 1688980957
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_585
timestamp 1688980957
transform 1 0 54924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_597
timestamp 1688980957
transform 1 0 56028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_609
timestamp 1688980957
transform 1 0 57132 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_615
timestamp 1688980957
transform 1 0 57684 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_617
timestamp 1688980957
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_629
timestamp 1688980957
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_641
timestamp 1688980957
transform 1 0 60076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_653
timestamp 1688980957
transform 1 0 61180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_665
timestamp 1688980957
transform 1 0 62284 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_671
timestamp 1688980957
transform 1 0 62836 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_673
timestamp 1688980957
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_685
timestamp 1688980957
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_697
timestamp 1688980957
transform 1 0 65228 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_709
timestamp 1688980957
transform 1 0 66332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_721
timestamp 1688980957
transform 1 0 67436 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_727
timestamp 1688980957
transform 1 0 67988 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_729
timestamp 1688980957
transform 1 0 68172 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_3
timestamp 1688980957
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_15
timestamp 1688980957
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_27
timestamp 1688980957
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_29
timestamp 1688980957
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_41
timestamp 1688980957
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_53
timestamp 1688980957
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_65
timestamp 1688980957
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_77
timestamp 1688980957
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_83
timestamp 1688980957
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_85
timestamp 1688980957
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_97
timestamp 1688980957
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_109
timestamp 1688980957
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_121
timestamp 1688980957
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_133
timestamp 1688980957
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_139
timestamp 1688980957
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_141
timestamp 1688980957
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_153
timestamp 1688980957
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_165
timestamp 1688980957
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_177
timestamp 1688980957
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_189
timestamp 1688980957
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_195
timestamp 1688980957
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_197
timestamp 1688980957
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_209
timestamp 1688980957
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_221
timestamp 1688980957
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_233
timestamp 1688980957
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_245
timestamp 1688980957
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_251
timestamp 1688980957
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_253
timestamp 1688980957
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_265
timestamp 1688980957
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_277
timestamp 1688980957
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_289
timestamp 1688980957
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_301
timestamp 1688980957
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_307
timestamp 1688980957
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_309
timestamp 1688980957
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_321
timestamp 1688980957
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_333
timestamp 1688980957
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_345
timestamp 1688980957
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_357
timestamp 1688980957
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_363
timestamp 1688980957
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_365
timestamp 1688980957
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_377
timestamp 1688980957
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_389
timestamp 1688980957
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_401
timestamp 1688980957
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_413
timestamp 1688980957
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_419
timestamp 1688980957
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_421
timestamp 1688980957
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_433
timestamp 1688980957
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_445
timestamp 1688980957
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_457
timestamp 1688980957
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_469
timestamp 1688980957
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_475
timestamp 1688980957
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_477
timestamp 1688980957
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_489
timestamp 1688980957
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_501
timestamp 1688980957
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_513
timestamp 1688980957
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_525
timestamp 1688980957
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_531
timestamp 1688980957
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_533
timestamp 1688980957
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_545
timestamp 1688980957
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_557
timestamp 1688980957
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_569
timestamp 1688980957
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_581
timestamp 1688980957
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_587
timestamp 1688980957
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_589
timestamp 1688980957
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_601
timestamp 1688980957
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_613
timestamp 1688980957
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_625
timestamp 1688980957
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_637
timestamp 1688980957
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_643
timestamp 1688980957
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_645
timestamp 1688980957
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_657
timestamp 1688980957
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_669
timestamp 1688980957
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_681
timestamp 1688980957
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_693
timestamp 1688980957
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_699
timestamp 1688980957
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_701
timestamp 1688980957
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_713
timestamp 1688980957
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_725
timestamp 1688980957
transform 1 0 67804 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_6
timestamp 1688980957
transform 1 0 1656 0 -1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_13
timestamp 1688980957
transform 1 0 2300 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_25
timestamp 1688980957
transform 1 0 3404 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_29
timestamp 1688980957
transform 1 0 3772 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_37
timestamp 1688980957
transform 1 0 4508 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_41
timestamp 1688980957
transform 1 0 4876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_53
timestamp 1688980957
transform 1 0 5980 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_57
timestamp 1688980957
transform 1 0 6348 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_65
timestamp 1688980957
transform 1 0 7084 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_69
timestamp 1688980957
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_81
timestamp 1688980957
transform 1 0 8556 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_85
timestamp 1688980957
transform 1 0 8924 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_93
timestamp 1688980957
transform 1 0 9660 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_97
timestamp 1688980957
transform 1 0 10028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_109
timestamp 1688980957
transform 1 0 11132 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_113
timestamp 1688980957
transform 1 0 11500 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_121
timestamp 1688980957
transform 1 0 12236 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_125
timestamp 1688980957
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_137
timestamp 1688980957
transform 1 0 13708 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_141
timestamp 1688980957
transform 1 0 14076 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_149
timestamp 1688980957
transform 1 0 14812 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_153
timestamp 1688980957
transform 1 0 15180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_165
timestamp 1688980957
transform 1 0 16284 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_169
timestamp 1688980957
transform 1 0 16652 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_177
timestamp 1688980957
transform 1 0 17388 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_181
timestamp 1688980957
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_193
timestamp 1688980957
transform 1 0 18860 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_197
timestamp 1688980957
transform 1 0 19228 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_205
timestamp 1688980957
transform 1 0 19964 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_209
timestamp 1688980957
transform 1 0 20332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_221
timestamp 1688980957
transform 1 0 21436 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_225
timestamp 1688980957
transform 1 0 21804 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_233
timestamp 1688980957
transform 1 0 22540 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_237
timestamp 1688980957
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_249
timestamp 1688980957
transform 1 0 24012 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_253
timestamp 1688980957
transform 1 0 24380 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_261
timestamp 1688980957
transform 1 0 25116 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_265
timestamp 1688980957
transform 1 0 25484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_277
timestamp 1688980957
transform 1 0 26588 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_281
timestamp 1688980957
transform 1 0 26956 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_289
timestamp 1688980957
transform 1 0 27692 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_293
timestamp 1688980957
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_305
timestamp 1688980957
transform 1 0 29164 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_309
timestamp 1688980957
transform 1 0 29532 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_317
timestamp 1688980957
transform 1 0 30268 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_321
timestamp 1688980957
transform 1 0 30636 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_333
timestamp 1688980957
transform 1 0 31740 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_337
timestamp 1688980957
transform 1 0 32108 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_345
timestamp 1688980957
transform 1 0 32844 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_349
timestamp 1688980957
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_361
timestamp 1688980957
transform 1 0 34316 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_365
timestamp 1688980957
transform 1 0 34684 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_377
timestamp 1688980957
transform 1 0 35788 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_389
timestamp 1688980957
transform 1 0 36892 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_393
timestamp 1688980957
transform 1 0 37260 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_401
timestamp 1688980957
transform 1 0 37996 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_405
timestamp 1688980957
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_417
timestamp 1688980957
transform 1 0 39468 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_421
timestamp 1688980957
transform 1 0 39836 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_429
timestamp 1688980957
transform 1 0 40572 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_433
timestamp 1688980957
transform 1 0 40940 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_445
timestamp 1688980957
transform 1 0 42044 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_449
timestamp 1688980957
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_461
timestamp 1688980957
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_473
timestamp 1688980957
transform 1 0 44620 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_477
timestamp 1688980957
transform 1 0 44988 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_485
timestamp 1688980957
transform 1 0 45724 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_489
timestamp 1688980957
transform 1 0 46092 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_501
timestamp 1688980957
transform 1 0 47196 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_505
timestamp 1688980957
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_517
timestamp 1688980957
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_529
timestamp 1688980957
transform 1 0 49772 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_533
timestamp 1688980957
transform 1 0 50140 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_545
timestamp 1688980957
transform 1 0 51244 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_557
timestamp 1688980957
transform 1 0 52348 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_561
timestamp 1688980957
transform 1 0 52716 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_569
timestamp 1688980957
transform 1 0 53452 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_573
timestamp 1688980957
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_585
timestamp 1688980957
transform 1 0 54924 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_589
timestamp 1688980957
transform 1 0 55292 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_597
timestamp 1688980957
transform 1 0 56028 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_601
timestamp 1688980957
transform 1 0 56396 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_613
timestamp 1688980957
transform 1 0 57500 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_617
timestamp 1688980957
transform 1 0 57868 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_625
timestamp 1688980957
transform 1 0 58604 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_629
timestamp 1688980957
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_641
timestamp 1688980957
transform 1 0 60076 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_645
timestamp 1688980957
transform 1 0 60444 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_653
timestamp 1688980957
transform 1 0 61180 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_657
timestamp 1688980957
transform 1 0 61548 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_669
timestamp 1688980957
transform 1 0 62652 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_673
timestamp 1688980957
transform 1 0 63020 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_681
timestamp 1688980957
transform 1 0 63756 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_685
timestamp 1688980957
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_697
timestamp 1688980957
transform 1 0 65228 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_701
timestamp 1688980957
transform 1 0 65596 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_713
timestamp 1688980957
transform 1 0 66700 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_725
timestamp 1688980957
transform 1 0 67804 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_729
timestamp 1688980957
transform 1 0 68172 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37168 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 44160 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 37720 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 36984 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 30360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 31832 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 30820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 41584 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 40940 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 32200 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 39008 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 41676 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 40296 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 42228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 49220 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 28336 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 44344 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 36616 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 35604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 33856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 33396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 29440 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 38548 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 33764 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 33304 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 31188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 31004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 42780 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 38548 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 33764 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 42228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 42780 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 38640 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 43424 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 35328 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 25024 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 40572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 40388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 25944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 26680 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 45356 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 38824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 48392 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 32292 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 42412 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 41676 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 27232 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 44252 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 44988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 45724 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 35328 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 35328 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 35880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 46276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 37812 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform 1 0 37812 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 36616 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 38824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 38088 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 31372 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 25668 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 33304 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 32568 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 38640 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 31004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 30268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform 1 0 45080 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 43700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 33212 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 44068 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 35972 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 27968 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 45724 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 45448 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 51704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 50692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 32384 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 29900 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 50140 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform 1 0 43516 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 46000 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform 1 0 48484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 48760 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 37168 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 41032 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 31096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform 1 0 32108 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 31096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform 1 0 36984 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 36064 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform 1 0 39560 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 48300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform 1 0 42504 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform 1 0 45908 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 44252 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform 1 0 46000 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform 1 0 35328 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 35052 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform 1 0 34500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform 1 0 41492 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform 1 0 31096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform 1 0 42412 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform 1 0 42412 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform 1 0 53268 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform 1 0 50876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform 1 0 35696 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform 1 0 36248 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform 1 0 41308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform 1 0 31924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 32292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 52716 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform 1 0 27600 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 51152 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform 1 0 48116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform 1 0 38272 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform 1 0 39836 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform 1 0 27876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform 1 0 36800 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform 1 0 30728 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 25576 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform 1 0 50508 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform 1 0 45724 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 27600 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform 1 0 29440 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 27232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform 1 0 24840 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform 1 0 24564 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform 1 0 38640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform 1 0 24656 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform 1 0 30452 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform 1 0 40020 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 47932 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform 1 0 46644 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform 1 0 40940 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform 1 0 36248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform 1 0 27784 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1688980957
transform 1 0 68172 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1688980957
transform 1 0 48392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1688980957
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1688980957
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1688980957
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1688980957
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1688980957
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1688980957
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1688980957
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1688980957
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1688980957
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1688980957
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1688980957
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1688980957
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1688980957
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1688980957
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1688980957
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1688980957
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1688980957
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1688980957
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1688980957
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1688980957
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1688980957
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1688980957
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1688980957
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1688980957
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1688980957
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1688980957
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1688980957
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1688980957
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1688980957
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1688980957
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1688980957
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1688980957
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1688980957
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1688980957
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1688980957
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1688980957
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1688980957
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1688980957
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1688980957
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1688980957
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1688980957
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1688980957
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1688980957
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1688980957
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1688980957
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1688980957
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1688980957
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1688980957
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1688980957
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1688980957
transform -1 0 68816 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1688980957
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1688980957
transform -1 0 68816 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1688980957
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1688980957
transform -1 0 68816 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1688980957
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1688980957
transform -1 0 68816 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1688980957
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1688980957
transform -1 0 68816 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1688980957
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1688980957
transform -1 0 68816 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1688980957
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1688980957
transform -1 0 68816 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1688980957
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1688980957
transform -1 0 68816 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1688980957
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1688980957
transform -1 0 68816 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1688980957
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1688980957
transform -1 0 68816 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1688980957
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1688980957
transform -1 0 68816 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1688980957
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1688980957
transform -1 0 68816 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1688980957
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1688980957
transform -1 0 68816 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1688980957
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1688980957
transform -1 0 68816 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1688980957
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1688980957
transform -1 0 68816 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1688980957
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1688980957
transform -1 0 68816 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1688980957
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1688980957
transform -1 0 68816 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1688980957
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1688980957
transform -1 0 68816 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1688980957
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1688980957
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1688980957
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1688980957
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1688980957
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1688980957
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1688980957
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1688980957
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1688980957
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1688980957
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1688980957
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1688980957
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1688980957
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1688980957
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1688980957
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1688980957
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1688980957
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1688980957
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1688980957
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1688980957
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1688980957
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1688980957
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1688980957
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1688980957
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1688980957
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1688980957
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1688980957
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1688980957
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1688980957
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1688980957
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1688980957
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1688980957
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1688980957
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1688980957
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1688980957
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1688980957
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1688980957
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1688980957
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1688980957
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1688980957
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1688980957
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1688980957
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1688980957
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1688980957
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1688980957
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1688980957
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1688980957
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1688980957
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1688980957
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1688980957
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1688980957
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1688980957
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1688980957
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1688980957
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1688980957
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1688980957
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1688980957
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1688980957
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1688980957
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1688980957
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1688980957
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1688980957
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1688980957
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1688980957
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1688980957
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1688980957
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1688980957
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1688980957
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1688980957
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1688980957
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1688980957
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1688980957
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1688980957
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1688980957
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1688980957
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1688980957
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1688980957
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1688980957
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1688980957
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1688980957
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1688980957
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1688980957
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1688980957
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1688980957
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1688980957
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1688980957
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1688980957
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1688980957
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1688980957
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1688980957
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1688980957
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1688980957
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1688980957
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1688980957
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1688980957
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1688980957
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1688980957
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1688980957
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1688980957
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1688980957
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1688980957
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1688980957
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1688980957
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1688980957
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1688980957
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1688980957
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1688980957
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1688980957
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1688980957
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1688980957
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1688980957
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1688980957
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1688980957
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1688980957
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1688980957
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1688980957
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1688980957
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1688980957
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1688980957
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1688980957
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1688980957
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1688980957
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1688980957
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1688980957
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1688980957
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1688980957
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1688980957
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1688980957
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1688980957
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1688980957
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1688980957
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1688980957
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1688980957
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1688980957
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1688980957
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1688980957
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1688980957
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1688980957
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1688980957
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1688980957
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1688980957
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1688980957
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1688980957
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1688980957
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1688980957
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1688980957
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1688980957
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1688980957
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1688980957
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1688980957
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1688980957
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1688980957
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1688980957
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1688980957
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1688980957
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1688980957
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1688980957
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1688980957
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1688980957
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1688980957
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1688980957
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1688980957
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1688980957
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1688980957
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1688980957
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1688980957
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1688980957
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1688980957
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1688980957
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1688980957
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1688980957
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1688980957
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1688980957
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1688980957
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1688980957
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1688980957
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1688980957
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1688980957
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1688980957
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1688980957
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1688980957
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1688980957
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1688980957
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1688980957
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1688980957
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1688980957
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1688980957
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1688980957
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1688980957
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1688980957
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1688980957
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1688980957
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1688980957
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1688980957
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1688980957
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1688980957
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1688980957
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1688980957
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1688980957
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1688980957
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1688980957
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1688980957
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1688980957
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1688980957
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1688980957
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1688980957
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1688980957
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1688980957
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1688980957
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1688980957
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1688980957
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1688980957
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1688980957
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1688980957
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1688980957
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1688980957
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1688980957
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1688980957
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1688980957
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1688980957
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1688980957
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1688980957
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1688980957
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1688980957
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1688980957
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1688980957
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1688980957
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1688980957
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1688980957
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1688980957
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1688980957
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1688980957
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1688980957
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1688980957
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1688980957
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1688980957
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1688980957
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1688980957
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1688980957
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1688980957
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1688980957
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1688980957
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1688980957
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1688980957
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1688980957
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1688980957
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1688980957
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1688980957
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1688980957
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1688980957
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1688980957
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1688980957
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1688980957
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1688980957
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1688980957
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1688980957
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1688980957
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1688980957
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1688980957
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1688980957
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1688980957
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1688980957
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1688980957
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1688980957
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1688980957
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1688980957
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1688980957
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1688980957
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1688980957
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1688980957
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1688980957
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1688980957
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1688980957
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1688980957
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1688980957
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1688980957
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1688980957
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1688980957
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1688980957
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1688980957
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1688980957
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1688980957
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1688980957
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1688980957
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1688980957
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1688980957
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1688980957
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1688980957
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1688980957
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1688980957
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1688980957
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1688980957
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1688980957
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1688980957
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1688980957
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1688980957
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1688980957
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1688980957
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1688980957
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1688980957
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1688980957
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1688980957
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1688980957
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1688980957
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1688980957
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1688980957
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1688980957
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1688980957
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1688980957
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1688980957
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1688980957
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1688980957
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1688980957
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1688980957
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1688980957
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1688980957
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1688980957
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1688980957
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1688980957
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1688980957
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1688980957
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1688980957
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1688980957
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1688980957
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1688980957
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1688980957
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1688980957
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1688980957
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1688980957
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1688980957
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1688980957
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1688980957
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1688980957
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1688980957
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1688980957
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1688980957
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1688980957
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1688980957
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1688980957
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1688980957
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1688980957
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1688980957
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1688980957
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1688980957
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1688980957
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1688980957
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1688980957
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1688980957
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1688980957
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1688980957
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1688980957
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1688980957
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1688980957
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1688980957
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1688980957
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1688980957
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1688980957
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1688980957
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1688980957
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1688980957
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1688980957
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1688980957
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1688980957
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1688980957
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1688980957
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1688980957
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1688980957
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1688980957
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1688980957
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1688980957
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1688980957
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1688980957
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1688980957
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1688980957
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1688980957
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1688980957
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1688980957
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1688980957
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1688980957
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1688980957
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1688980957
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1688980957
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1688980957
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1688980957
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1688980957
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1688980957
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1688980957
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1688980957
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1688980957
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1688980957
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1688980957
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1688980957
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1688980957
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1688980957
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1688980957
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1688980957
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1688980957
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1688980957
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1688980957
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1688980957
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1688980957
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1688980957
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1688980957
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1688980957
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1688980957
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1688980957
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1688980957
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1688980957
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1688980957
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1688980957
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1688980957
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1688980957
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1688980957
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1688980957
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1688980957
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1688980957
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1688980957
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1688980957
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1688980957
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1688980957
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1688980957
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1688980957
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1688980957
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1688980957
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1688980957
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1688980957
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1688980957
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1688980957
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1688980957
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1688980957
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1688980957
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1688980957
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1688980957
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1688980957
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1688980957
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1688980957
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1688980957
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1688980957
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1688980957
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1688980957
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1688980957
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1688980957
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1688980957
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1688980957
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1688980957
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1688980957
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1688980957
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1688980957
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1688980957
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1688980957
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1688980957
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1688980957
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1688980957
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1688980957
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1688980957
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1688980957
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1688980957
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1688980957
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1688980957
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1688980957
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1688980957
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1688980957
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1688980957
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1688980957
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1688980957
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1688980957
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1688980957
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1688980957
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1688980957
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1688980957
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1688980957
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1688980957
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1688980957
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1688980957
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1688980957
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1688980957
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1688980957
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1688980957
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1688980957
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1688980957
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1688980957
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1688980957
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1688980957
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1688980957
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1688980957
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1688980957
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1688980957
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1688980957
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1688980957
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1688980957
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1688980957
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1688980957
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1688980957
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1688980957
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1688980957
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1688980957
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1688980957
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1688980957
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1688980957
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1688980957
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1688980957
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1688980957
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1688980957
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1688980957
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1688980957
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1688980957
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1688980957
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1688980957
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1688980957
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1688980957
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1688980957
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1688980957
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1688980957
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1688980957
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1688980957
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1688980957
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1688980957
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1688980957
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1688980957
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1688980957
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1688980957
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1688980957
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1688980957
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1688980957
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1688980957
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1688980957
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1688980957
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1688980957
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1688980957
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1688980957
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1688980957
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1688980957
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1688980957
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1688980957
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1688980957
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1688980957
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1688980957
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1688980957
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1688980957
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1688980957
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1688980957
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1688980957
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1688980957
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1688980957
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1688980957
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1688980957
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1688980957
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1688980957
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1688980957
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1688980957
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1688980957
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1688980957
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1688980957
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1688980957
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1688980957
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1688980957
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1688980957
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1688980957
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1688980957
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1688980957
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1688980957
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1688980957
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1688980957
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1688980957
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1688980957
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1688980957
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1688980957
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1688980957
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1688980957
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1688980957
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1688980957
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1688980957
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1688980957
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1688980957
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1688980957
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1688980957
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1688980957
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1688980957
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1688980957
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1688980957
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1688980957
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1688980957
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1688980957
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1688980957
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1688980957
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1688980957
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1688980957
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1688980957
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1688980957
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1688980957
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1688980957
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1688980957
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1688980957
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1688980957
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1688980957
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1688980957
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1688980957
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1688980957
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1688980957
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1688980957
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1688980957
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1688980957
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1688980957
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1688980957
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1688980957
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1688980957
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1688980957
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1688980957
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1688980957
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1688980957
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1688980957
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1688980957
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1688980957
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1688980957
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1688980957
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1688980957
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1688980957
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1688980957
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1688980957
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1688980957
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1688980957
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1688980957
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1688980957
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1688980957
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1688980957
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1688980957
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1688980957
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1688980957
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1688980957
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1688980957
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1688980957
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1688980957
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1688980957
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1688980957
transform 1 0 60352 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1688980957
transform 1 0 65504 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1688980957
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1688980957
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1688980957
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1688980957
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1688980957
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1688980957
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1688980957
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1688980957
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1688980957
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1688980957
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1688980957
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1688980957
transform 1 0 62928 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1688980957
transform 1 0 68080 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1688980957
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1688980957
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1688980957
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1688980957
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1688980957
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1688980957
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1688980957
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1688980957
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1688980957
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1688980957
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1688980957
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1688980957
transform 1 0 60352 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1688980957
transform 1 0 65504 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1688980957
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1688980957
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1688980957
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1688980957
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1688980957
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1688980957
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1688980957
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1688980957
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1688980957
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1688980957
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1688980957
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1688980957
transform 1 0 62928 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1688980957
transform 1 0 68080 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1688980957
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1688980957
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1688980957
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1688980957
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1688980957
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1688980957
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1688980957
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1688980957
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1688980957
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1688980957
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1688980957
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1688980957
transform 1 0 60352 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1688980957
transform 1 0 65504 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1688980957
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1688980957
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1688980957
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1688980957
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1688980957
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1688980957
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1688980957
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1688980957
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1688980957
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1688980957
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1688980957
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1688980957
transform 1 0 62928 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1688980957
transform 1 0 68080 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1688980957
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1688980957
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1688980957
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1688980957
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1688980957
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1688980957
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1688980957
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1688980957
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1688980957
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1688980957
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1688980957
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1688980957
transform 1 0 60352 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1688980957
transform 1 0 65504 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1688980957
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1688980957
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1688980957
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1688980957
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1688980957
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1688980957
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1688980957
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1688980957
transform 1 0 42320 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1688980957
transform 1 0 47472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1688980957
transform 1 0 52624 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1688980957
transform 1 0 57776 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1688980957
transform 1 0 62928 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1688980957
transform 1 0 68080 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1688980957
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1688980957
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1688980957
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1688980957
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1688980957
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1688980957
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1688980957
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1688980957
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1688980957
transform 1 0 44896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1688980957
transform 1 0 50048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1688980957
transform 1 0 55200 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1688980957
transform 1 0 60352 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1688980957
transform 1 0 65504 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1688980957
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1688980957
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1688980957
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1688980957
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1688980957
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1688980957
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1688980957
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1688980957
transform 1 0 42320 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1688980957
transform 1 0 47472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1688980957
transform 1 0 52624 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1688980957
transform 1 0 57776 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1688980957
transform 1 0 62928 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1688980957
transform 1 0 68080 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1688980957
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1688980957
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1688980957
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1688980957
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1688980957
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1688980957
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1688980957
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1688980957
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1688980957
transform 1 0 44896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1688980957
transform 1 0 50048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1688980957
transform 1 0 55200 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1688980957
transform 1 0 60352 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1688980957
transform 1 0 65504 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1688980957
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1688980957
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1688980957
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1688980957
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1688980957
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1688980957
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1688980957
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1688980957
transform 1 0 42320 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1688980957
transform 1 0 47472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1688980957
transform 1 0 52624 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1688980957
transform 1 0 57776 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1688980957
transform 1 0 62928 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1688980957
transform 1 0 68080 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1688980957
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1688980957
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1688980957
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1688980957
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1688980957
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1688980957
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1688980957
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1688980957
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1688980957
transform 1 0 44896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1688980957
transform 1 0 50048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1688980957
transform 1 0 55200 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1688980957
transform 1 0 60352 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1688980957
transform 1 0 65504 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1688980957
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1688980957
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1688980957
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1688980957
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1688980957
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1688980957
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1688980957
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1688980957
transform 1 0 42320 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1688980957
transform 1 0 47472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1688980957
transform 1 0 52624 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1688980957
transform 1 0 57776 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1688980957
transform 1 0 62928 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1688980957
transform 1 0 68080 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1688980957
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1688980957
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1688980957
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1688980957
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1688980957
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1688980957
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1688980957
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1688980957
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1688980957
transform 1 0 44896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1688980957
transform 1 0 50048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1688980957
transform 1 0 55200 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1688980957
transform 1 0 60352 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1688980957
transform 1 0 65504 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1688980957
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1688980957
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1688980957
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1688980957
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1688980957
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1688980957
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1688980957
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1688980957
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1688980957
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1688980957
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1688980957
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1688980957
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1688980957
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1688980957
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1688980957
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1688980957
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1688980957
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1688980957
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1688980957
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1688980957
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1688980957
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1688980957
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1688980957
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1688980957
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1688980957
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1688980957
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1688980957
transform 1 0 3680 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1688980957
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1688980957
transform 1 0 8832 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1688980957
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1688980957
transform 1 0 13984 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1688980957
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1688980957
transform 1 0 19136 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1688980957
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1688980957
transform 1 0 24288 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1688980957
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1688980957
transform 1 0 29440 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1688980957
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1688980957
transform 1 0 34592 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1688980957
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1688980957
transform 1 0 39744 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1688980957
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1688980957
transform 1 0 44896 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1688980957
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1688980957
transform 1 0 50048 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1688980957
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1688980957
transform 1 0 55200 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1688980957
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1688980957
transform 1 0 60352 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1688980957
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1688980957
transform 1 0 65504 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1688980957
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire6
timestamp 1688980957
transform 1 0 29624 0 1 7616
box -38 -48 314 592
<< labels >>
flabel metal2 s 18 69200 74 70000 0 FreeSans 224 90 0 0 audio_sample[0]
port 0 nsew signal input
flabel metal3 s 69200 68688 70000 68808 0 FreeSans 480 0 0 0 audio_sample[10]
port 1 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 audio_sample[11]
port 2 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 audio_sample[12]
port 3 nsew signal input
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 audio_sample[13]
port 4 nsew signal input
flabel metal2 s 43166 69200 43222 70000 0 FreeSans 224 90 0 0 audio_sample[14]
port 5 nsew signal input
flabel metal2 s 66350 69200 66406 70000 0 FreeSans 224 90 0 0 audio_sample[15]
port 6 nsew signal input
flabel metal2 s 50894 69200 50950 70000 0 FreeSans 224 90 0 0 audio_sample[1]
port 7 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 audio_sample[2]
port 8 nsew signal input
flabel metal2 s 35438 69200 35494 70000 0 FreeSans 224 90 0 0 audio_sample[3]
port 9 nsew signal input
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 audio_sample[4]
port 10 nsew signal input
flabel metal3 s 69200 38768 70000 38888 0 FreeSans 480 0 0 0 audio_sample[5]
port 11 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 audio_sample[6]
port 12 nsew signal input
flabel metal3 s 0 53728 800 53848 0 FreeSans 480 0 0 0 audio_sample[7]
port 13 nsew signal input
flabel metal2 s 48318 69200 48374 70000 0 FreeSans 224 90 0 0 audio_sample[8]
port 14 nsew signal input
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 audio_sample[9]
port 15 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal3 s 69200 60528 70000 60648 0 FreeSans 480 0 0 0 done
port 17 nsew signal tristate
flabel metal3 s 0 59168 800 59288 0 FreeSans 480 0 0 0 io_oeb[0]
port 18 nsew signal tristate
flabel metal3 s 69200 22448 70000 22568 0 FreeSans 480 0 0 0 io_oeb[10]
port 19 nsew signal tristate
flabel metal3 s 69200 57808 70000 57928 0 FreeSans 480 0 0 0 io_oeb[11]
port 20 nsew signal tristate
flabel metal2 s 58622 69200 58678 70000 0 FreeSans 224 90 0 0 io_oeb[12]
port 21 nsew signal tristate
flabel metal3 s 69200 14288 70000 14408 0 FreeSans 480 0 0 0 io_oeb[13]
port 22 nsew signal tristate
flabel metal3 s 69200 65968 70000 66088 0 FreeSans 480 0 0 0 io_oeb[14]
port 23 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 io_oeb[15]
port 24 nsew signal tristate
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 io_oeb[16]
port 25 nsew signal tristate
flabel metal3 s 69200 11568 70000 11688 0 FreeSans 480 0 0 0 io_oeb[17]
port 26 nsew signal tristate
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 io_oeb[18]
port 27 nsew signal tristate
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 io_oeb[19]
port 28 nsew signal tristate
flabel metal2 s 19982 69200 20038 70000 0 FreeSans 224 90 0 0 io_oeb[1]
port 29 nsew signal tristate
flabel metal2 s 38014 69200 38070 70000 0 FreeSans 224 90 0 0 io_oeb[20]
port 30 nsew signal tristate
flabel metal2 s 63774 69200 63830 70000 0 FreeSans 224 90 0 0 io_oeb[21]
port 31 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 32 nsew signal tristate
flabel metal3 s 69200 52368 70000 52488 0 FreeSans 480 0 0 0 io_oeb[23]
port 33 nsew signal tristate
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_oeb[24]
port 34 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 io_oeb[25]
port 35 nsew signal tristate
flabel metal3 s 69200 3408 70000 3528 0 FreeSans 480 0 0 0 io_oeb[26]
port 36 nsew signal tristate
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 37 nsew signal tristate
flabel metal3 s 69200 30608 70000 30728 0 FreeSans 480 0 0 0 io_oeb[28]
port 38 nsew signal tristate
flabel metal3 s 69200 25168 70000 25288 0 FreeSans 480 0 0 0 io_oeb[29]
port 39 nsew signal tristate
flabel metal2 s 22558 69200 22614 70000 0 FreeSans 224 90 0 0 io_oeb[2]
port 40 nsew signal tristate
flabel metal2 s 25134 69200 25190 70000 0 FreeSans 224 90 0 0 io_oeb[30]
port 41 nsew signal tristate
flabel metal3 s 69200 55088 70000 55208 0 FreeSans 480 0 0 0 io_oeb[31]
port 42 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 io_oeb[32]
port 43 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 44 nsew signal tristate
flabel metal3 s 69200 8848 70000 8968 0 FreeSans 480 0 0 0 io_oeb[34]
port 45 nsew signal tristate
flabel metal3 s 69200 688 70000 808 0 FreeSans 480 0 0 0 io_oeb[35]
port 46 nsew signal tristate
flabel metal3 s 69200 36048 70000 36168 0 FreeSans 480 0 0 0 io_oeb[36]
port 47 nsew signal tristate
flabel metal3 s 0 51008 800 51128 0 FreeSans 480 0 0 0 io_oeb[37]
port 48 nsew signal tristate
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 49 nsew signal tristate
flabel metal2 s 27710 69200 27766 70000 0 FreeSans 224 90 0 0 io_oeb[4]
port 50 nsew signal tristate
flabel metal3 s 69200 63248 70000 63368 0 FreeSans 480 0 0 0 io_oeb[5]
port 51 nsew signal tristate
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 52 nsew signal tristate
flabel metal2 s 32862 69200 32918 70000 0 FreeSans 224 90 0 0 io_oeb[7]
port 53 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 54 nsew signal tristate
flabel metal3 s 69200 17008 70000 17128 0 FreeSans 480 0 0 0 io_oeb[9]
port 55 nsew signal tristate
flabel metal3 s 69200 44208 70000 44328 0 FreeSans 480 0 0 0 io_out[0]
port 56 nsew signal tristate
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 io_out[10]
port 57 nsew signal tristate
flabel metal2 s 40590 69200 40646 70000 0 FreeSans 224 90 0 0 io_out[11]
port 58 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 io_out[12]
port 59 nsew signal tristate
flabel metal2 s 17406 69200 17462 70000 0 FreeSans 224 90 0 0 io_out[13]
port 60 nsew signal tristate
flabel metal3 s 0 64608 800 64728 0 FreeSans 480 0 0 0 io_out[14]
port 61 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 io_out[15]
port 62 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 io_out[16]
port 63 nsew signal tristate
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 io_out[17]
port 64 nsew signal tristate
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 io_out[18]
port 65 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 io_out[19]
port 66 nsew signal tristate
flabel metal3 s 69200 19728 70000 19848 0 FreeSans 480 0 0 0 io_out[1]
port 67 nsew signal tristate
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 io_out[20]
port 68 nsew signal tristate
flabel metal3 s 0 56448 800 56568 0 FreeSans 480 0 0 0 io_out[21]
port 69 nsew signal tristate
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 io_out[22]
port 70 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_out[23]
port 71 nsew signal tristate
flabel metal3 s 69200 27888 70000 28008 0 FreeSans 480 0 0 0 io_out[24]
port 72 nsew signal tristate
flabel metal3 s 69200 46928 70000 47048 0 FreeSans 480 0 0 0 io_out[25]
port 73 nsew signal tristate
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 io_out[26]
port 74 nsew signal tristate
flabel metal3 s 69200 49648 70000 49768 0 FreeSans 480 0 0 0 io_out[27]
port 75 nsew signal tristate
flabel metal2 s 7102 69200 7158 70000 0 FreeSans 224 90 0 0 io_out[28]
port 76 nsew signal tristate
flabel metal2 s 9678 69200 9734 70000 0 FreeSans 224 90 0 0 io_out[29]
port 77 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 io_out[2]
port 78 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 io_out[30]
port 79 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 io_out[31]
port 80 nsew signal tristate
flabel metal2 s 12254 69200 12310 70000 0 FreeSans 224 90 0 0 io_out[32]
port 81 nsew signal tristate
flabel metal2 s 30286 69200 30342 70000 0 FreeSans 224 90 0 0 io_out[33]
port 82 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 io_out[34]
port 83 nsew signal tristate
flabel metal3 s 0 67328 800 67448 0 FreeSans 480 0 0 0 io_out[35]
port 84 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 io_out[36]
port 85 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 io_out[37]
port 86 nsew signal tristate
flabel metal2 s 61198 69200 61254 70000 0 FreeSans 224 90 0 0 io_out[3]
port 87 nsew signal tristate
flabel metal2 s 45742 69200 45798 70000 0 FreeSans 224 90 0 0 io_out[4]
port 88 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 io_out[5]
port 89 nsew signal tristate
flabel metal2 s 68926 69200 68982 70000 0 FreeSans 224 90 0 0 io_out[6]
port 90 nsew signal tristate
flabel metal3 s 69200 6128 70000 6248 0 FreeSans 480 0 0 0 io_out[7]
port 91 nsew signal tristate
flabel metal2 s 1950 69200 2006 70000 0 FreeSans 224 90 0 0 io_out[8]
port 92 nsew signal tristate
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 io_out[9]
port 93 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 psram_ce_n
port 94 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 psram_d[0]
port 95 nsew signal bidirectional
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 psram_d[1]
port 96 nsew signal bidirectional
flabel metal3 s 69200 41488 70000 41608 0 FreeSans 480 0 0 0 psram_d[2]
port 97 nsew signal bidirectional
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 psram_d[3]
port 98 nsew signal bidirectional
flabel metal2 s 56046 69200 56102 70000 0 FreeSans 224 90 0 0 psram_douten[0]
port 99 nsew signal tristate
flabel metal2 s 53470 69200 53526 70000 0 FreeSans 224 90 0 0 psram_douten[1]
port 100 nsew signal tristate
flabel metal2 s 4526 69200 4582 70000 0 FreeSans 224 90 0 0 psram_douten[2]
port 101 nsew signal tristate
flabel metal2 s 14830 69200 14886 70000 0 FreeSans 224 90 0 0 psram_douten[3]
port 102 nsew signal tristate
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 psram_sck
port 103 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 rst
port 104 nsew signal input
flabel metal3 s 0 61888 800 62008 0 FreeSans 480 0 0 0 sample_valid
port 105 nsew signal input
flabel metal3 s 69200 33328 70000 33448 0 FreeSans 480 0 0 0 start
port 106 nsew signal input
flabel metal4 s 4208 2128 4528 67504 0 FreeSans 1920 90 0 0 vccd1
port 107 nsew power bidirectional
flabel metal4 s 34928 2128 35248 67504 0 FreeSans 1920 90 0 0 vccd1
port 107 nsew power bidirectional
flabel metal4 s 65648 2128 65968 67504 0 FreeSans 1920 90 0 0 vccd1
port 107 nsew power bidirectional
flabel metal4 s 19568 2128 19888 67504 0 FreeSans 1920 90 0 0 vssd1
port 108 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 67504 0 FreeSans 1920 90 0 0 vssd1
port 108 nsew ground bidirectional
rlabel via1 34960 66912 34960 66912 0 vccd1
rlabel metal1 34960 67456 34960 67456 0 vssd1
rlabel metal2 33166 14790 33166 14790 0 _0000_
rlabel metal1 33023 13906 33023 13906 0 _0001_
rlabel metal1 29654 15062 29654 15062 0 _0002_
rlabel metal1 28791 17170 28791 17170 0 _0003_
rlabel metal2 37674 13090 37674 13090 0 _0004_
rlabel metal1 38175 11730 38175 11730 0 _0005_
rlabel metal1 41331 12954 41331 12954 0 _0006_
rlabel metal1 40112 10506 40112 10506 0 _0007_
rlabel metal1 40556 15402 40556 15402 0 _0008_
rlabel metal1 40326 16490 40326 16490 0 _0009_
rlabel metal1 34679 19414 34679 19414 0 _0010_
rlabel metal2 32614 20774 32614 20774 0 _0011_
rlabel metal1 33023 15402 33023 15402 0 _0012_
rlabel metal1 29716 13498 29716 13498 0 _0013_
rlabel metal1 32568 11730 32568 11730 0 _0014_
rlabel metal1 33856 12750 33856 12750 0 _0015_
rlabel metal2 31050 14756 31050 14756 0 _0016_
rlabel metal1 29348 15674 29348 15674 0 _0017_
rlabel via1 25801 16558 25801 16558 0 _0018_
rlabel metal1 30171 16558 30171 16558 0 _0019_
rlabel metal2 36478 14790 36478 14790 0 _0020_
rlabel metal1 35144 11866 35144 11866 0 _0021_
rlabel metal1 37076 11186 37076 11186 0 _0022_
rlabel metal1 36064 12750 36064 12750 0 _0023_
rlabel metal1 39606 13430 39606 13430 0 _0024_
rlabel metal1 39192 11322 39192 11322 0 _0025_
rlabel metal1 40567 9622 40567 9622 0 _0026_
rlabel metal1 40434 12716 40434 12716 0 _0027_
rlabel metal1 42550 15130 42550 15130 0 _0028_
rlabel metal1 39376 15674 39376 15674 0 _0029_
rlabel metal1 39688 17170 39688 17170 0 _0030_
rlabel metal1 36386 18938 36386 18938 0 _0031_
rlabel metal1 35558 21896 35558 21896 0 _0032_
rlabel metal2 33350 20604 33350 20604 0 _0033_
rlabel metal1 29164 21114 29164 21114 0 _0034_
rlabel metal1 29072 19482 29072 19482 0 _0035_
rlabel metal1 42591 20842 42591 20842 0 _0036_
rlabel metal1 37244 13974 37244 13974 0 _0037_
rlabel metal1 33529 11798 33529 11798 0 _0038_
rlabel metal1 42959 13974 42959 13974 0 _0039_
rlabel metal1 40429 19822 40429 19822 0 _0040_
rlabel metal1 41068 13906 41068 13906 0 _0041_
rlabel metal1 34776 14586 34776 14586 0 _0042_
rlabel metal1 43976 16218 43976 16218 0 _0043_
rlabel metal2 31970 7684 31970 7684 0 _0044_
rlabel metal2 30958 9894 30958 9894 0 _0045_
rlabel metal1 37904 8602 37904 8602 0 _0046_
rlabel metal2 43378 9860 43378 9860 0 _0047_
rlabel metal1 44390 13362 44390 13362 0 _0048_
rlabel metal1 43516 15538 43516 15538 0 _0049_
rlabel via2 39238 15419 39238 15419 0 _0050_
rlabel metal2 38134 15912 38134 15912 0 _0051_
rlabel via2 38226 16507 38226 16507 0 _0052_
rlabel metal2 33350 8024 33350 8024 0 _0053_
rlabel metal1 32292 3162 32292 3162 0 _0054_
rlabel metal1 33120 4046 33120 4046 0 _0055_
rlabel metal2 30406 2856 30406 2856 0 _0056_
rlabel metal1 28520 2618 28520 2618 0 _0057_
rlabel metal2 27094 4386 27094 4386 0 _0058_
rlabel metal1 26496 5338 26496 5338 0 _0059_
rlabel metal1 26680 6426 26680 6426 0 _0060_
rlabel metal2 29302 7650 29302 7650 0 _0061_
rlabel metal1 31648 7514 31648 7514 0 _0062_
rlabel metal2 32246 9758 32246 9758 0 _0063_
rlabel metal2 23966 13736 23966 13736 0 _0064_
rlabel metal1 26588 12410 26588 12410 0 _0065_
rlabel metal2 23690 12648 23690 12648 0 _0066_
rlabel metal1 23644 10778 23644 10778 0 _0067_
rlabel metal1 23644 9146 23644 9146 0 _0068_
rlabel metal2 24518 8296 24518 8296 0 _0069_
rlabel metal2 26358 7650 26358 7650 0 _0070_
rlabel metal1 29401 8874 29401 8874 0 _0071_
rlabel metal1 30820 9486 30820 9486 0 _0072_
rlabel metal2 33810 6494 33810 6494 0 _0073_
rlabel metal1 38456 8602 38456 8602 0 _0074_
rlabel metal1 36340 2618 36340 2618 0 _0075_
rlabel metal1 35282 4794 35282 4794 0 _0076_
rlabel metal2 34822 3944 34822 3944 0 _0077_
rlabel metal1 38502 2618 38502 2618 0 _0078_
rlabel metal1 41446 3577 41446 3577 0 _0079_
rlabel metal2 40710 2856 40710 2856 0 _0080_
rlabel metal1 42879 4522 42879 4522 0 _0081_
rlabel metal1 43431 5610 43431 5610 0 _0082_
rlabel metal1 40158 7480 40158 7480 0 _0083_
rlabel metal2 34454 9384 34454 9384 0 _0084_
rlabel metal1 43976 9622 43976 9622 0 _0085_
rlabel metal2 44482 5032 44482 5032 0 _0086_
rlabel metal1 48859 5610 48859 5610 0 _0087_
rlabel metal1 47065 4590 47065 4590 0 _0088_
rlabel metal2 44298 6562 44298 6562 0 _0089_
rlabel metal2 48806 6562 48806 6562 0 _0090_
rlabel metal1 51297 8534 51297 8534 0 _0091_
rlabel metal2 47334 9112 47334 9112 0 _0092_
rlabel metal1 50975 9622 50975 9622 0 _0093_
rlabel metal1 44811 8534 44811 8534 0 _0094_
rlabel metal2 40710 8738 40710 8738 0 _0095_
rlabel metal2 44574 13090 44574 13090 0 _0096_
rlabel metal2 47794 11526 47794 11526 0 _0097_
rlabel metal2 47150 12002 47150 12002 0 _0098_
rlabel metal2 51474 10914 51474 10914 0 _0099_
rlabel metal1 50975 10710 50975 10710 0 _0100_
rlabel metal2 53590 13090 53590 13090 0 _0101_
rlabel metal2 49910 15198 49910 15198 0 _0102_
rlabel metal2 51474 16286 51474 16286 0 _0103_
rlabel metal1 53176 14586 53176 14586 0 _0104_
rlabel metal1 49963 17238 49963 17238 0 _0105_
rlabel metal1 44857 12138 44857 12138 0 _0106_
rlabel metal1 44482 15130 44482 15130 0 _0107_
rlabel metal2 51106 18054 51106 18054 0 _0108_
rlabel metal1 49036 18598 49036 18598 0 _0109_
rlabel metal2 51106 19346 51106 19346 0 _0110_
rlabel metal2 49818 21726 49818 21726 0 _0111_
rlabel metal1 49411 23018 49411 23018 0 _0112_
rlabel metal2 45126 22814 45126 22814 0 _0113_
rlabel metal2 44574 21352 44574 21352 0 _0114_
rlabel metal2 46966 23290 46966 23290 0 _0115_
rlabel metal2 43562 20264 43562 20264 0 _0116_
rlabel metal1 38405 21998 38405 21998 0 _0117_
rlabel metal1 39958 20842 39958 20842 0 _0118_
rlabel metal1 37612 19754 37612 19754 0 _0119_
rlabel metal2 35834 18054 35834 18054 0 _0120_
rlabel metal1 37388 17646 37388 17646 0 _0121_
rlabel metal1 38824 17102 38824 17102 0 _0122_
rlabel metal1 34587 22610 34587 22610 0 _0123_
rlabel metal1 36156 23834 36156 23834 0 _0124_
rlabel metal1 34638 23630 34638 23630 0 _0125_
rlabel metal2 37766 23698 37766 23698 0 _0126_
rlabel metal1 39095 23698 39095 23698 0 _0127_
rlabel via1 35645 16558 35645 16558 0 _0128_
rlabel metal1 31786 19244 31786 19244 0 _0129_
rlabel metal1 31183 17646 31183 17646 0 _0130_
rlabel metal1 32798 17714 32798 17714 0 _0131_
rlabel via1 33989 17170 33989 17170 0 _0132_
rlabel metal1 46230 15538 46230 15538 0 _0133_
rlabel metal1 46736 14382 46736 14382 0 _0134_
rlabel metal1 33488 19958 33488 19958 0 _0135_
rlabel metal1 30636 20026 30636 20026 0 _0136_
rlabel metal1 30360 23834 30360 23834 0 _0137_
rlabel metal2 31326 23936 31326 23936 0 _0138_
rlabel via1 32701 23018 32701 23018 0 _0139_
rlabel via1 30493 21998 30493 21998 0 _0140_
rlabel metal1 28653 24854 28653 24854 0 _0141_
rlabel metal1 26951 23018 26951 23018 0 _0142_
rlabel metal1 30360 18122 30360 18122 0 _0143_
rlabel metal1 27319 17578 27319 17578 0 _0144_
rlabel metal1 26077 18734 26077 18734 0 _0145_
rlabel metal1 25622 20978 25622 20978 0 _0146_
rlabel metal1 26353 21522 26353 21522 0 _0147_
rlabel metal1 45678 12954 45678 12954 0 _0148_
rlabel metal1 44834 19754 44834 19754 0 _0149_
rlabel metal1 45034 16626 45034 16626 0 _0150_
rlabel metal1 31086 3706 31086 3706 0 _0151_
rlabel metal2 32154 5372 32154 5372 0 _0152_
rlabel metal1 29762 3094 29762 3094 0 _0153_
rlabel metal1 27784 3094 27784 3094 0 _0154_
rlabel metal1 26581 4794 26581 4794 0 _0155_
rlabel metal1 25852 5338 25852 5338 0 _0156_
rlabel metal1 27547 6970 27547 6970 0 _0157_
rlabel metal1 28428 7514 28428 7514 0 _0158_
rlabel metal1 30953 8942 30953 8942 0 _0159_
rlabel metal1 30268 12954 30268 12954 0 _0160_
rlabel metal1 23322 13498 23322 13498 0 _0161_
rlabel metal1 25898 11866 25898 11866 0 _0162_
rlabel metal1 23736 12750 23736 12750 0 _0163_
rlabel metal2 24426 10982 24426 10982 0 _0164_
rlabel metal1 23184 9486 23184 9486 0 _0165_
rlabel metal2 23506 8942 23506 8942 0 _0166_
rlabel metal1 25622 7752 25622 7752 0 _0167_
rlabel metal1 27830 9010 27830 9010 0 _0168_
rlabel via1 27825 12818 27825 12818 0 _0169_
rlabel metal1 29210 14382 29210 14382 0 _0170_
rlabel metal1 29516 11798 29516 11798 0 _0171_
rlabel metal2 33074 6052 33074 6052 0 _0172_
rlabel metal1 35512 2618 35512 2618 0 _0173_
rlabel metal2 36110 4964 36110 4964 0 _0174_
rlabel metal1 35052 4046 35052 4046 0 _0175_
rlabel metal2 37582 3434 37582 3434 0 _0176_
rlabel metal1 40388 3434 40388 3434 0 _0177_
rlabel metal1 39836 2618 39836 2618 0 _0178_
rlabel metal1 40802 4726 40802 4726 0 _0179_
rlabel metal2 41998 5474 41998 5474 0 _0180_
rlabel via1 36657 7854 36657 7854 0 _0181_
rlabel metal2 36110 9316 36110 9316 0 _0182_
rlabel metal2 33074 9758 33074 9758 0 _0183_
rlabel metal1 26307 15062 26307 15062 0 _0184_
rlabel metal1 24467 14994 24467 14994 0 _0185_
rlabel metal1 43884 4794 43884 4794 0 _0186_
rlabel metal2 47426 5916 47426 5916 0 _0187_
rlabel metal1 45901 4794 45901 4794 0 _0188_
rlabel metal1 44153 6970 44153 6970 0 _0189_
rlabel metal1 48707 6970 48707 6970 0 _0190_
rlabel metal1 49726 8058 49726 8058 0 _0191_
rlabel metal1 47189 9146 47189 9146 0 _0192_
rlabel metal2 49174 9248 49174 9248 0 _0193_
rlabel metal2 41998 8670 41998 8670 0 _0194_
rlabel metal1 42182 10234 42182 10234 0 _0195_
rlabel metal1 39596 9146 39596 9146 0 _0196_
rlabel metal2 34730 8262 34730 8262 0 _0197_
rlabel viali 35101 7718 35101 7718 0 _0198_
rlabel metal1 47610 11322 47610 11322 0 _0199_
rlabel metal1 47472 13158 47472 13158 0 _0200_
rlabel metal2 51290 11424 51290 11424 0 _0201_
rlabel metal2 49542 11118 49542 11118 0 _0202_
rlabel metal1 52118 13226 52118 13226 0 _0203_
rlabel metal1 49358 14586 49358 14586 0 _0204_
rlabel metal1 51152 15470 51152 15470 0 _0205_
rlabel metal1 52900 14926 52900 14926 0 _0206_
rlabel metal1 46184 16626 46184 16626 0 _0207_
rlabel metal1 43792 11866 43792 11866 0 _0208_
rlabel via1 41165 7378 41165 7378 0 _0209_
rlabel metal1 42632 7378 42632 7378 0 _0210_
rlabel metal1 49634 17850 49634 17850 0 _0211_
rlabel metal1 47702 18190 47702 18190 0 _0212_
rlabel metal1 49910 19890 49910 19890 0 _0213_
rlabel metal1 49312 21114 49312 21114 0 _0214_
rlabel metal1 47932 22202 47932 22202 0 _0215_
rlabel metal1 44528 22202 44528 22202 0 _0216_
rlabel metal1 45908 21454 45908 21454 0 _0217_
rlabel metal1 46552 23630 46552 23630 0 _0218_
rlabel metal1 41124 18394 41124 18394 0 _0219_
rlabel metal1 42678 18258 42678 18258 0 _0220_
rlabel metal1 45678 18190 45678 18190 0 _0221_
rlabel metal1 42458 6698 42458 6698 0 _0222_
rlabel metal2 41170 18598 41170 18598 0 _0223_
rlabel metal1 44666 18802 44666 18802 0 _0224_
rlabel metal2 46966 20502 46966 20502 0 _0225_
rlabel metal1 47518 19754 47518 19754 0 _0226_
rlabel metal1 46552 18734 46552 18734 0 _0227_
rlabel viali 43838 19333 43838 19333 0 _0228_
rlabel metal1 46460 19346 46460 19346 0 _0229_
rlabel metal1 48898 21522 48898 21522 0 _0230_
rlabel metal1 47886 21522 47886 21522 0 _0231_
rlabel metal1 46414 21930 46414 21930 0 _0232_
rlabel via1 46506 21437 46506 21437 0 _0233_
rlabel metal1 50255 19754 50255 19754 0 _0234_
rlabel viali 46703 21522 46703 21522 0 _0235_
rlabel metal1 46782 22406 46782 22406 0 _0236_
rlabel metal1 48254 21658 48254 21658 0 _0237_
rlabel metal2 47104 21658 47104 21658 0 _0238_
rlabel metal2 49726 19244 49726 19244 0 _0239_
rlabel metal2 47334 22440 47334 22440 0 _0240_
rlabel metal2 44850 22039 44850 22039 0 _0241_
rlabel metal1 48070 21964 48070 21964 0 _0242_
rlabel metal1 49542 20944 49542 20944 0 _0243_
rlabel viali 49450 20911 49450 20911 0 _0244_
rlabel metal2 49634 20026 49634 20026 0 _0245_
rlabel metal2 50186 19584 50186 19584 0 _0246_
rlabel metal1 47104 18258 47104 18258 0 _0247_
rlabel metal2 46782 18411 46782 18411 0 _0248_
rlabel metal1 49818 17646 49818 17646 0 _0249_
rlabel metal1 44666 11628 44666 11628 0 _0250_
rlabel metal1 44850 11526 44850 11526 0 _0251_
rlabel metal1 46460 8466 46460 8466 0 _0252_
rlabel metal1 46744 7786 46744 7786 0 _0253_
rlabel metal2 46506 9724 46506 9724 0 _0254_
rlabel metal1 45954 9622 45954 9622 0 _0255_
rlabel metal2 46782 9520 46782 9520 0 _0256_
rlabel metal1 40066 12954 40066 12954 0 _0257_
rlabel metal1 49634 13702 49634 13702 0 _0258_
rlabel metal2 51290 14110 51290 14110 0 _0259_
rlabel metal1 50278 13770 50278 13770 0 _0260_
rlabel metal1 40296 15470 40296 15470 0 _0261_
rlabel metal1 51750 14348 51750 14348 0 _0262_
rlabel metal1 50976 12070 50976 12070 0 _0263_
rlabel metal1 51658 13192 51658 13192 0 _0264_
rlabel metal1 51520 14382 51520 14382 0 _0265_
rlabel metal1 51658 14824 51658 14824 0 _0266_
rlabel metal1 52394 15368 52394 15368 0 _0267_
rlabel metal1 52164 12818 52164 12818 0 _0268_
rlabel metal1 52279 15470 52279 15470 0 _0269_
rlabel metal1 51934 14960 51934 14960 0 _0270_
rlabel metal2 51796 12716 51796 12716 0 _0271_
rlabel metal1 52210 14042 52210 14042 0 _0272_
rlabel metal1 51704 13294 51704 13294 0 _0273_
rlabel metal1 51566 13328 51566 13328 0 _0274_
rlabel metal1 50232 14042 50232 14042 0 _0275_
rlabel metal1 49818 11662 49818 11662 0 _0276_
rlabel metal1 49726 11764 49726 11764 0 _0277_
rlabel metal2 51566 11679 51566 11679 0 _0278_
rlabel metal1 51474 11696 51474 11696 0 _0279_
rlabel metal1 48530 13260 48530 13260 0 _0280_
rlabel metal1 47518 11152 47518 11152 0 _0281_
rlabel metal1 39192 9486 39192 9486 0 _0282_
rlabel metal1 39698 9350 39698 9350 0 _0283_
rlabel metal1 39054 5814 39054 5814 0 _0284_
rlabel metal1 39744 6086 39744 6086 0 _0285_
rlabel metal1 37858 5678 37858 5678 0 _0286_
rlabel metal1 38318 5746 38318 5746 0 _0287_
rlabel metal1 39008 5882 39008 5882 0 _0288_
rlabel metal1 37904 8466 37904 8466 0 _0289_
rlabel metal1 45724 8942 45724 8942 0 _0290_
rlabel metal1 48346 5270 48346 5270 0 _0291_
rlabel metal1 48438 8024 48438 8024 0 _0292_
rlabel metal2 47978 9078 47978 9078 0 _0293_
rlabel metal1 48622 8976 48622 8976 0 _0294_
rlabel metal1 48806 9078 48806 9078 0 _0295_
rlabel metal1 48024 7378 48024 7378 0 _0296_
rlabel metal2 48990 9282 48990 9282 0 _0297_
rlabel metal2 48806 8772 48806 8772 0 _0298_
rlabel via1 48446 7786 48446 7786 0 _0299_
rlabel metal1 49450 7514 49450 7514 0 _0300_
rlabel metal2 45402 7752 45402 7752 0 _0301_
rlabel metal1 48898 7786 48898 7786 0 _0302_
rlabel metal1 49818 7922 49818 7922 0 _0303_
rlabel metal1 48944 7378 48944 7378 0 _0304_
rlabel metal1 45448 6766 45448 6766 0 _0305_
rlabel metal1 45218 6698 45218 6698 0 _0306_
rlabel metal1 46414 5100 46414 5100 0 _0307_
rlabel metal1 46322 5236 46322 5236 0 _0308_
rlabel metal1 46736 6358 46736 6358 0 _0309_
rlabel metal1 44206 4666 44206 4666 0 _0310_
rlabel metal2 33534 10234 33534 10234 0 _0311_
rlabel metal1 33350 10234 33350 10234 0 _0312_
rlabel metal1 26818 11866 26818 11866 0 _0313_
rlabel metal1 28152 10982 28152 10982 0 _0314_
rlabel metal2 27370 10948 27370 10948 0 _0315_
rlabel metal1 28198 11050 28198 11050 0 _0316_
rlabel metal1 27462 11050 27462 11050 0 _0317_
rlabel metal1 27876 11322 27876 11322 0 _0318_
rlabel metal1 32798 9928 32798 9928 0 _0319_
rlabel metal1 40296 6698 40296 6698 0 _0320_
rlabel metal1 39422 4148 39422 4148 0 _0321_
rlabel metal1 39468 4250 39468 4250 0 _0322_
rlabel metal1 40112 5882 40112 5882 0 _0323_
rlabel metal1 40480 5678 40480 5678 0 _0324_
rlabel metal1 40848 6358 40848 6358 0 _0325_
rlabel metal1 39146 2448 39146 2448 0 _0326_
rlabel metal2 40250 6154 40250 6154 0 _0327_
rlabel metal2 41262 5712 41262 5712 0 _0328_
rlabel metal2 41538 5814 41538 5814 0 _0329_
rlabel metal2 40986 5372 40986 5372 0 _0330_
rlabel metal2 39054 4352 39054 4352 0 _0331_
rlabel metal1 40250 4522 40250 4522 0 _0332_
rlabel metal1 39836 2414 39836 2414 0 _0333_
rlabel metal1 39284 2346 39284 2346 0 _0334_
rlabel metal1 38042 3706 38042 3706 0 _0335_
rlabel metal1 36248 5270 36248 5270 0 _0336_
rlabel metal1 36294 4658 36294 4658 0 _0337_
rlabel metal1 36202 4216 36202 4216 0 _0338_
rlabel metal1 36064 4114 36064 4114 0 _0339_
rlabel metal1 36386 4624 36386 4624 0 _0340_
rlabel metal1 35880 2414 35880 2414 0 _0341_
rlabel metal1 33626 5746 33626 5746 0 _0342_
rlabel metal1 33580 5882 33580 5882 0 _0343_
rlabel metal2 31970 5610 31970 5610 0 _0344_
rlabel metal1 29670 6256 29670 6256 0 _0345_
rlabel metal1 31142 5814 31142 5814 0 _0346_
rlabel metal1 30590 5610 30590 5610 0 _0347_
rlabel metal1 31326 5202 31326 5202 0 _0348_
rlabel metal1 32338 13328 32338 13328 0 _0349_
rlabel metal1 27324 10030 27324 10030 0 _0350_
rlabel metal2 25714 11254 25714 11254 0 _0351_
rlabel metal1 26312 9418 26312 9418 0 _0352_
rlabel metal1 26956 9622 26956 9622 0 _0353_
rlabel metal1 27232 8942 27232 8942 0 _0354_
rlabel metal1 26772 10030 26772 10030 0 _0355_
rlabel metal1 25024 12818 25024 12818 0 _0356_
rlabel metal1 25139 12138 25139 12138 0 _0357_
rlabel metal1 26772 8874 26772 8874 0 _0358_
rlabel metal2 26818 9316 26818 9316 0 _0359_
rlabel metal1 26312 8466 26312 8466 0 _0360_
rlabel metal1 26036 10030 26036 10030 0 _0361_
rlabel metal2 24886 9758 24886 9758 0 _0362_
rlabel metal1 25024 9622 25024 9622 0 _0363_
rlabel metal1 26174 10778 26174 10778 0 _0364_
rlabel metal1 23966 10098 23966 10098 0 _0365_
rlabel metal1 24794 10710 24794 10710 0 _0366_
rlabel metal1 24656 10642 24656 10642 0 _0367_
rlabel metal1 24886 12206 24886 12206 0 _0368_
rlabel metal1 27002 12308 27002 12308 0 _0369_
rlabel viali 26174 11729 26174 11729 0 _0370_
rlabel metal1 24196 12954 24196 12954 0 _0371_
rlabel metal1 28980 3502 28980 3502 0 _0372_
rlabel metal1 28290 3434 28290 3434 0 _0373_
rlabel metal2 28934 5712 28934 5712 0 _0374_
rlabel metal1 29164 6426 29164 6426 0 _0375_
rlabel metal2 31786 6596 31786 6596 0 _0376_
rlabel metal1 32292 6630 32292 6630 0 _0377_
rlabel metal1 28014 6358 28014 6358 0 _0378_
rlabel metal1 28842 6800 28842 6800 0 _0379_
rlabel metal1 29118 7344 29118 7344 0 _0380_
rlabel metal1 28704 5542 28704 5542 0 _0381_
rlabel metal1 27922 5610 27922 5610 0 _0382_
rlabel metal2 31602 4352 31602 4352 0 _0383_
rlabel metal1 27968 5202 27968 5202 0 _0384_
rlabel metal1 26174 5236 26174 5236 0 _0385_
rlabel via2 29486 5355 29486 5355 0 _0386_
rlabel metal1 27278 5134 27278 5134 0 _0387_
rlabel metal1 28382 3570 28382 3570 0 _0388_
rlabel metal2 30130 3910 30130 3910 0 _0389_
rlabel metal1 30544 4794 30544 4794 0 _0390_
rlabel metal1 32660 5338 32660 5338 0 _0391_
rlabel metal1 30866 3162 30866 3162 0 _0392_
rlabel metal1 45310 15130 45310 15130 0 _0393_
rlabel metal1 45310 16524 45310 16524 0 _0394_
rlabel metal1 44896 18598 44896 18598 0 _0395_
rlabel metal1 46276 12818 46276 12818 0 _0396_
rlabel metal1 46184 12750 46184 12750 0 _0397_
rlabel metal2 35374 14756 35374 14756 0 _0398_
rlabel metal1 31878 24171 31878 24171 0 _0399_
rlabel metal1 39606 14552 39606 14552 0 _0400_
rlabel metal1 33074 20264 33074 20264 0 _0401_
rlabel metal1 35374 22066 35374 22066 0 _0402_
rlabel metal1 39606 16728 39606 16728 0 _0403_
rlabel metal1 39284 15470 39284 15470 0 _0404_
rlabel metal1 32039 16082 32039 16082 0 _0405_
rlabel metal1 32154 16218 32154 16218 0 _0406_
rlabel metal1 34132 14926 34132 14926 0 _0407_
rlabel metal1 45494 14518 45494 14518 0 _0408_
rlabel metal1 34684 12818 34684 12818 0 _0409_
rlabel metal2 40158 13804 40158 13804 0 _0410_
rlabel metal1 37030 14926 37030 14926 0 _0411_
rlabel metal2 40894 20196 40894 20196 0 _0412_
rlabel metal1 42504 16558 42504 16558 0 _0413_
rlabel metal1 43746 16082 43746 16082 0 _0414_
rlabel metal1 34316 14314 34316 14314 0 _0415_
rlabel metal1 34868 14042 34868 14042 0 _0416_
rlabel metal1 39882 13430 39882 13430 0 _0417_
rlabel metal1 41492 20026 41492 20026 0 _0418_
rlabel metal1 40710 20468 40710 20468 0 _0419_
rlabel metal2 42918 14382 42918 14382 0 _0420_
rlabel metal1 36064 17170 36064 17170 0 _0421_
rlabel metal1 33994 14790 33994 14790 0 _0422_
rlabel metal2 38686 13430 38686 13430 0 _0423_
rlabel metal1 36708 13974 36708 13974 0 _0424_
rlabel metal1 43838 20944 43838 20944 0 _0425_
rlabel metal1 44206 18802 44206 18802 0 _0426_
rlabel metal2 46138 19686 46138 19686 0 _0427_
rlabel metal1 27876 18938 27876 18938 0 _0428_
rlabel metal2 28750 19890 28750 19890 0 _0429_
rlabel metal1 28750 23188 28750 23188 0 _0430_
rlabel metal1 29854 20978 29854 20978 0 _0431_
rlabel via1 29770 19686 29770 19686 0 _0432_
rlabel metal1 29578 19346 29578 19346 0 _0433_
rlabel metal1 27876 19686 27876 19686 0 _0434_
rlabel metal1 33120 19686 33120 19686 0 _0435_
rlabel metal1 34454 19924 34454 19924 0 _0436_
rlabel metal1 33956 18598 33956 18598 0 _0437_
rlabel metal2 33718 20213 33718 20213 0 _0438_
rlabel metal1 40434 20434 40434 20434 0 _0439_
rlabel metal1 37598 23018 37598 23018 0 _0440_
rlabel metal1 38740 21590 38740 21590 0 _0441_
rlabel metal2 38318 19720 38318 19720 0 _0442_
rlabel metal1 36846 20978 36846 20978 0 _0443_
rlabel metal1 36892 21488 36892 21488 0 _0444_
rlabel metal1 35834 21590 35834 21590 0 _0445_
rlabel metal1 35604 21998 35604 21998 0 _0446_
rlabel metal1 39698 21046 39698 21046 0 _0447_
rlabel metal1 38962 19822 38962 19822 0 _0448_
rlabel metal1 37536 19822 37536 19822 0 _0449_
rlabel metal2 36294 19482 36294 19482 0 _0450_
rlabel metal1 40848 15946 40848 15946 0 _0451_
rlabel metal1 30958 13396 30958 13396 0 _0452_
rlabel metal1 33488 12818 33488 12818 0 _0453_
rlabel metal2 33258 12517 33258 12517 0 _0454_
rlabel metal2 40802 11866 40802 11866 0 _0455_
rlabel via1 42090 10115 42090 10115 0 _0456_
rlabel metal2 28658 15980 28658 15980 0 _0457_
rlabel via1 40437 12070 40437 12070 0 _0458_
rlabel metal1 39514 13498 39514 13498 0 _0459_
rlabel metal1 26726 16082 26726 16082 0 _0460_
rlabel metal2 26634 16694 26634 16694 0 _0461_
rlabel metal1 38134 12614 38134 12614 0 _0462_
rlabel metal1 38226 11220 38226 11220 0 _0463_
rlabel metal1 37214 12274 37214 12274 0 _0464_
rlabel metal1 45126 10778 45126 10778 0 _0465_
rlabel metal1 38226 10098 38226 10098 0 _0466_
rlabel metal1 36018 9894 36018 9894 0 _0467_
rlabel metal1 35420 6630 35420 6630 0 _0468_
rlabel metal1 39238 3060 39238 3060 0 _0469_
rlabel metal1 44298 10778 44298 10778 0 _0470_
rlabel metal1 40710 9928 40710 9928 0 _0471_
rlabel metal1 36386 10234 36386 10234 0 _0472_
rlabel metal1 33626 7514 33626 7514 0 _0473_
rlabel metal1 32798 3026 32798 3026 0 _0474_
rlabel metal1 25714 14246 25714 14246 0 _0475_
rlabel metal1 28658 11186 28658 11186 0 _0476_
rlabel metal1 29394 11254 29394 11254 0 _0477_
rlabel metal2 27462 12410 27462 12410 0 _0478_
rlabel metal1 30130 11254 30130 11254 0 _0479_
rlabel metal2 37306 6256 37306 6256 0 _0480_
rlabel metal1 36064 6290 36064 6290 0 _0481_
rlabel viali 36848 6290 36848 6290 0 _0482_
rlabel metal1 36662 6256 36662 6256 0 _0483_
rlabel metal1 37076 5678 37076 5678 0 _0484_
rlabel metal1 37352 5610 37352 5610 0 _0485_
rlabel metal2 38870 8432 38870 8432 0 _0486_
rlabel metal1 49588 12614 49588 12614 0 _0487_
rlabel metal2 48898 13345 48898 13345 0 _0488_
rlabel metal1 48438 15334 48438 15334 0 _0489_
rlabel metal1 48346 13464 48346 13464 0 _0490_
rlabel metal2 49818 13736 49818 13736 0 _0491_
rlabel metal1 50140 12682 50140 12682 0 _0492_
rlabel metal1 48760 12886 48760 12886 0 _0493_
rlabel metal1 47472 13702 47472 13702 0 _0494_
rlabel metal1 47334 18938 47334 18938 0 _0495_
rlabel metal1 46966 17306 46966 17306 0 _0496_
rlabel metal1 46736 19482 46736 19482 0 _0497_
rlabel metal1 47978 20298 47978 20298 0 _0498_
rlabel metal1 47242 19890 47242 19890 0 _0499_
rlabel metal1 48760 20298 48760 20298 0 _0500_
rlabel metal1 47012 19822 47012 19822 0 _0501_
rlabel metal1 46276 19890 46276 19890 0 _0502_
rlabel metal1 46182 7854 46182 7854 0 _0503_
rlabel metal1 44666 7242 44666 7242 0 _0504_
rlabel metal1 46414 5678 46414 5678 0 _0505_
rlabel metal2 46414 6868 46414 6868 0 _0506_
rlabel metal2 45862 9554 45862 9554 0 _0507_
rlabel metal1 46368 10234 46368 10234 0 _0508_
rlabel metal1 37582 10608 37582 10608 0 _0509_
rlabel metal2 37398 10846 37398 10846 0 _0510_
rlabel metal1 30176 7378 30176 7378 0 _0511_
rlabel metal1 30866 5202 30866 5202 0 _0512_
rlabel metal1 30774 5338 30774 5338 0 _0513_
rlabel metal1 30406 6324 30406 6324 0 _0514_
rlabel metal1 29946 6358 29946 6358 0 _0515_
rlabel metal2 30406 6562 30406 6562 0 _0516_
rlabel metal1 31947 8330 31947 8330 0 _0517_
rlabel metal1 29762 10574 29762 10574 0 _0518_
rlabel metal1 38732 7854 38732 7854 0 _0519_
rlabel metal1 42964 8466 42964 8466 0 _0520_
rlabel metal2 48438 17034 48438 17034 0 _0521_
rlabel metal1 42826 19482 42826 19482 0 _0522_
rlabel metal1 31970 12648 31970 12648 0 _0523_
rlabel metal1 32660 13498 32660 13498 0 _0524_
rlabel metal1 39974 16558 39974 16558 0 _0525_
rlabel metal1 28612 16218 28612 16218 0 _0526_
rlabel metal2 29118 15300 29118 15300 0 _0527_
rlabel metal1 28474 16762 28474 16762 0 _0528_
rlabel metal1 40250 10676 40250 10676 0 _0529_
rlabel metal1 41814 12818 41814 12818 0 _0530_
rlabel metal1 32798 19890 32798 19890 0 _0531_
rlabel metal1 34500 18938 34500 18938 0 _0532_
rlabel metal1 38870 11322 38870 11322 0 _0533_
rlabel metal2 37858 12619 37858 12619 0 _0534_
rlabel metal2 37490 22372 37490 22372 0 _0535_
rlabel metal1 40204 20298 40204 20298 0 _0536_
rlabel metal1 38456 20434 38456 20434 0 _0537_
rlabel metal1 36018 17612 36018 17612 0 _0538_
rlabel viali 36941 18190 36941 18190 0 _0539_
rlabel metal2 38870 17714 38870 17714 0 _0540_
rlabel metal1 38824 17170 38824 17170 0 _0541_
rlabel metal1 34914 23290 34914 23290 0 _0542_
rlabel metal2 35650 23426 35650 23426 0 _0543_
rlabel metal1 34914 23120 34914 23120 0 _0544_
rlabel metal1 35190 23732 35190 23732 0 _0545_
rlabel metal1 36110 23732 36110 23732 0 _0546_
rlabel metal1 34914 23664 34914 23664 0 _0547_
rlabel metal1 36892 23290 36892 23290 0 _0548_
rlabel metal1 37766 23120 37766 23120 0 _0549_
rlabel metal1 38916 23018 38916 23018 0 _0550_
rlabel metal1 35742 17136 35742 17136 0 _0551_
rlabel metal1 33948 19482 33948 19482 0 _0552_
rlabel metal2 32890 19040 32890 19040 0 _0553_
rlabel metal1 34099 18394 34099 18394 0 _0554_
rlabel metal1 31832 17306 31832 17306 0 _0555_
rlabel metal1 32614 18122 32614 18122 0 _0556_
rlabel metal1 33672 18122 33672 18122 0 _0557_
rlabel metal1 46874 15878 46874 15878 0 _0558_
rlabel metal1 33534 19890 33534 19890 0 _0559_
rlabel metal2 29118 23426 29118 23426 0 _0560_
rlabel metal1 28796 23290 28796 23290 0 _0561_
rlabel metal1 32338 23732 32338 23732 0 _0562_
rlabel metal1 31418 23528 31418 23528 0 _0563_
rlabel metal1 30590 23732 30590 23732 0 _0564_
rlabel metal1 32522 22406 32522 22406 0 _0565_
rlabel metal1 31510 23630 31510 23630 0 _0566_
rlabel metal1 32660 22474 32660 22474 0 _0567_
rlabel via1 31878 23171 31878 23171 0 _0568_
rlabel metal1 29762 23086 29762 23086 0 _0569_
rlabel metal1 30636 21318 30636 21318 0 _0570_
rlabel metal1 30828 21658 30828 21658 0 _0571_
rlabel metal2 31050 21869 31050 21869 0 _0572_
rlabel metal2 28934 24820 28934 24820 0 _0573_
rlabel metal1 29946 24378 29946 24378 0 _0574_
rlabel metal1 28612 23766 28612 23766 0 _0575_
rlabel metal1 28290 23630 28290 23630 0 _0576_
rlabel metal1 27646 22610 27646 22610 0 _0577_
rlabel metal1 27278 22746 27278 22746 0 _0578_
rlabel metal1 28336 18122 28336 18122 0 _0579_
rlabel metal1 29210 18088 29210 18088 0 _0580_
rlabel metal1 30682 18156 30682 18156 0 _0581_
rlabel metal1 28152 17646 28152 17646 0 _0582_
rlabel metal1 27278 19278 27278 19278 0 _0583_
rlabel metal1 27002 19414 27002 19414 0 _0584_
rlabel metal1 27002 19278 27002 19278 0 _0585_
rlabel metal1 26818 20944 26818 20944 0 _0586_
rlabel metal2 26542 20434 26542 20434 0 _0587_
rlabel metal1 26910 21114 26910 21114 0 _0588_
rlabel metal1 30314 2448 30314 2448 0 _0589_
rlabel metal1 43378 18734 43378 18734 0 _0590_
rlabel metal2 32660 14348 32660 14348 0 _0591_
rlabel metal1 32154 12886 32154 12886 0 _0592_
rlabel metal1 31188 12750 31188 12750 0 _0593_
rlabel metal1 40618 2482 40618 2482 0 _0594_
rlabel metal1 26772 15674 26772 15674 0 _0595_
rlabel metal1 30038 14416 30038 14416 0 _0596_
rlabel metal1 34638 17000 34638 17000 0 _0597_
rlabel metal1 30731 11866 30731 11866 0 _0598_
rlabel metal2 40066 8364 40066 8364 0 _0599_
rlabel metal1 36386 10574 36386 10574 0 _0600_
rlabel metal1 36570 8908 36570 8908 0 _0601_
rlabel metal1 26864 15470 26864 15470 0 _0602_
rlabel metal2 26358 15351 26358 15351 0 _0603_
rlabel metal2 51474 8976 51474 8976 0 _0604_
rlabel metal1 41906 7854 41906 7854 0 _0605_
rlabel metal2 42550 10506 42550 10506 0 _0606_
rlabel metal1 35742 8466 35742 8466 0 _0607_
rlabel metal1 36202 6970 36202 6970 0 _0608_
rlabel viali 44486 14994 44486 14994 0 _0609_
rlabel metal1 41574 7922 41574 7922 0 _0610_
rlabel metal3 37559 13804 37559 13804 0 clk
rlabel metal1 34316 20434 34316 20434 0 clknet_0_clk
rlabel metal1 27462 3094 27462 3094 0 clknet_4_0_0_clk
rlabel metal1 45356 4658 45356 4658 0 clknet_4_10_0_clk
rlabel metal2 52026 12240 52026 12240 0 clknet_4_11_0_clk
rlabel metal1 40158 16048 40158 16048 0 clknet_4_12_0_clk
rlabel metal1 37490 19958 37490 19958 0 clknet_4_13_0_clk
rlabel metal2 52302 15470 52302 15470 0 clknet_4_14_0_clk
rlabel metal2 47610 19006 47610 19006 0 clknet_4_15_0_clk
rlabel metal1 22540 12750 22540 12750 0 clknet_4_1_0_clk
rlabel metal1 35098 2890 35098 2890 0 clknet_4_2_0_clk
rlabel metal1 36110 13294 36110 13294 0 clknet_4_3_0_clk
rlabel metal1 25208 14926 25208 14926 0 clknet_4_4_0_clk
rlabel metal1 30130 21998 30130 21998 0 clknet_4_5_0_clk
rlabel metal2 37306 14960 37306 14960 0 clknet_4_6_0_clk
rlabel metal1 33994 24820 33994 24820 0 clknet_4_7_0_clk
rlabel metal1 37858 7378 37858 7378 0 clknet_4_8_0_clk
rlabel metal1 39698 13294 39698 13294 0 clknet_4_9_0_clk
rlabel metal1 30958 12206 30958 12206 0 conv1.addr\[8\]
rlabel metal1 33948 8466 33948 8466 0 conv1.data_valid
rlabel metal1 33764 15130 33764 15130 0 conv1.done
rlabel metal2 33442 7616 33442 7616 0 conv1.psram_ce_n
rlabel metal1 32430 2958 32430 2958 0 conv1.psram_ctrl.counter\[0\]
rlabel metal1 33488 5134 33488 5134 0 conv1.psram_ctrl.counter\[1\]
rlabel metal1 30636 3434 30636 3434 0 conv1.psram_ctrl.counter\[2\]
rlabel metal2 29578 6630 29578 6630 0 conv1.psram_ctrl.counter\[3\]
rlabel metal1 29624 5202 29624 5202 0 conv1.psram_ctrl.counter\[4\]
rlabel via1 29946 5763 29946 5763 0 conv1.psram_ctrl.counter\[5\]
rlabel metal1 27646 6800 27646 6800 0 conv1.psram_ctrl.counter\[6\]
rlabel metal1 30130 6290 30130 6290 0 conv1.psram_ctrl.counter\[7\]
rlabel metal1 30590 12682 30590 12682 0 conv1.psram_ctrl.has_wait_states
rlabel metal1 30728 7786 30728 7786 0 conv1.psram_ctrl.nstate
rlabel metal1 28796 6358 28796 6358 0 conv1.psram_ctrl.sck
rlabel metal1 31694 9044 31694 9044 0 conv1.psram_ctrl.start
rlabel metal1 32476 8058 32476 8058 0 conv1.psram_ctrl.state
rlabel metal2 33994 14892 33994 14892 0 conv1.state\[0\]
rlabel metal2 32246 12478 32246 12478 0 conv1.state\[1\]
rlabel metal1 32062 12172 32062 12172 0 conv1.state\[2\]
rlabel metal1 32660 12818 32660 12818 0 conv1.state\[3\]
rlabel metal1 32752 14042 32752 14042 0 conv1.state\[5\]
rlabel metal1 26358 15130 26358 15130 0 conv2.addr\[8\]
rlabel metal2 25162 14586 25162 14586 0 conv2.addr\[9\]
rlabel metal1 31050 15130 31050 15130 0 conv2.data_out_valid
rlabel metal1 35006 15028 35006 15028 0 conv2.data_valid
rlabel metal1 33350 10676 33350 10676 0 conv2.psram_ce_n
rlabel metal1 26956 12818 26956 12818 0 conv2.psram_ctrl.counter\[0\]
rlabel metal1 25898 12954 25898 12954 0 conv2.psram_ctrl.counter\[1\]
rlabel metal1 27416 12070 27416 12070 0 conv2.psram_ctrl.counter\[2\]
rlabel metal1 28290 11118 28290 11118 0 conv2.psram_ctrl.counter\[3\]
rlabel metal2 25806 10591 25806 10591 0 conv2.psram_ctrl.counter\[4\]
rlabel metal1 27968 10574 27968 10574 0 conv2.psram_ctrl.counter\[5\]
rlabel metal2 27002 9010 27002 9010 0 conv2.psram_ctrl.counter\[6\]
rlabel metal1 27922 8568 27922 8568 0 conv2.psram_ctrl.counter\[7\]
rlabel metal1 29256 14246 29256 14246 0 conv2.psram_ctrl.has_wait_states
rlabel metal1 29440 9622 29440 9622 0 conv2.psram_ctrl.nstate
rlabel metal1 33534 10608 33534 10608 0 conv2.psram_ctrl.sck
rlabel metal1 29118 12614 29118 12614 0 conv2.psram_ctrl.start
rlabel metal2 29302 10370 29302 10370 0 conv2.psram_ctrl.state
rlabel metal1 31050 16082 31050 16082 0 conv2.state\[0\]
rlabel metal1 28842 15878 28842 15878 0 conv2.state\[1\]
rlabel metal1 28290 15402 28290 15402 0 conv2.state\[2\]
rlabel metal1 29486 16116 29486 16116 0 conv2.state\[3\]
rlabel metal1 28658 16626 28658 16626 0 conv2.state\[5\]
rlabel via2 68402 60571 68402 60571 0 done
rlabel metal2 36294 6766 36294 6766 0 fc1.addr\[10\]
rlabel metal2 35834 7310 35834 7310 0 fc1.addr\[8\]
rlabel metal1 39008 13294 39008 13294 0 fc1.data_out_valid
rlabel metal1 38778 9588 38778 9588 0 fc1.psram_ce_n
rlabel metal1 37444 6766 37444 6766 0 fc1.psram_ctrl.counter\[0\]
rlabel metal1 38272 3434 38272 3434 0 fc1.psram_ctrl.counter\[1\]
rlabel metal2 36846 4284 36846 4284 0 fc1.psram_ctrl.counter\[2\]
rlabel metal1 38042 6222 38042 6222 0 fc1.psram_ctrl.counter\[3\]
rlabel metal1 36754 6256 36754 6256 0 fc1.psram_ctrl.counter\[4\]
rlabel metal1 39330 2924 39330 2924 0 fc1.psram_ctrl.counter\[5\]
rlabel metal2 41170 5372 41170 5372 0 fc1.psram_ctrl.counter\[6\]
rlabel metal1 41354 5576 41354 5576 0 fc1.psram_ctrl.counter\[7\]
rlabel metal1 36386 8874 36386 8874 0 fc1.psram_ctrl.has_wait_states
rlabel metal1 38502 7480 38502 7480 0 fc1.psram_ctrl.nstate
rlabel metal2 38962 9724 38962 9724 0 fc1.psram_ctrl.sck
rlabel metal1 38686 7956 38686 7956 0 fc1.psram_ctrl.start
rlabel metal2 39974 6970 39974 6970 0 fc1.psram_ctrl.state
rlabel metal2 36754 14620 36754 14620 0 fc1.state\[0\]
rlabel metal1 36892 12206 36892 12206 0 fc1.state\[1\]
rlabel metal1 37306 11322 37306 11322 0 fc1.state\[2\]
rlabel metal1 36570 12886 36570 12886 0 fc1.state\[3\]
rlabel metal1 38272 11866 38272 11866 0 fc1.state\[5\]
rlabel metal1 43700 7514 43700 7514 0 fc2.addr\[10\]
rlabel metal1 42274 7480 42274 7480 0 fc2.addr\[8\]
rlabel metal1 43102 12954 43102 12954 0 fc2.done
rlabel metal1 45080 11730 45080 11730 0 fc2.psram_ce_n
rlabel metal1 46092 6290 46092 6290 0 fc2.psram_ctrl.counter\[0\]
rlabel metal1 48898 6154 48898 6154 0 fc2.psram_ctrl.counter\[1\]
rlabel metal1 48530 5168 48530 5168 0 fc2.psram_ctrl.counter\[2\]
rlabel metal1 45908 6766 45908 6766 0 fc2.psram_ctrl.counter\[3\]
rlabel metal1 48346 7276 48346 7276 0 fc2.psram_ctrl.counter\[4\]
rlabel metal1 46092 10030 46092 10030 0 fc2.psram_ctrl.counter\[5\]
rlabel metal1 48254 9486 48254 9486 0 fc2.psram_ctrl.counter\[6\]
rlabel metal1 49220 10030 49220 10030 0 fc2.psram_ctrl.counter\[7\]
rlabel metal1 42366 10200 42366 10200 0 fc2.psram_ctrl.has_wait_states
rlabel metal1 43056 8534 43056 8534 0 fc2.psram_ctrl.nstate
rlabel metal2 45126 9248 45126 9248 0 fc2.psram_ctrl.sck
rlabel metal1 44114 9044 44114 9044 0 fc2.psram_ctrl.start
rlabel metal1 45218 8330 45218 8330 0 fc2.psram_ctrl.state
rlabel metal1 40066 14450 40066 14450 0 fc2.state\[0\]
rlabel metal1 41078 11764 41078 11764 0 fc2.state\[1\]
rlabel metal1 41584 9418 41584 9418 0 fc2.state\[2\]
rlabel metal1 40618 13158 40618 13158 0 fc2.state\[3\]
rlabel metal2 41262 11764 41262 11764 0 fc2.state\[5\]
rlabel metal1 47472 14926 47472 14926 0 maxpool.addr\[11\]
rlabel metal1 48208 15470 48208 15470 0 maxpool.addr\[8\]
rlabel metal1 42274 15572 42274 15572 0 maxpool.done
rlabel metal2 44850 13668 44850 13668 0 maxpool.psram_ce_n
rlabel metal1 49404 12818 49404 12818 0 maxpool.psram_ctrl.counter\[0\]
rlabel metal1 49174 13226 49174 13226 0 maxpool.psram_ctrl.counter\[1\]
rlabel metal1 52256 11730 52256 11730 0 maxpool.psram_ctrl.counter\[2\]
rlabel metal1 51060 12138 51060 12138 0 maxpool.psram_ctrl.counter\[3\]
rlabel metal1 52854 12852 52854 12852 0 maxpool.psram_ctrl.counter\[4\]
rlabel metal1 51290 13804 51290 13804 0 maxpool.psram_ctrl.counter\[5\]
rlabel metal1 51888 16218 51888 16218 0 maxpool.psram_ctrl.counter\[6\]
rlabel metal1 53958 15470 53958 15470 0 maxpool.psram_ctrl.counter\[7\]
rlabel metal1 48392 16762 48392 16762 0 maxpool.psram_ctrl.nstate
rlabel metal1 48760 13838 48760 13838 0 maxpool.psram_ctrl.sck
rlabel metal1 48530 16660 48530 16660 0 maxpool.psram_ctrl.start
rlabel metal1 49036 16626 49036 16626 0 maxpool.psram_ctrl.state
rlabel metal1 45862 13804 45862 13804 0 maxpool.start
rlabel metal2 43838 15470 43838 15470 0 maxpool.state\[0\]
rlabel metal1 41584 16626 41584 16626 0 maxpool.state\[2\]
rlabel metal1 40020 15878 40020 15878 0 maxpool.state\[3\]
rlabel metal2 40894 16592 40894 16592 0 maxpool.state\[4\]
rlabel metal2 36110 20604 36110 20604 0 mfcc.dct.data_valid
rlabel metal1 37214 16660 37214 16660 0 mfcc.dct.dct_valid
rlabel metal1 36110 23188 36110 23188 0 mfcc.dct.input_counter\[0\]
rlabel metal1 35742 23596 35742 23596 0 mfcc.dct.input_counter\[1\]
rlabel metal1 35374 24310 35374 24310 0 mfcc.dct.input_counter\[2\]
rlabel metal1 38226 23528 38226 23528 0 mfcc.dct.input_counter\[3\]
rlabel metal2 38594 23324 38594 23324 0 mfcc.dct.input_counter\[4\]
rlabel metal1 38594 21624 38594 21624 0 mfcc.dct.output_counter\[0\]
rlabel metal1 39698 20468 39698 20468 0 mfcc.dct.output_counter\[1\]
rlabel metal1 38870 20298 38870 20298 0 mfcc.dct.output_counter\[2\]
rlabel metal1 37582 18088 37582 18088 0 mfcc.dct.output_counter\[3\]
rlabel metal1 37628 18258 37628 18258 0 mfcc.dct.output_counter\[4\]
rlabel metal1 38686 18326 38686 18326 0 mfcc.dct.output_counter\[5\]
rlabel metal2 36662 20995 36662 20995 0 mfcc.dct.state\[0\]
rlabel metal1 37030 21386 37030 21386 0 mfcc.dct.state\[1\]
rlabel metal1 32338 19856 32338 19856 0 mfcc.log.data_valid
rlabel metal1 33580 19210 33580 19210 0 mfcc.log.shift_count\[0\]
rlabel metal2 32154 18020 32154 18020 0 mfcc.log.shift_count\[1\]
rlabel metal1 33534 17646 33534 17646 0 mfcc.log.shift_count\[2\]
rlabel metal2 34730 17918 34730 17918 0 mfcc.log.shift_count\[3\]
rlabel metal1 32660 20774 32660 20774 0 mfcc.log.state\[0\]
rlabel metal1 33994 19346 33994 19346 0 mfcc.log.state\[1\]
rlabel metal1 33764 21454 33764 21454 0 mfcc.log.state\[2\]
rlabel metal1 29532 18258 29532 18258 0 mfcc.mel.coeff_counter\[0\]
rlabel metal1 27370 18938 27370 18938 0 mfcc.mel.coeff_counter\[1\]
rlabel metal1 27232 18598 27232 18598 0 mfcc.mel.coeff_counter\[2\]
rlabel metal1 27094 20332 27094 20332 0 mfcc.mel.coeff_counter\[3\]
rlabel metal1 27462 21318 27462 21318 0 mfcc.mel.coeff_counter\[4\]
rlabel via1 31970 23613 31970 23613 0 mfcc.mel.filter_counter\[0\]
rlabel metal1 32499 24378 32499 24378 0 mfcc.mel.filter_counter\[1\]
rlabel metal1 32476 22610 32476 22610 0 mfcc.mel.filter_counter\[2\]
rlabel metal1 31418 22542 31418 22542 0 mfcc.mel.filter_counter\[3\]
rlabel metal2 29210 23426 29210 23426 0 mfcc.mel.filter_counter\[4\]
rlabel via1 28934 23087 28934 23087 0 mfcc.mel.filter_counter\[5\]
rlabel metal1 28934 22141 28934 22141 0 mfcc.mel.state\[0\]
rlabel metal1 29578 19788 29578 19788 0 mfcc.mel.state\[1\]
rlabel metal1 38870 15878 38870 15878 0 mfcc.mfcc_valid
rlabel metal2 1794 19584 1794 19584 0 net1
rlabel metal2 58650 1588 58650 1588 0 net10
rlabel metal1 38042 8500 38042 8500 0 net100
rlabel metal1 41354 12138 41354 12138 0 net101
rlabel metal2 39238 11322 39238 11322 0 net102
rlabel metal1 41998 13328 41998 13328 0 net103
rlabel metal1 39831 13974 39831 13974 0 net104
rlabel viali 48346 14383 48346 14383 0 net105
rlabel metal1 29072 16490 29072 16490 0 net106
rlabel metal1 29854 15436 29854 15436 0 net107
rlabel metal1 44252 19346 44252 19346 0 net108
rlabel metal1 36800 14382 36800 14382 0 net109
rlabel metal2 28014 68255 28014 68255 0 net11
rlabel metal2 36294 13090 36294 13090 0 net110
rlabel metal1 34592 14586 34592 14586 0 net111
rlabel metal2 34086 13090 34086 13090 0 net112
rlabel metal1 30130 21012 30130 21012 0 net113
rlabel metal1 38732 22950 38732 22950 0 net114
rlabel metal2 33442 21216 33442 21216 0 net115
rlabel metal1 33626 20570 33626 20570 0 net116
rlabel metal1 31832 14994 31832 14994 0 net117
rlabel metal2 31694 15266 31694 15266 0 net118
rlabel metal1 43608 20910 43608 20910 0 net119
rlabel via2 68494 63325 68494 63325 0 net12
rlabel metal2 39238 14212 39238 14212 0 net120
rlabel metal1 34086 16082 34086 16082 0 net121
rlabel metal2 42918 16082 42918 16082 0 net122
rlabel metal1 43097 16082 43097 16082 0 net123
rlabel metal1 39008 17850 39008 17850 0 net124
rlabel metal1 34960 17714 34960 17714 0 net125
rlabel metal1 43194 7888 43194 7888 0 net126
rlabel metal1 36708 6766 36708 6766 0 net127
rlabel metal1 35599 7446 35599 7446 0 net128
rlabel metal2 26266 14858 26266 14858 0 net129
rlabel metal2 68310 1027 68310 1027 0 net13
rlabel metal1 40802 12818 40802 12818 0 net130
rlabel metal2 41078 13090 41078 13090 0 net131
rlabel metal1 26864 14246 26864 14246 0 net132
rlabel metal1 27048 14994 27048 14994 0 net133
rlabel metal1 45448 19482 45448 19482 0 net134
rlabel metal1 39330 17238 39330 17238 0 net135
rlabel metal1 48714 9554 48714 9554 0 net136
rlabel metal1 32568 22746 32568 22746 0 net137
rlabel metal1 42320 7786 42320 7786 0 net138
rlabel metal1 41078 7922 41078 7922 0 net139
rlabel metal2 33166 67371 33166 67371 0 net14
rlabel metal2 27646 21692 27646 21692 0 net140
rlabel metal1 44666 18394 44666 18394 0 net141
rlabel metal1 45678 18326 45678 18326 0 net142
rlabel metal1 45903 17578 45903 17578 0 net143
rlabel metal1 29670 10710 29670 10710 0 net144
rlabel metal1 35604 23154 35604 23154 0 net145
rlabel metal1 35880 8806 35880 8806 0 net146
rlabel metal1 34776 7854 34776 7854 0 net147
rlabel metal1 47242 14416 47242 14416 0 net148
rlabel metal1 46782 14586 46782 14586 0 net149
rlabel metal2 25162 1588 25162 1588 0 net15
rlabel metal1 37996 21658 37996 21658 0 net150
rlabel metal1 38548 22610 38548 22610 0 net151
rlabel metal1 27140 8534 27140 8534 0 net152
rlabel metal2 32430 17850 32430 17850 0 net153
rlabel metal1 42136 5270 42136 5270 0 net154
rlabel metal1 37260 23086 37260 23086 0 net155
rlabel metal1 37720 23222 37720 23222 0 net156
rlabel metal1 39146 20570 39146 20570 0 net157
rlabel metal1 37122 19856 37122 19856 0 net158
rlabel metal2 32062 20264 32062 20264 0 net159
rlabel via2 68494 17051 68494 17051 0 net16
rlabel metal1 26358 19856 26358 19856 0 net160
rlabel metal1 25525 20502 25525 20502 0 net161
rlabel metal1 33120 17578 33120 17578 0 net162
rlabel metal1 32885 17170 32885 17170 0 net163
rlabel metal1 38778 7786 38778 7786 0 net164
rlabel metal1 31418 11866 31418 11866 0 net165
rlabel metal1 29210 12172 29210 12172 0 net166
rlabel metal1 45586 15674 45586 15674 0 net167
rlabel metal1 44344 14926 44344 14926 0 net168
rlabel metal1 33396 18666 33396 18666 0 net169
rlabel via2 68494 22491 68494 22491 0 net17
rlabel metal1 44206 8874 44206 8874 0 net170
rlabel via1 36184 18734 36184 18734 0 net171
rlabel metal2 36662 19618 36662 19618 0 net172
rlabel metal1 28152 15130 28152 15130 0 net173
rlabel metal1 28469 14314 28469 14314 0 net174
rlabel metal1 46874 21556 46874 21556 0 net175
rlabel metal1 43930 21624 43930 21624 0 net176
rlabel metal1 52256 15538 52256 15538 0 net177
rlabel metal2 50462 15844 50462 15844 0 net178
rlabel metal2 32062 12937 32062 12937 0 net179
rlabel via2 68494 57885 68494 57885 0 net18
rlabel metal1 29941 12886 29941 12886 0 net180
rlabel metal1 50462 9894 50462 9894 0 net181
rlabel metal1 46276 17034 46276 17034 0 net182
rlabel metal1 46858 16490 46858 16490 0 net183
rlabel metal1 48990 16762 48990 16762 0 net184
rlabel metal2 48254 22202 48254 22202 0 net185
rlabel metal1 36570 17646 36570 17646 0 net186
rlabel metal1 41630 11118 41630 11118 0 net187
rlabel metal2 43102 10914 43102 10914 0 net188
rlabel metal1 31648 13362 31648 13362 0 net189
rlabel metal2 58926 68255 58926 68255 0 net19
rlabel metal2 32798 12104 32798 12104 0 net190
rlabel metal1 32660 8602 32660 8602 0 net191
rlabel metal2 31786 23868 31786 23868 0 net192
rlabel metal1 37490 10030 37490 10030 0 net193
rlabel metal2 36754 9826 36754 9826 0 net194
rlabel metal1 40066 20570 40066 20570 0 net195
rlabel metal1 35374 10676 35374 10676 0 net196
rlabel metal2 36662 9452 36662 9452 0 net197
rlabel metal1 49220 7446 49220 7446 0 net198
rlabel metal1 43332 18598 43332 18598 0 net199
rlabel metal2 68402 27421 68402 27421 0 net2
rlabel via2 68494 14365 68494 14365 0 net20
rlabel metal1 47104 22066 47104 22066 0 net200
rlabel metal1 46000 23018 46000 23018 0 net201
rlabel metal2 44942 16320 44942 16320 0 net202
rlabel metal1 46858 15402 46858 15402 0 net203
rlabel metal1 29532 24106 29532 24106 0 net204
rlabel metal1 35466 23698 35466 23698 0 net205
rlabel metal2 33626 20060 33626 20060 0 net206
rlabel metal1 34904 20910 34904 20910 0 net207
rlabel metal1 40250 14960 40250 14960 0 net208
rlabel metal1 30912 23630 30912 23630 0 net209
rlabel via2 68494 66011 68494 66011 0 net21
rlabel metal2 41906 11084 41906 11084 0 net210
rlabel metal2 41906 8908 41906 8908 0 net211
rlabel metal1 52026 15062 52026 15062 0 net212
rlabel metal1 50738 21420 50738 21420 0 net213
rlabel metal1 36800 10642 36800 10642 0 net214
rlabel metal1 36013 11050 36013 11050 0 net215
rlabel metal1 40986 9996 40986 9996 0 net216
rlabel metal1 32844 12274 32844 12274 0 net217
rlabel metal1 32287 11050 32287 11050 0 net218
rlabel metal1 39560 3366 39560 3366 0 net219
rlabel metal3 820 12988 820 12988 0 net22
rlabel metal2 51382 13124 51382 13124 0 net220
rlabel metal1 27876 17646 27876 17646 0 net221
rlabel metal2 51888 12580 51888 12580 0 net222
rlabel metal1 48530 12954 48530 12954 0 net223
rlabel metal1 36478 4488 36478 4488 0 net224
rlabel metal1 39882 4624 39882 4624 0 net225
rlabel metal1 46782 5100 46782 5100 0 net226
rlabel metal1 28612 6766 28612 6766 0 net227
rlabel metal1 37030 4114 37030 4114 0 net228
rlabel metal1 30544 4046 30544 4046 0 net229
rlabel metal3 820 29308 820 29308 0 net23
rlabel metal1 32944 20570 32944 20570 0 net230
rlabel metal1 33534 5338 33534 5338 0 net231
rlabel metal1 32331 4794 32331 4794 0 net232
rlabel metal1 25714 12274 25714 12274 0 net233
rlabel metal1 50600 11730 50600 11730 0 net234
rlabel metal1 46046 6834 46046 6834 0 net235
rlabel metal1 27876 5270 27876 5270 0 net236
rlabel metal1 27554 15640 27554 15640 0 net237
rlabel metal1 27876 13906 27876 13906 0 net238
rlabel metal1 25162 9146 25162 9146 0 net239
rlabel via2 68494 11611 68494 11611 0 net24
rlabel metal1 36110 24242 36110 24242 0 net240
rlabel metal1 24702 9894 24702 9894 0 net241
rlabel metal1 39330 3944 39330 3944 0 net242
rlabel metal2 25070 10778 25070 10778 0 net243
rlabel metal1 30866 11254 30866 11254 0 net244
rlabel metal2 41630 19482 41630 19482 0 net245
rlabel metal1 47748 6358 47748 6358 0 net246
rlabel metal1 47104 17850 47104 17850 0 net247
rlabel metal1 41722 11730 41722 11730 0 net248
rlabel metal1 35972 11730 35972 11730 0 net249
rlabel metal3 820 37468 820 37468 0 net25
rlabel metal2 28750 15164 28750 15164 0 net250
rlabel metal3 820 48348 820 48348 0 net26
rlabel metal2 38318 68255 38318 68255 0 net27
rlabel metal2 64078 68255 64078 68255 0 net28
rlabel metal2 7130 1588 7130 1588 0 net29
rlabel metal1 68034 60690 68034 60690 0 net3
rlabel via2 68494 52445 68494 52445 0 net30
rlabel metal3 820 45628 820 45628 0 net31
rlabel metal3 820 7548 820 7548 0 net32
rlabel via2 68494 3485 68494 3485 0 net33
rlabel metal2 53498 1588 53498 1588 0 net34
rlabel via2 68494 30685 68494 30685 0 net35
rlabel via2 68494 25245 68494 25245 0 net36
rlabel metal2 25438 68255 25438 68255 0 net37
rlabel via2 68494 55131 68494 55131 0 net38
rlabel metal3 820 10268 820 10268 0 net39
rlabel metal1 22126 2346 22126 2346 0 net4
rlabel metal2 17434 1588 17434 1588 0 net40
rlabel via2 68494 8925 68494 8925 0 net41
rlabel metal1 68356 2482 68356 2482 0 net42
rlabel via2 68494 36125 68494 36125 0 net43
rlabel metal3 820 51068 820 51068 0 net44
rlabel via2 68494 44251 68494 44251 0 net45
rlabel via2 68494 19805 68494 19805 0 net46
rlabel metal2 35466 823 35466 823 0 net47
rlabel metal2 61502 68255 61502 68255 0 net48
rlabel metal2 46046 68255 46046 68255 0 net49
rlabel metal1 48438 2414 48438 2414 0 net5
rlabel metal2 30314 1588 30314 1588 0 net50
rlabel metal1 68724 67218 68724 67218 0 net51
rlabel via2 68494 6171 68494 6171 0 net52
rlabel metal2 2254 68255 2254 68255 0 net53
rlabel metal3 820 26588 820 26588 0 net54
rlabel metal3 820 34748 820 34748 0 net55
rlabel metal2 40894 68255 40894 68255 0 net56
rlabel metal2 32890 1588 32890 1588 0 net57
rlabel metal2 17710 68255 17710 68255 0 net58
rlabel metal3 751 64668 751 64668 0 net59
rlabel metal1 29486 7412 29486 7412 0 net6
rlabel metal2 45770 1588 45770 1588 0 net60
rlabel metal2 4554 1588 4554 1588 0 net61
rlabel metal3 820 32028 820 32028 0 net62
rlabel metal2 66378 1588 66378 1588 0 net63
rlabel metal3 820 2108 820 2108 0 net64
rlabel metal2 50922 1588 50922 1588 0 net65
rlabel metal3 1142 56508 1142 56508 0 net66
rlabel metal3 820 42908 820 42908 0 net67
rlabel metal3 820 15708 820 15708 0 net68
rlabel via2 68494 27931 68494 27931 0 net69
rlabel metal3 1142 59228 1142 59228 0 net7
rlabel via2 68494 47005 68494 47005 0 net70
rlabel metal2 56074 1588 56074 1588 0 net71
rlabel via2 68494 49725 68494 49725 0 net72
rlabel metal2 7406 68255 7406 68255 0 net73
rlabel metal2 9982 68255 9982 68255 0 net74
rlabel metal2 46 1656 46 1656 0 net75
rlabel metal2 43194 1588 43194 1588 0 net76
rlabel metal1 12512 67218 12512 67218 0 net77
rlabel metal1 30498 67218 30498 67218 0 net78
rlabel metal3 820 18428 820 18428 0 net79
rlabel metal2 20286 68255 20286 68255 0 net8
rlabel metal1 1288 67218 1288 67218 0 net80
rlabel metal2 9706 1588 9706 1588 0 net81
rlabel metal2 1978 1588 1978 1588 0 net82
rlabel metal3 820 23868 820 23868 0 net83
rlabel via2 68494 41565 68494 41565 0 net84
rlabel metal2 38042 823 38042 823 0 net85
rlabel metal2 53774 68255 53774 68255 0 net86
rlabel metal2 4830 68255 4830 68255 0 net87
rlabel metal2 15134 68255 15134 68255 0 net88
rlabel metal2 56166 68323 56166 68323 0 net89
rlabel metal2 22862 68255 22862 68255 0 net9
rlabel metal2 37858 17000 37858 17000 0 net90
rlabel metal1 43470 9486 43470 9486 0 net91
rlabel metal2 37352 12716 37352 12716 0 net92
rlabel metal1 35098 11764 35098 11764 0 net93
rlabel metal1 31050 9622 31050 9622 0 net94
rlabel metal1 32292 13226 32292 13226 0 net95
rlabel metal1 29670 13260 29670 13260 0 net96
rlabel metal1 41055 16150 41055 16150 0 net97
rlabel metal1 39422 17612 39422 17612 0 net98
rlabel metal1 32292 7378 32292 7378 0 net99
rlabel metal2 12282 1571 12282 1571 0 psram_ce_n
rlabel metal1 26864 2822 26864 2822 0 psram_d[0]
rlabel metal2 48346 1520 48346 1520 0 psram_sck
rlabel metal3 820 21148 820 21148 0 rst
rlabel metal2 46414 19312 46414 19312 0 softmax.addr\[11\]
rlabel metal1 45908 17850 45908 17850 0 softmax.addr\[8\]
rlabel metal1 44620 18122 44620 18122 0 softmax.data_valid
rlabel metal1 44896 14994 44896 14994 0 softmax.psram_ce_n
rlabel metal1 51750 18360 51750 18360 0 softmax.psram_ctrl.counter\[0\]
rlabel metal2 47794 18836 47794 18836 0 softmax.psram_ctrl.counter\[1\]
rlabel metal1 47702 19924 47702 19924 0 softmax.psram_ctrl.counter\[2\]
rlabel metal2 47978 20060 47978 20060 0 softmax.psram_ctrl.counter\[3\]
rlabel metal1 48208 20434 48208 20434 0 softmax.psram_ctrl.counter\[4\]
rlabel metal1 46322 20808 46322 20808 0 softmax.psram_ctrl.counter\[5\]
rlabel metal1 45402 21522 45402 21522 0 softmax.psram_ctrl.counter\[6\]
rlabel metal1 46782 20944 46782 20944 0 softmax.psram_ctrl.counter\[7\]
rlabel metal1 42642 20026 42642 20026 0 softmax.psram_ctrl.nstate
rlabel metal1 45448 14994 45448 14994 0 softmax.psram_ctrl.sck
rlabel metal1 43562 19346 43562 19346 0 softmax.psram_ctrl.start
rlabel metal1 44344 20366 44344 20366 0 softmax.psram_ctrl.state
rlabel metal1 44620 18258 44620 18258 0 softmax.start
rlabel metal1 68540 33490 68540 33490 0 start
rlabel metal1 42550 20774 42550 20774 0 state\[0\]
rlabel metal1 39238 14042 39238 14042 0 state\[1\]
rlabel metal1 40802 19686 40802 19686 0 state\[4\]
rlabel metal1 42550 14280 42550 14280 0 state\[5\]
<< properties >>
string FIXED_BBOX 0 0 70000 70000
<< end >>
