magic
tech sky130A
magscale 1 2
timestamp 1715939645
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 14 2128 68986 67504
<< metal2 >>
rect 18 69200 74 70000
rect 1950 69200 2006 70000
rect 4526 69200 4582 70000
rect 7102 69200 7158 70000
rect 9678 69200 9734 70000
rect 12254 69200 12310 70000
rect 14830 69200 14886 70000
rect 17406 69200 17462 70000
rect 19982 69200 20038 70000
rect 22558 69200 22614 70000
rect 25134 69200 25190 70000
rect 27710 69200 27766 70000
rect 30286 69200 30342 70000
rect 32862 69200 32918 70000
rect 35438 69200 35494 70000
rect 38014 69200 38070 70000
rect 40590 69200 40646 70000
rect 43166 69200 43222 70000
rect 45742 69200 45798 70000
rect 48318 69200 48374 70000
rect 50894 69200 50950 70000
rect 53470 69200 53526 70000
rect 56046 69200 56102 70000
rect 58622 69200 58678 70000
rect 61198 69200 61254 70000
rect 63774 69200 63830 70000
rect 66350 69200 66406 70000
rect 68926 69200 68982 70000
rect 18 0 74 800
rect 1950 0 2006 800
rect 4526 0 4582 800
rect 7102 0 7158 800
rect 9678 0 9734 800
rect 12254 0 12310 800
rect 14830 0 14886 800
rect 17406 0 17462 800
rect 19982 0 20038 800
rect 22558 0 22614 800
rect 25134 0 25190 800
rect 27710 0 27766 800
rect 30286 0 30342 800
rect 32862 0 32918 800
rect 35438 0 35494 800
rect 38014 0 38070 800
rect 40590 0 40646 800
rect 43166 0 43222 800
rect 45742 0 45798 800
rect 48318 0 48374 800
rect 50894 0 50950 800
rect 53470 0 53526 800
rect 56046 0 56102 800
rect 58622 0 58678 800
rect 61198 0 61254 800
rect 63774 0 63830 800
rect 66350 0 66406 800
rect 68282 0 68338 800
<< obsm2 >>
rect 130 69144 1894 69306
rect 2062 69144 4470 69306
rect 4638 69144 7046 69306
rect 7214 69144 9622 69306
rect 9790 69144 12198 69306
rect 12366 69144 14774 69306
rect 14942 69144 17350 69306
rect 17518 69144 19926 69306
rect 20094 69144 22502 69306
rect 22670 69144 25078 69306
rect 25246 69144 27654 69306
rect 27822 69144 30230 69306
rect 30398 69144 32806 69306
rect 32974 69144 35382 69306
rect 35550 69144 37958 69306
rect 38126 69144 40534 69306
rect 40702 69144 43110 69306
rect 43278 69144 45686 69306
rect 45854 69144 48262 69306
rect 48430 69144 50838 69306
rect 51006 69144 53414 69306
rect 53582 69144 55990 69306
rect 56158 69144 58566 69306
rect 58734 69144 61142 69306
rect 61310 69144 63718 69306
rect 63886 69144 66294 69306
rect 66462 69144 68870 69306
rect 20 856 68980 69144
rect 130 711 1894 856
rect 2062 711 4470 856
rect 4638 711 7046 856
rect 7214 711 9622 856
rect 9790 711 12198 856
rect 12366 711 14774 856
rect 14942 711 17350 856
rect 17518 711 19926 856
rect 20094 711 22502 856
rect 22670 711 25078 856
rect 25246 711 27654 856
rect 27822 711 30230 856
rect 30398 711 32806 856
rect 32974 711 35382 856
rect 35550 711 37958 856
rect 38126 711 40534 856
rect 40702 711 43110 856
rect 43278 711 45686 856
rect 45854 711 48262 856
rect 48430 711 50838 856
rect 51006 711 53414 856
rect 53582 711 55990 856
rect 56158 711 58566 856
rect 58734 711 61142 856
rect 61310 711 63718 856
rect 63886 711 66294 856
rect 66462 711 68226 856
rect 68394 711 68980 856
<< metal3 >>
rect 69200 68688 70000 68808
rect 0 67328 800 67448
rect 69200 65968 70000 66088
rect 0 64608 800 64728
rect 69200 63248 70000 63368
rect 0 61888 800 62008
rect 69200 60528 70000 60648
rect 0 59168 800 59288
rect 69200 57808 70000 57928
rect 0 56448 800 56568
rect 69200 55088 70000 55208
rect 0 53728 800 53848
rect 69200 52368 70000 52488
rect 0 51008 800 51128
rect 69200 49648 70000 49768
rect 0 48288 800 48408
rect 69200 46928 70000 47048
rect 0 45568 800 45688
rect 69200 44208 70000 44328
rect 0 42848 800 42968
rect 69200 41488 70000 41608
rect 0 40128 800 40248
rect 69200 38768 70000 38888
rect 0 37408 800 37528
rect 69200 36048 70000 36168
rect 0 34688 800 34808
rect 69200 33328 70000 33448
rect 0 31968 800 32088
rect 69200 30608 70000 30728
rect 0 29248 800 29368
rect 69200 27888 70000 28008
rect 0 26528 800 26648
rect 69200 25168 70000 25288
rect 0 23808 800 23928
rect 69200 22448 70000 22568
rect 0 21088 800 21208
rect 69200 19728 70000 19848
rect 0 18368 800 18488
rect 69200 17008 70000 17128
rect 0 15648 800 15768
rect 69200 14288 70000 14408
rect 0 12928 800 13048
rect 69200 11568 70000 11688
rect 0 10208 800 10328
rect 69200 8848 70000 8968
rect 0 7488 800 7608
rect 69200 6128 70000 6248
rect 0 4768 800 4888
rect 69200 3408 70000 3528
rect 0 2048 800 2168
rect 69200 688 70000 808
<< obsm3 >>
rect 880 67248 69200 67489
rect 798 66168 69200 67248
rect 798 65888 69120 66168
rect 798 64808 69200 65888
rect 880 64528 69200 64808
rect 798 63448 69200 64528
rect 798 63168 69120 63448
rect 798 62088 69200 63168
rect 880 61808 69200 62088
rect 798 60728 69200 61808
rect 798 60448 69120 60728
rect 798 59368 69200 60448
rect 880 59088 69200 59368
rect 798 58008 69200 59088
rect 798 57728 69120 58008
rect 798 56648 69200 57728
rect 880 56368 69200 56648
rect 798 55288 69200 56368
rect 798 55008 69120 55288
rect 798 53928 69200 55008
rect 880 53648 69200 53928
rect 798 52568 69200 53648
rect 798 52288 69120 52568
rect 798 51208 69200 52288
rect 880 50928 69200 51208
rect 798 49848 69200 50928
rect 798 49568 69120 49848
rect 798 48488 69200 49568
rect 880 48208 69200 48488
rect 798 47128 69200 48208
rect 798 46848 69120 47128
rect 798 45768 69200 46848
rect 880 45488 69200 45768
rect 798 44408 69200 45488
rect 798 44128 69120 44408
rect 798 43048 69200 44128
rect 880 42768 69200 43048
rect 798 41688 69200 42768
rect 798 41408 69120 41688
rect 798 40328 69200 41408
rect 880 40048 69200 40328
rect 798 38968 69200 40048
rect 798 38688 69120 38968
rect 798 37608 69200 38688
rect 880 37328 69200 37608
rect 798 36248 69200 37328
rect 798 35968 69120 36248
rect 798 34888 69200 35968
rect 880 34608 69200 34888
rect 798 33528 69200 34608
rect 798 33248 69120 33528
rect 798 32168 69200 33248
rect 880 31888 69200 32168
rect 798 30808 69200 31888
rect 798 30528 69120 30808
rect 798 29448 69200 30528
rect 880 29168 69200 29448
rect 798 28088 69200 29168
rect 798 27808 69120 28088
rect 798 26728 69200 27808
rect 880 26448 69200 26728
rect 798 25368 69200 26448
rect 798 25088 69120 25368
rect 798 24008 69200 25088
rect 880 23728 69200 24008
rect 798 22648 69200 23728
rect 798 22368 69120 22648
rect 798 21288 69200 22368
rect 880 21008 69200 21288
rect 798 19928 69200 21008
rect 798 19648 69120 19928
rect 798 18568 69200 19648
rect 880 18288 69200 18568
rect 798 17208 69200 18288
rect 798 16928 69120 17208
rect 798 15848 69200 16928
rect 880 15568 69200 15848
rect 798 14488 69200 15568
rect 798 14208 69120 14488
rect 798 13128 69200 14208
rect 880 12848 69200 13128
rect 798 11768 69200 12848
rect 798 11488 69120 11768
rect 798 10408 69200 11488
rect 880 10128 69200 10408
rect 798 9048 69200 10128
rect 798 8768 69120 9048
rect 798 7688 69200 8768
rect 880 7408 69200 7688
rect 798 6328 69200 7408
rect 798 6048 69120 6328
rect 798 4968 69200 6048
rect 880 4688 69200 4968
rect 798 3608 69200 4688
rect 798 3328 69120 3608
rect 798 2248 69200 3328
rect 880 1968 69200 2248
rect 798 888 69200 1968
rect 798 715 69120 888
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 37595 3299 37661 13837
<< labels >>
rlabel metal2 s 18 69200 74 70000 6 audio_sample[0]
port 1 nsew signal input
rlabel metal3 s 69200 68688 70000 68808 6 audio_sample[10]
port 2 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 audio_sample[11]
port 3 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 audio_sample[12]
port 4 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 audio_sample[13]
port 5 nsew signal input
rlabel metal2 s 43166 69200 43222 70000 6 audio_sample[14]
port 6 nsew signal input
rlabel metal2 s 66350 69200 66406 70000 6 audio_sample[15]
port 7 nsew signal input
rlabel metal2 s 50894 69200 50950 70000 6 audio_sample[1]
port 8 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 audio_sample[2]
port 9 nsew signal input
rlabel metal2 s 35438 69200 35494 70000 6 audio_sample[3]
port 10 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 audio_sample[4]
port 11 nsew signal input
rlabel metal3 s 69200 38768 70000 38888 6 audio_sample[5]
port 12 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 audio_sample[6]
port 13 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 audio_sample[7]
port 14 nsew signal input
rlabel metal2 s 48318 69200 48374 70000 6 audio_sample[8]
port 15 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 audio_sample[9]
port 16 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 clk
port 17 nsew signal input
rlabel metal3 s 69200 60528 70000 60648 6 done
port 18 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 io_oeb[0]
port 19 nsew signal output
rlabel metal3 s 69200 22448 70000 22568 6 io_oeb[10]
port 20 nsew signal output
rlabel metal3 s 69200 57808 70000 57928 6 io_oeb[11]
port 21 nsew signal output
rlabel metal2 s 58622 69200 58678 70000 6 io_oeb[12]
port 22 nsew signal output
rlabel metal3 s 69200 14288 70000 14408 6 io_oeb[13]
port 23 nsew signal output
rlabel metal3 s 69200 65968 70000 66088 6 io_oeb[14]
port 24 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 io_oeb[15]
port 25 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 io_oeb[16]
port 26 nsew signal output
rlabel metal3 s 69200 11568 70000 11688 6 io_oeb[17]
port 27 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 io_oeb[18]
port 28 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_oeb[19]
port 29 nsew signal output
rlabel metal2 s 19982 69200 20038 70000 6 io_oeb[1]
port 30 nsew signal output
rlabel metal2 s 38014 69200 38070 70000 6 io_oeb[20]
port 31 nsew signal output
rlabel metal2 s 63774 69200 63830 70000 6 io_oeb[21]
port 32 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 io_oeb[22]
port 33 nsew signal output
rlabel metal3 s 69200 52368 70000 52488 6 io_oeb[23]
port 34 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 io_oeb[24]
port 35 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 io_oeb[25]
port 36 nsew signal output
rlabel metal3 s 69200 3408 70000 3528 6 io_oeb[26]
port 37 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 io_oeb[27]
port 38 nsew signal output
rlabel metal3 s 69200 30608 70000 30728 6 io_oeb[28]
port 39 nsew signal output
rlabel metal3 s 69200 25168 70000 25288 6 io_oeb[29]
port 40 nsew signal output
rlabel metal2 s 22558 69200 22614 70000 6 io_oeb[2]
port 41 nsew signal output
rlabel metal2 s 25134 69200 25190 70000 6 io_oeb[30]
port 42 nsew signal output
rlabel metal3 s 69200 55088 70000 55208 6 io_oeb[31]
port 43 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 io_oeb[32]
port 44 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 io_oeb[33]
port 45 nsew signal output
rlabel metal3 s 69200 8848 70000 8968 6 io_oeb[34]
port 46 nsew signal output
rlabel metal3 s 69200 688 70000 808 6 io_oeb[35]
port 47 nsew signal output
rlabel metal3 s 69200 36048 70000 36168 6 io_oeb[36]
port 48 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 io_oeb[37]
port 49 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 io_oeb[3]
port 50 nsew signal output
rlabel metal2 s 27710 69200 27766 70000 6 io_oeb[4]
port 51 nsew signal output
rlabel metal3 s 69200 63248 70000 63368 6 io_oeb[5]
port 52 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 io_oeb[6]
port 53 nsew signal output
rlabel metal2 s 32862 69200 32918 70000 6 io_oeb[7]
port 54 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 io_oeb[8]
port 55 nsew signal output
rlabel metal3 s 69200 17008 70000 17128 6 io_oeb[9]
port 56 nsew signal output
rlabel metal3 s 69200 44208 70000 44328 6 io_out[0]
port 57 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 io_out[10]
port 58 nsew signal output
rlabel metal2 s 40590 69200 40646 70000 6 io_out[11]
port 59 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 io_out[12]
port 60 nsew signal output
rlabel metal2 s 17406 69200 17462 70000 6 io_out[13]
port 61 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 io_out[14]
port 62 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 io_out[15]
port 63 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 io_out[16]
port 64 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_out[17]
port 65 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 io_out[18]
port 66 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 io_out[19]
port 67 nsew signal output
rlabel metal3 s 69200 19728 70000 19848 6 io_out[1]
port 68 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 io_out[20]
port 69 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 io_out[21]
port 70 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 io_out[22]
port 71 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 io_out[23]
port 72 nsew signal output
rlabel metal3 s 69200 27888 70000 28008 6 io_out[24]
port 73 nsew signal output
rlabel metal3 s 69200 46928 70000 47048 6 io_out[25]
port 74 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 io_out[26]
port 75 nsew signal output
rlabel metal3 s 69200 49648 70000 49768 6 io_out[27]
port 76 nsew signal output
rlabel metal2 s 7102 69200 7158 70000 6 io_out[28]
port 77 nsew signal output
rlabel metal2 s 9678 69200 9734 70000 6 io_out[29]
port 78 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 io_out[2]
port 79 nsew signal output
rlabel metal2 s 18 0 74 800 6 io_out[30]
port 80 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 io_out[31]
port 81 nsew signal output
rlabel metal2 s 12254 69200 12310 70000 6 io_out[32]
port 82 nsew signal output
rlabel metal2 s 30286 69200 30342 70000 6 io_out[33]
port 83 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_out[34]
port 84 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 io_out[35]
port 85 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 io_out[36]
port 86 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 io_out[37]
port 87 nsew signal output
rlabel metal2 s 61198 69200 61254 70000 6 io_out[3]
port 88 nsew signal output
rlabel metal2 s 45742 69200 45798 70000 6 io_out[4]
port 89 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 io_out[5]
port 90 nsew signal output
rlabel metal2 s 68926 69200 68982 70000 6 io_out[6]
port 91 nsew signal output
rlabel metal3 s 69200 6128 70000 6248 6 io_out[7]
port 92 nsew signal output
rlabel metal2 s 1950 69200 2006 70000 6 io_out[8]
port 93 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 io_out[9]
port 94 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 psram_ce_n
port 95 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 psram_d[0]
port 96 nsew signal bidirectional
rlabel metal3 s 0 23808 800 23928 6 psram_d[1]
port 97 nsew signal bidirectional
rlabel metal3 s 69200 41488 70000 41608 6 psram_d[2]
port 98 nsew signal bidirectional
rlabel metal2 s 38014 0 38070 800 6 psram_d[3]
port 99 nsew signal bidirectional
rlabel metal2 s 56046 69200 56102 70000 6 psram_douten[0]
port 100 nsew signal output
rlabel metal2 s 53470 69200 53526 70000 6 psram_douten[1]
port 101 nsew signal output
rlabel metal2 s 4526 69200 4582 70000 6 psram_douten[2]
port 102 nsew signal output
rlabel metal2 s 14830 69200 14886 70000 6 psram_douten[3]
port 103 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 psram_sck
port 104 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 rst
port 105 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 sample_valid
port 106 nsew signal input
rlabel metal3 s 69200 33328 70000 33448 6 start
port 107 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 108 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 108 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 108 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 109 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 109 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3495338
string GDS_FILE /home/iamme/asic_tools/caravel_user_project/openlane/cnn_kws_accel/runs/24_05_17_12_34/results/signoff/cnn_kws_accel.magic.gds
string GDS_START 470050
<< end >>

