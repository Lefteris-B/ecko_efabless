magic
tech sky130A
magscale 1 2
timestamp 1715980346
<< viali >>
rect 13001 67201 13035 67235
rect 30389 67201 30423 67235
rect 39405 67201 39439 67235
rect 1409 64957 1443 64991
rect 68477 56117 68511 56151
rect 1777 46529 1811 46563
rect 1501 46325 1535 46359
rect 1777 37281 1811 37315
rect 1501 37145 1535 37179
rect 21005 29121 21039 29155
rect 22661 29121 22695 29155
rect 24041 29121 24075 29155
rect 24777 29121 24811 29155
rect 23949 29053 23983 29087
rect 22753 28985 22787 29019
rect 24133 28985 24167 29019
rect 21097 28917 21131 28951
rect 23305 28917 23339 28951
rect 24869 28917 24903 28951
rect 24409 28577 24443 28611
rect 20085 28509 20119 28543
rect 22201 28509 22235 28543
rect 20361 28441 20395 28475
rect 22109 28441 22143 28475
rect 22477 28441 22511 28475
rect 24685 28441 24719 28475
rect 26433 28441 26467 28475
rect 23949 28373 23983 28407
rect 20453 28169 20487 28203
rect 20729 28169 20763 28203
rect 22201 28169 22235 28203
rect 21097 28101 21131 28135
rect 22687 28101 22721 28135
rect 20637 28033 20671 28067
rect 21189 28033 21223 28067
rect 22385 28033 22419 28067
rect 22477 28033 22511 28067
rect 22569 28033 22603 28067
rect 22845 28033 22879 28067
rect 25697 28033 25731 28067
rect 68385 28033 68419 28067
rect 21373 27965 21407 27999
rect 23213 27965 23247 27999
rect 25421 27965 25455 27999
rect 23949 27897 23983 27931
rect 23765 27829 23799 27863
rect 68293 27829 68327 27863
rect 22937 27625 22971 27659
rect 25053 27625 25087 27659
rect 23121 27489 23155 27523
rect 23305 27489 23339 27523
rect 24409 27489 24443 27523
rect 25237 27489 25271 27523
rect 26157 27489 26191 27523
rect 20821 27421 20855 27455
rect 21005 27421 21039 27455
rect 23213 27421 23247 27455
rect 23397 27421 23431 27455
rect 24547 27421 24581 27455
rect 24869 27421 24903 27455
rect 25145 27421 25179 27455
rect 25329 27421 25363 27455
rect 25421 27421 25455 27455
rect 27997 27421 28031 27455
rect 30113 27421 30147 27455
rect 30481 27421 30515 27455
rect 24685 27353 24719 27387
rect 24777 27353 24811 27387
rect 26424 27353 26458 27387
rect 28264 27353 28298 27387
rect 20913 27285 20947 27319
rect 25513 27285 25547 27319
rect 27537 27285 27571 27319
rect 29377 27285 29411 27319
rect 29561 27285 29595 27319
rect 30297 27285 30331 27319
rect 19625 27081 19659 27115
rect 21439 27081 21473 27115
rect 22661 27081 22695 27115
rect 23029 27081 23063 27115
rect 23121 27081 23155 27115
rect 24685 27081 24719 27115
rect 24777 27081 24811 27115
rect 26709 27081 26743 27115
rect 28641 27081 28675 27115
rect 21649 27013 21683 27047
rect 23213 27013 23247 27047
rect 24199 27013 24233 27047
rect 24409 27013 24443 27047
rect 25237 27013 25271 27047
rect 25421 27013 25455 27047
rect 27077 27013 27111 27047
rect 27905 27013 27939 27047
rect 30196 27013 30230 27047
rect 17877 26945 17911 26979
rect 20085 26945 20119 26979
rect 22293 26945 22327 26979
rect 22477 26945 22511 26979
rect 22753 26945 22787 26979
rect 23489 26945 23523 26979
rect 24317 26945 24351 26979
rect 24501 26945 24535 26979
rect 24961 26945 24995 26979
rect 25145 26945 25179 26979
rect 25605 26945 25639 26979
rect 25697 26945 25731 26979
rect 25881 26945 25915 26979
rect 26617 26945 26651 26979
rect 26801 26945 26835 26979
rect 27353 26945 27387 26979
rect 27629 26945 27663 26979
rect 27721 26945 27755 26979
rect 28457 26945 28491 26979
rect 28825 26945 28859 26979
rect 29101 26945 29135 26979
rect 29285 26945 29319 26979
rect 32853 26945 32887 26979
rect 18153 26877 18187 26911
rect 20177 26877 20211 26911
rect 20361 26877 20395 26911
rect 21097 26877 21131 26911
rect 23581 26877 23615 26911
rect 24041 26877 24075 26911
rect 25789 26877 25823 26911
rect 27077 26877 27111 26911
rect 27261 26877 27295 26911
rect 29929 26877 29963 26911
rect 32597 26877 32631 26911
rect 34621 26877 34655 26911
rect 21281 26809 21315 26843
rect 23397 26809 23431 26843
rect 33977 26809 34011 26843
rect 19717 26741 19751 26775
rect 20545 26741 20579 26775
rect 21465 26741 21499 26775
rect 22293 26741 22327 26775
rect 22845 26741 22879 26775
rect 23489 26741 23523 26775
rect 23857 26741 23891 26775
rect 27445 26741 27479 26775
rect 31309 26741 31343 26775
rect 34069 26741 34103 26775
rect 18153 26537 18187 26571
rect 18797 26537 18831 26571
rect 19809 26537 19843 26571
rect 21373 26537 21407 26571
rect 22753 26537 22787 26571
rect 23121 26537 23155 26571
rect 25329 26537 25363 26571
rect 27445 26537 27479 26571
rect 28549 26537 28583 26571
rect 29561 26537 29595 26571
rect 33517 26537 33551 26571
rect 19533 26469 19567 26503
rect 21833 26469 21867 26503
rect 28181 26469 28215 26503
rect 31861 26469 31895 26503
rect 25421 26401 25455 26435
rect 31309 26401 31343 26435
rect 32413 26401 32447 26435
rect 32597 26401 32631 26435
rect 32965 26401 32999 26435
rect 33057 26401 33091 26435
rect 12173 26333 12207 26367
rect 14289 26333 14323 26367
rect 18245 26333 18279 26367
rect 18705 26333 18739 26367
rect 19441 26333 19475 26367
rect 19717 26333 19751 26367
rect 19993 26333 20027 26367
rect 20177 26333 20211 26367
rect 20269 26333 20303 26367
rect 20637 26333 20671 26367
rect 20821 26333 20855 26367
rect 21097 26333 21131 26367
rect 21557 26333 21591 26367
rect 21741 26333 21775 26367
rect 21833 26333 21867 26367
rect 22017 26333 22051 26367
rect 22845 26333 22879 26367
rect 22937 26333 22971 26367
rect 25145 26333 25179 26367
rect 27721 26333 27755 26367
rect 29745 26333 29779 26367
rect 29837 26333 29871 26367
rect 30021 26333 30055 26367
rect 30113 26333 30147 26367
rect 30573 26333 30607 26367
rect 30665 26333 30699 26367
rect 31033 26333 31067 26367
rect 31493 26333 31527 26367
rect 31769 26333 31803 26367
rect 31861 26333 31895 26367
rect 31953 26333 31987 26367
rect 32321 26333 32355 26367
rect 32505 26333 32539 26367
rect 32781 26333 32815 26367
rect 32873 26333 32907 26367
rect 33241 26333 33275 26367
rect 33517 26333 33551 26367
rect 12449 26265 12483 26299
rect 14197 26265 14231 26299
rect 19349 26265 19383 26299
rect 21005 26265 21039 26299
rect 22661 26265 22695 26299
rect 27997 26265 28031 26299
rect 28549 26265 28583 26299
rect 30757 26265 30791 26299
rect 30895 26265 30929 26299
rect 32137 26265 32171 26299
rect 33333 26265 33367 26299
rect 13921 26197 13955 26231
rect 24961 26197 24995 26231
rect 27629 26197 27663 26231
rect 27813 26197 27847 26231
rect 28733 26197 28767 26231
rect 30389 26197 30423 26231
rect 31677 26197 31711 26231
rect 12357 25993 12391 26027
rect 19901 25993 19935 26027
rect 21189 25993 21223 26027
rect 21925 25993 21959 26027
rect 22661 25993 22695 26027
rect 28273 25993 28307 26027
rect 18429 25925 18463 25959
rect 20821 25925 20855 25959
rect 28089 25925 28123 25959
rect 11989 25857 12023 25891
rect 12725 25857 12759 25891
rect 14013 25857 14047 25891
rect 18153 25857 18187 25891
rect 20637 25857 20671 25891
rect 21373 25857 21407 25891
rect 21557 25857 21591 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22569 25857 22603 25891
rect 22753 25857 22787 25891
rect 23305 25857 23339 25891
rect 24777 25857 24811 25891
rect 24961 25857 24995 25891
rect 25145 25857 25179 25891
rect 25697 25857 25731 25891
rect 26801 25857 26835 25891
rect 27169 25857 27203 25891
rect 27353 25857 27387 25891
rect 27629 25857 27663 25891
rect 27721 25857 27755 25891
rect 29193 25857 29227 25891
rect 30113 25857 30147 25891
rect 31217 25857 31251 25891
rect 31309 25857 31343 25891
rect 12817 25789 12851 25823
rect 13001 25789 13035 25823
rect 14289 25789 14323 25823
rect 25053 25789 25087 25823
rect 25421 25789 25455 25823
rect 29929 25789 29963 25823
rect 30297 25789 30331 25823
rect 31125 25789 31159 25823
rect 12173 25721 12207 25755
rect 25237 25721 25271 25755
rect 25605 25721 25639 25755
rect 26985 25721 27019 25755
rect 15761 25653 15795 25687
rect 21005 25653 21039 25687
rect 23121 25653 23155 25687
rect 24593 25653 24627 25687
rect 25329 25653 25363 25687
rect 26709 25653 26743 25687
rect 27537 25653 27571 25687
rect 28089 25653 28123 25687
rect 29377 25653 29411 25687
rect 30941 25653 30975 25687
rect 13645 25449 13679 25483
rect 14381 25449 14415 25483
rect 16313 25449 16347 25483
rect 23581 25449 23615 25483
rect 25145 25449 25179 25483
rect 27537 25449 27571 25483
rect 29285 25449 29319 25483
rect 31861 25449 31895 25483
rect 32137 25449 32171 25483
rect 13461 25381 13495 25415
rect 14657 25381 14691 25415
rect 27445 25381 27479 25415
rect 32505 25381 32539 25415
rect 10149 25313 10183 25347
rect 11897 25313 11931 25347
rect 12725 25313 12759 25347
rect 15301 25313 15335 25347
rect 19257 25313 19291 25347
rect 22109 25313 22143 25347
rect 24409 25313 24443 25347
rect 26065 25313 26099 25347
rect 27721 25313 27755 25347
rect 27997 25313 28031 25347
rect 31125 25313 31159 25347
rect 13277 25245 13311 25279
rect 13369 25245 13403 25279
rect 13553 25245 13587 25279
rect 13645 25245 13679 25279
rect 13829 25245 13863 25279
rect 14565 25245 14599 25279
rect 16037 25245 16071 25279
rect 16405 25245 16439 25279
rect 16681 25245 16715 25279
rect 18705 25245 18739 25279
rect 22017 25245 22051 25279
rect 22201 25245 22235 25279
rect 22477 25245 22511 25279
rect 22845 25245 22879 25279
rect 23029 25245 23063 25279
rect 23305 25245 23339 25279
rect 23397 25245 23431 25279
rect 23857 25245 23891 25279
rect 24961 25245 24995 25279
rect 25324 25245 25358 25279
rect 25641 25245 25675 25279
rect 25789 25245 25823 25279
rect 26332 25245 26366 25279
rect 27813 25245 27847 25279
rect 27905 25245 27939 25279
rect 28641 25245 28675 25279
rect 28825 25245 28859 25279
rect 28917 25245 28951 25279
rect 29101 25245 29135 25279
rect 30941 25245 30975 25279
rect 31217 25245 31251 25279
rect 31309 25245 31343 25279
rect 31677 25245 31711 25279
rect 33885 25245 33919 25279
rect 36093 25245 36127 25279
rect 36277 25245 36311 25279
rect 10425 25177 10459 25211
rect 13093 25177 13127 25211
rect 15025 25177 15059 25211
rect 15485 25177 15519 25211
rect 16926 25177 16960 25211
rect 18153 25177 18187 25211
rect 19533 25177 19567 25211
rect 22569 25177 22603 25211
rect 22661 25177 22695 25211
rect 23213 25177 23247 25211
rect 23673 25177 23707 25211
rect 25421 25177 25455 25211
rect 25513 25177 25547 25211
rect 30674 25177 30708 25211
rect 31493 25177 31527 25211
rect 31585 25177 31619 25211
rect 31953 25177 31987 25211
rect 33618 25177 33652 25211
rect 12173 25109 12207 25143
rect 12909 25109 12943 25143
rect 15117 25109 15151 25143
rect 18061 25109 18095 25143
rect 21005 25109 21039 25143
rect 22293 25109 22327 25143
rect 24041 25109 24075 25143
rect 28733 25109 28767 25143
rect 29561 25109 29595 25143
rect 32153 25109 32187 25143
rect 32321 25109 32355 25143
rect 36185 25109 36219 25143
rect 11161 24905 11195 24939
rect 11989 24905 12023 24939
rect 12357 24905 12391 24939
rect 15393 24905 15427 24939
rect 16497 24905 16531 24939
rect 19441 24905 19475 24939
rect 19625 24905 19659 24939
rect 22477 24905 22511 24939
rect 25421 24905 25455 24939
rect 25697 24905 25731 24939
rect 29535 24905 29569 24939
rect 30941 24905 30975 24939
rect 32229 24905 32263 24939
rect 33057 24905 33091 24939
rect 11529 24837 11563 24871
rect 11745 24837 11779 24871
rect 22293 24837 22327 24871
rect 23213 24837 23247 24871
rect 23949 24837 23983 24871
rect 29745 24837 29779 24871
rect 31953 24837 31987 24871
rect 35992 24837 36026 24871
rect 23443 24803 23477 24837
rect 11069 24769 11103 24803
rect 12173 24769 12207 24803
rect 12449 24769 12483 24803
rect 13093 24769 13127 24803
rect 14013 24769 14047 24803
rect 14280 24769 14314 24803
rect 16313 24769 16347 24803
rect 16681 24769 16715 24803
rect 16937 24769 16971 24803
rect 18705 24769 18739 24803
rect 19257 24769 19291 24803
rect 19533 24769 19567 24803
rect 21465 24769 21499 24803
rect 22017 24769 22051 24803
rect 22201 24769 22235 24803
rect 22385 24769 22419 24803
rect 25605 24769 25639 24803
rect 25789 24769 25823 24803
rect 28273 24769 28307 24803
rect 28457 24769 28491 24803
rect 30849 24769 30883 24803
rect 31033 24769 31067 24803
rect 31493 24769 31527 24803
rect 31677 24769 31711 24803
rect 32413 24769 32447 24803
rect 32505 24769 32539 24803
rect 32597 24769 32631 24803
rect 32873 24769 32907 24803
rect 34253 24769 34287 24803
rect 34520 24769 34554 24803
rect 35725 24769 35759 24803
rect 8309 24701 8343 24735
rect 8585 24701 8619 24735
rect 10057 24701 10091 24735
rect 10425 24701 10459 24735
rect 13277 24701 13311 24735
rect 20545 24701 20579 24735
rect 23029 24701 23063 24735
rect 23673 24701 23707 24735
rect 28549 24701 28583 24735
rect 32781 24701 32815 24735
rect 37289 24701 37323 24735
rect 11897 24633 11931 24667
rect 23581 24633 23615 24667
rect 29377 24633 29411 24667
rect 31309 24633 31343 24667
rect 37105 24633 37139 24667
rect 10977 24565 11011 24599
rect 11713 24565 11747 24599
rect 12909 24565 12943 24599
rect 18061 24565 18095 24599
rect 18153 24565 18187 24599
rect 19901 24565 19935 24599
rect 20913 24565 20947 24599
rect 21925 24565 21959 24599
rect 23397 24565 23431 24599
rect 28089 24565 28123 24599
rect 29561 24565 29595 24599
rect 31861 24565 31895 24599
rect 35633 24565 35667 24599
rect 37933 24565 37967 24599
rect 9413 24361 9447 24395
rect 10701 24361 10735 24395
rect 12633 24361 12667 24395
rect 13185 24361 13219 24395
rect 14473 24361 14507 24395
rect 16497 24361 16531 24395
rect 19625 24361 19659 24395
rect 22385 24361 22419 24395
rect 24685 24361 24719 24395
rect 30573 24361 30607 24395
rect 30757 24361 30791 24395
rect 32413 24361 32447 24395
rect 34989 24361 35023 24395
rect 37289 24361 37323 24395
rect 16865 24293 16899 24327
rect 15485 24225 15519 24259
rect 16957 24225 16991 24259
rect 17509 24225 17543 24259
rect 19073 24225 19107 24259
rect 20269 24225 20303 24259
rect 20729 24225 20763 24259
rect 27445 24225 27479 24259
rect 31953 24225 31987 24259
rect 32137 24225 32171 24259
rect 32689 24225 32723 24259
rect 37197 24225 37231 24259
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 10885 24157 10919 24191
rect 10977 24157 11011 24191
rect 11253 24157 11287 24191
rect 11345 24157 11379 24191
rect 11529 24157 11563 24191
rect 12173 24157 12207 24191
rect 12449 24157 12483 24191
rect 13093 24157 13127 24191
rect 13277 24157 13311 24191
rect 14473 24157 14507 24191
rect 14657 24157 14691 24191
rect 15393 24157 15427 24191
rect 16037 24157 16071 24191
rect 16313 24157 16347 24191
rect 16497 24157 16531 24191
rect 16589 24157 16623 24191
rect 16865 24157 16899 24191
rect 20453 24157 20487 24191
rect 22661 24157 22695 24191
rect 22753 24157 22787 24191
rect 24593 24157 24627 24191
rect 25421 24157 25455 24191
rect 27353 24157 27387 24191
rect 28273 24157 28307 24191
rect 28365 24157 28399 24191
rect 30297 24157 30331 24191
rect 32045 24157 32079 24191
rect 32229 24157 32263 24191
rect 32873 24157 32907 24191
rect 32965 24157 32999 24191
rect 34437 24157 34471 24191
rect 35173 24157 35207 24191
rect 35449 24157 35483 24191
rect 35633 24157 35667 24191
rect 35725 24157 35759 24191
rect 36369 24157 36403 24191
rect 37013 24157 37047 24191
rect 37381 24157 37415 24191
rect 37473 24157 37507 24191
rect 11069 24089 11103 24123
rect 11437 24089 11471 24123
rect 12725 24089 12759 24123
rect 12909 24089 12943 24123
rect 18806 24089 18840 24123
rect 19993 24089 20027 24123
rect 22293 24089 22327 24123
rect 28089 24089 28123 24123
rect 34170 24089 34204 24123
rect 10609 24021 10643 24055
rect 12265 24021 12299 24055
rect 14749 24021 14783 24055
rect 16681 24021 16715 24055
rect 17693 24021 17727 24055
rect 20085 24021 20119 24055
rect 22201 24021 22235 24055
rect 22937 24021 22971 24055
rect 25329 24021 25363 24055
rect 26985 24021 27019 24055
rect 27905 24021 27939 24055
rect 28549 24021 28583 24055
rect 32689 24021 32723 24055
rect 33057 24021 33091 24055
rect 36461 24021 36495 24055
rect 9689 23817 9723 23851
rect 10149 23817 10183 23851
rect 10517 23817 10551 23851
rect 10701 23817 10735 23851
rect 11897 23817 11931 23851
rect 12909 23817 12943 23851
rect 16957 23817 16991 23851
rect 18521 23817 18555 23851
rect 21005 23817 21039 23851
rect 24593 23817 24627 23851
rect 25421 23817 25455 23851
rect 25697 23817 25731 23851
rect 27721 23817 27755 23851
rect 35817 23817 35851 23851
rect 11253 23749 11287 23783
rect 11529 23749 11563 23783
rect 11729 23749 11763 23783
rect 28834 23749 28868 23783
rect 33149 23749 33183 23783
rect 33885 23749 33919 23783
rect 10057 23681 10091 23715
rect 10333 23681 10367 23715
rect 10609 23681 10643 23715
rect 10885 23681 10919 23715
rect 11161 23681 11195 23715
rect 11345 23681 11379 23715
rect 12725 23681 12759 23715
rect 14657 23681 14691 23715
rect 14749 23681 14783 23715
rect 16497 23681 16531 23715
rect 17141 23681 17175 23715
rect 17601 23681 17635 23715
rect 17785 23681 17819 23715
rect 18061 23681 18095 23715
rect 18245 23681 18279 23715
rect 18337 23681 18371 23715
rect 19625 23681 19659 23715
rect 19892 23681 19926 23715
rect 22753 23681 22787 23715
rect 25329 23681 25363 23715
rect 25605 23681 25639 23715
rect 26249 23681 26283 23715
rect 26525 23681 26559 23715
rect 26709 23681 26743 23715
rect 34069 23681 34103 23715
rect 34161 23681 34195 23715
rect 36001 23681 36035 23715
rect 36185 23681 36219 23715
rect 36553 23681 36587 23715
rect 7941 23613 7975 23647
rect 8217 23613 8251 23647
rect 12541 23613 12575 23647
rect 14013 23613 14047 23647
rect 16221 23613 16255 23647
rect 17325 23613 17359 23647
rect 17877 23613 17911 23647
rect 22385 23613 22419 23647
rect 22661 23613 22695 23647
rect 25145 23613 25179 23647
rect 26985 23613 27019 23647
rect 27629 23613 27663 23647
rect 29101 23613 29135 23647
rect 29929 23613 29963 23647
rect 31033 23613 31067 23647
rect 33701 23613 33735 23647
rect 36093 23613 36127 23647
rect 36277 23613 36311 23647
rect 36829 23613 36863 23647
rect 11069 23545 11103 23579
rect 16405 23545 16439 23579
rect 30205 23545 30239 23579
rect 30389 23545 30423 23579
rect 36645 23545 36679 23579
rect 11713 23477 11747 23511
rect 14841 23477 14875 23511
rect 16313 23477 16347 23511
rect 17601 23477 17635 23511
rect 25605 23477 25639 23511
rect 26709 23477 26743 23511
rect 30481 23477 30515 23511
rect 33885 23477 33919 23511
rect 36737 23477 36771 23511
rect 9045 23273 9079 23307
rect 11161 23273 11195 23307
rect 11345 23273 11379 23307
rect 13001 23273 13035 23307
rect 18153 23273 18187 23307
rect 20361 23273 20395 23307
rect 25973 23273 26007 23307
rect 27445 23273 27479 23307
rect 27997 23273 28031 23307
rect 28181 23273 28215 23307
rect 28457 23273 28491 23307
rect 30941 23273 30975 23307
rect 31401 23273 31435 23307
rect 32597 23273 32631 23307
rect 32781 23273 32815 23307
rect 32965 23273 32999 23307
rect 35449 23273 35483 23307
rect 36093 23273 36127 23307
rect 17141 23205 17175 23239
rect 27629 23205 27663 23239
rect 35265 23205 35299 23239
rect 36185 23205 36219 23239
rect 12633 23137 12667 23171
rect 14565 23137 14599 23171
rect 17509 23137 17543 23171
rect 18245 23137 18279 23171
rect 29561 23137 29595 23171
rect 32229 23137 32263 23171
rect 33701 23137 33735 23171
rect 34069 23137 34103 23171
rect 35909 23137 35943 23171
rect 8953 23069 8987 23103
rect 10149 23069 10183 23103
rect 11621 23069 11655 23103
rect 11713 23069 11747 23103
rect 12449 23069 12483 23103
rect 12817 23069 12851 23103
rect 13185 23069 13219 23103
rect 14381 23069 14415 23103
rect 14473 23069 14507 23103
rect 16129 23069 16163 23103
rect 16865 23069 16899 23103
rect 17141 23069 17175 23103
rect 17693 23069 17727 23103
rect 18429 23069 18463 23103
rect 18613 23069 18647 23103
rect 18705 23069 18739 23103
rect 20177 23069 20211 23103
rect 20361 23069 20395 23103
rect 23213 23069 23247 23103
rect 24133 23069 24167 23103
rect 24593 23069 24627 23103
rect 26065 23069 26099 23103
rect 26332 23069 26366 23103
rect 31217 23069 31251 23103
rect 31493 23069 31527 23103
rect 31677 23069 31711 23103
rect 33517 23069 33551 23103
rect 33885 23069 33919 23103
rect 34161 23069 34195 23103
rect 34345 23069 34379 23103
rect 35725 23069 35759 23103
rect 36093 23069 36127 23103
rect 36553 23069 36587 23103
rect 37013 23069 37047 23103
rect 37280 23069 37314 23103
rect 11329 23001 11363 23035
rect 11529 23001 11563 23035
rect 14197 23001 14231 23035
rect 14832 23001 14866 23035
rect 23581 23001 23615 23035
rect 24860 23001 24894 23035
rect 27997 23001 28031 23035
rect 28273 23001 28307 23035
rect 29806 23001 29840 23035
rect 32413 23001 32447 23035
rect 34253 23001 34287 23035
rect 35633 23001 35667 23035
rect 35817 23001 35851 23035
rect 36369 23001 36403 23035
rect 36461 23001 36495 23035
rect 36737 23001 36771 23035
rect 10701 22933 10735 22967
rect 12541 22933 12575 22967
rect 12725 22933 12759 22967
rect 14295 22933 14329 22967
rect 15945 22933 15979 22967
rect 16773 22933 16807 22967
rect 16957 22933 16991 22967
rect 17785 22933 17819 22967
rect 18889 22933 18923 22967
rect 23305 22933 23339 22967
rect 28473 22933 28507 22967
rect 28641 22933 28675 22967
rect 31033 22933 31067 22967
rect 32623 22933 32657 22967
rect 35433 22933 35467 22967
rect 38393 22933 38427 22967
rect 11069 22729 11103 22763
rect 13093 22729 13127 22763
rect 13277 22729 13311 22763
rect 21925 22729 21959 22763
rect 24041 22729 24075 22763
rect 24317 22729 24351 22763
rect 28273 22729 28307 22763
rect 29377 22729 29411 22763
rect 31769 22729 31803 22763
rect 37289 22729 37323 22763
rect 10149 22661 10183 22695
rect 10287 22661 10321 22695
rect 10793 22661 10827 22695
rect 12173 22661 12207 22695
rect 14390 22661 14424 22695
rect 15853 22661 15887 22695
rect 18521 22661 18555 22695
rect 23049 22661 23083 22695
rect 26801 22661 26835 22695
rect 27905 22661 27939 22695
rect 33609 22661 33643 22695
rect 36429 22661 36463 22695
rect 36645 22661 36679 22695
rect 7941 22593 7975 22627
rect 9965 22593 9999 22627
rect 10057 22593 10091 22627
rect 10425 22593 10459 22627
rect 10701 22593 10735 22627
rect 10885 22593 10919 22627
rect 11345 22593 11379 22627
rect 11713 22593 11747 22627
rect 11989 22593 12023 22627
rect 12081 22593 12115 22627
rect 12357 22593 12391 22627
rect 12541 22593 12575 22627
rect 12633 22593 12667 22627
rect 12909 22593 12943 22627
rect 14657 22593 14691 22627
rect 15025 22593 15059 22627
rect 15209 22593 15243 22627
rect 15485 22593 15519 22627
rect 15761 22593 15795 22627
rect 16497 22593 16531 22627
rect 17601 22593 17635 22627
rect 17693 22593 17727 22627
rect 17877 22593 17911 22627
rect 18061 22593 18095 22627
rect 19257 22593 19291 22627
rect 19441 22593 19475 22627
rect 20545 22593 20579 22627
rect 20729 22593 20763 22627
rect 21281 22593 21315 22627
rect 23397 22593 23431 22627
rect 23581 22593 23615 22627
rect 23765 22593 23799 22627
rect 23857 22593 23891 22627
rect 25441 22593 25475 22627
rect 25697 22593 25731 22627
rect 27077 22593 27111 22627
rect 29561 22593 29595 22627
rect 29653 22593 29687 22627
rect 29837 22593 29871 22627
rect 29929 22593 29963 22627
rect 30656 22593 30690 22627
rect 32321 22593 32355 22627
rect 32781 22593 32815 22627
rect 33793 22593 33827 22627
rect 34060 22593 34094 22627
rect 37933 22593 37967 22627
rect 8217 22525 8251 22559
rect 9781 22525 9815 22559
rect 11253 22525 11287 22559
rect 11621 22525 11655 22559
rect 11897 22525 11931 22559
rect 12725 22525 12759 22559
rect 15117 22525 15151 22559
rect 17325 22525 17359 22559
rect 17417 22525 17451 22559
rect 19717 22525 19751 22559
rect 23305 22525 23339 22559
rect 26065 22525 26099 22559
rect 28825 22525 28859 22559
rect 30389 22525 30423 22559
rect 32597 22525 32631 22559
rect 35817 22525 35851 22559
rect 9689 22457 9723 22491
rect 10517 22457 10551 22491
rect 11805 22457 11839 22491
rect 15393 22457 15427 22491
rect 15669 22457 15703 22491
rect 17785 22457 17819 22491
rect 23673 22457 23707 22491
rect 35173 22457 35207 22491
rect 12909 22389 12943 22423
rect 16681 22389 16715 22423
rect 20637 22389 20671 22423
rect 21373 22389 21407 22423
rect 32137 22389 32171 22423
rect 32505 22389 32539 22423
rect 35265 22389 35299 22423
rect 36277 22389 36311 22423
rect 36461 22389 36495 22423
rect 9045 22185 9079 22219
rect 10241 22185 10275 22219
rect 12633 22185 12667 22219
rect 15485 22185 15519 22219
rect 16957 22185 16991 22219
rect 26433 22185 26467 22219
rect 33241 22185 33275 22219
rect 36001 22185 36035 22219
rect 38025 22185 38059 22219
rect 13185 22117 13219 22151
rect 23029 22117 23063 22151
rect 24225 22117 24259 22151
rect 24685 22117 24719 22151
rect 34713 22117 34747 22151
rect 35265 22117 35299 22151
rect 36461 22117 36495 22151
rect 10701 22049 10735 22083
rect 12817 22049 12851 22083
rect 13737 22049 13771 22083
rect 16865 22049 16899 22083
rect 24777 22049 24811 22083
rect 25421 22049 25455 22083
rect 27077 22049 27111 22083
rect 29377 22049 29411 22083
rect 31677 22049 31711 22083
rect 35173 22049 35207 22083
rect 35633 22049 35667 22083
rect 36277 22049 36311 22083
rect 36645 22049 36679 22083
rect 38669 22049 38703 22083
rect 8953 21981 8987 22015
rect 10425 21981 10459 22015
rect 10517 21981 10551 22015
rect 10609 21981 10643 22015
rect 12633 21981 12667 22015
rect 12909 21981 12943 22015
rect 13553 21981 13587 22015
rect 13645 21981 13679 22015
rect 16598 21981 16632 22015
rect 17601 21981 17635 22015
rect 17877 21981 17911 22015
rect 17969 21981 18003 22015
rect 18153 21981 18187 22015
rect 18245 21981 18279 22015
rect 18429 21981 18463 22015
rect 20361 21981 20395 22015
rect 20729 21981 20763 22015
rect 23029 21981 23063 22015
rect 23121 21981 23155 22015
rect 23949 21991 23983 22025
rect 24041 21981 24075 22015
rect 24409 21981 24443 22015
rect 26249 21981 26283 22015
rect 26433 21981 26467 22015
rect 26629 21981 26663 22015
rect 26893 21981 26927 22015
rect 27169 21981 27203 22015
rect 27813 21981 27847 22015
rect 31585 21981 31619 22015
rect 31769 21981 31803 22015
rect 31861 21981 31895 22015
rect 33333 21981 33367 22015
rect 34345 21981 34379 22015
rect 34529 21981 34563 22015
rect 34897 21981 34931 22015
rect 35081 21981 35115 22015
rect 35446 21975 35480 22009
rect 36553 21981 36587 22015
rect 38117 21981 38151 22015
rect 19257 21913 19291 21947
rect 20085 21913 20119 21947
rect 23305 21913 23339 21947
rect 24225 21913 24259 21947
rect 24685 21913 24719 21947
rect 27261 21913 27295 21947
rect 29132 21913 29166 21947
rect 32128 21913 32162 21947
rect 34069 21913 34103 21947
rect 34437 21913 34471 21947
rect 35985 21913 36019 21947
rect 36185 21913 36219 21947
rect 36912 21913 36946 21947
rect 13093 21845 13127 21879
rect 17693 21845 17727 21879
rect 19073 21845 19107 21879
rect 22155 21845 22189 21879
rect 24501 21845 24535 21879
rect 25697 21845 25731 21879
rect 26709 21845 26743 21879
rect 27997 21845 28031 21879
rect 35817 21845 35851 21879
rect 36277 21845 36311 21879
rect 9229 21641 9263 21675
rect 9689 21641 9723 21675
rect 18337 21641 18371 21675
rect 24133 21641 24167 21675
rect 28641 21641 28675 21675
rect 29469 21641 29503 21675
rect 34805 21641 34839 21675
rect 35081 21641 35115 21675
rect 11345 21573 11379 21607
rect 11805 21573 11839 21607
rect 11897 21573 11931 21607
rect 20913 21573 20947 21607
rect 27528 21573 27562 21607
rect 35449 21573 35483 21607
rect 36737 21573 36771 21607
rect 36921 21573 36955 21607
rect 8677 21505 8711 21539
rect 9597 21505 9631 21539
rect 10977 21505 11011 21539
rect 11161 21505 11195 21539
rect 11713 21505 11747 21539
rect 12015 21505 12049 21539
rect 12173 21505 12207 21539
rect 13369 21505 13403 21539
rect 13829 21505 13863 21539
rect 14013 21505 14047 21539
rect 17509 21505 17543 21539
rect 17693 21505 17727 21539
rect 19450 21505 19484 21539
rect 19717 21505 19751 21539
rect 23489 21505 23523 21539
rect 25513 21505 25547 21539
rect 25605 21505 25639 21539
rect 25789 21505 25823 21539
rect 27261 21505 27295 21539
rect 29653 21505 29687 21539
rect 30950 21505 30984 21539
rect 33425 21505 33459 21539
rect 33692 21505 33726 21539
rect 36645 21505 36679 21539
rect 9781 21437 9815 21471
rect 12633 21437 12667 21471
rect 20729 21437 20763 21471
rect 23673 21437 23707 21471
rect 24777 21437 24811 21471
rect 25881 21437 25915 21471
rect 26433 21437 26467 21471
rect 29285 21437 29319 21471
rect 31217 21437 31251 21471
rect 35541 21437 35575 21471
rect 35725 21437 35759 21471
rect 25329 21369 25363 21403
rect 36921 21369 36955 21403
rect 8493 21301 8527 21335
rect 11529 21301 11563 21335
rect 13921 21301 13955 21335
rect 17325 21301 17359 21335
rect 18245 21301 18279 21335
rect 20085 21301 20119 21335
rect 21005 21301 21039 21335
rect 23305 21301 23339 21335
rect 25789 21301 25823 21335
rect 28733 21301 28767 21335
rect 29837 21301 29871 21335
rect 17693 21097 17727 21131
rect 24225 21097 24259 21131
rect 27813 21097 27847 21131
rect 28181 21097 28215 21131
rect 29377 21097 29411 21131
rect 30205 21097 30239 21131
rect 34253 21097 34287 21131
rect 28365 21029 28399 21063
rect 32781 21029 32815 21063
rect 8953 20961 8987 20995
rect 10977 20961 11011 20995
rect 14105 20961 14139 20995
rect 14473 20961 14507 20995
rect 33425 20961 33459 20995
rect 35541 20961 35575 20995
rect 8769 20893 8803 20927
rect 11069 20893 11103 20927
rect 11345 20893 11379 20927
rect 11529 20893 11563 20927
rect 11897 20893 11931 20927
rect 12081 20893 12115 20927
rect 12265 20893 12299 20927
rect 12367 20903 12401 20937
rect 13369 20893 13403 20927
rect 17334 20893 17368 20927
rect 17601 20893 17635 20927
rect 19073 20893 19107 20927
rect 19257 20893 19291 20927
rect 19533 20893 19567 20927
rect 21005 20893 21039 20927
rect 22845 20893 22879 20927
rect 24593 20893 24627 20927
rect 24685 20893 24719 20927
rect 26074 20893 26108 20927
rect 26341 20893 26375 20927
rect 26433 20893 26467 20927
rect 26700 20893 26734 20927
rect 28273 20893 28307 20927
rect 28641 20893 28675 20927
rect 28733 20893 28767 20927
rect 29193 20893 29227 20927
rect 29653 20893 29687 20927
rect 30665 20893 30699 20927
rect 31401 20893 31435 20927
rect 33885 20893 33919 20927
rect 33977 20893 34011 20927
rect 34161 20893 34195 20927
rect 34437 20893 34471 20927
rect 35081 20893 35115 20927
rect 35265 20893 35299 20927
rect 37197 20893 37231 20927
rect 38577 20893 38611 20927
rect 30159 20859 30193 20893
rect 10701 20825 10735 20859
rect 11207 20825 11241 20859
rect 11437 20825 11471 20859
rect 12541 20825 12575 20859
rect 18806 20825 18840 20859
rect 19800 20825 19834 20859
rect 21272 20825 21306 20859
rect 23112 20825 23146 20859
rect 30389 20825 30423 20859
rect 31668 20825 31702 20859
rect 34897 20825 34931 20859
rect 35173 20825 35207 20859
rect 35383 20825 35417 20859
rect 8677 20757 8711 20791
rect 11713 20757 11747 20791
rect 15899 20757 15933 20791
rect 16221 20757 16255 20791
rect 19349 20757 19383 20791
rect 20913 20757 20947 20791
rect 22385 20757 22419 20791
rect 24409 20757 24443 20791
rect 24961 20757 24995 20791
rect 27905 20757 27939 20791
rect 28549 20757 28583 20791
rect 28825 20757 28859 20791
rect 29745 20757 29779 20791
rect 30021 20757 30055 20791
rect 30573 20757 30607 20791
rect 32873 20757 32907 20791
rect 37841 20757 37875 20791
rect 37933 20757 37967 20791
rect 10977 20553 11011 20587
rect 11345 20553 11379 20587
rect 11713 20553 11747 20587
rect 12357 20553 12391 20587
rect 14749 20553 14783 20587
rect 18245 20553 18279 20587
rect 19993 20553 20027 20587
rect 23029 20553 23063 20587
rect 24685 20553 24719 20587
rect 26157 20553 26191 20587
rect 27721 20553 27755 20587
rect 30021 20553 30055 20587
rect 32137 20553 32171 20587
rect 35173 20553 35207 20587
rect 35909 20553 35943 20587
rect 36829 20553 36863 20587
rect 38669 20553 38703 20587
rect 8217 20485 8251 20519
rect 9965 20485 9999 20519
rect 11253 20485 11287 20519
rect 16313 20485 16347 20519
rect 17785 20485 17819 20519
rect 28457 20485 28491 20519
rect 37556 20485 37590 20519
rect 10425 20417 10459 20451
rect 11069 20417 11103 20451
rect 11345 20417 11379 20451
rect 11621 20417 11655 20451
rect 11805 20417 11839 20451
rect 12449 20417 12483 20451
rect 13001 20417 13035 20451
rect 13461 20417 13495 20451
rect 13553 20417 13587 20451
rect 13921 20417 13955 20451
rect 14013 20417 14047 20451
rect 14657 20417 14691 20451
rect 15393 20417 15427 20451
rect 15669 20417 15703 20451
rect 15945 20417 15979 20451
rect 16037 20417 16071 20451
rect 16221 20417 16255 20451
rect 16405 20417 16439 20451
rect 16681 20417 16715 20451
rect 17601 20417 17635 20451
rect 17877 20417 17911 20451
rect 17969 20417 18003 20451
rect 18429 20417 18463 20451
rect 18613 20417 18647 20451
rect 20269 20417 20303 20451
rect 20821 20417 20855 20451
rect 22293 20417 22327 20451
rect 23305 20417 23339 20451
rect 23397 20417 23431 20451
rect 23489 20417 23523 20451
rect 23765 20417 23799 20451
rect 24777 20417 24811 20451
rect 25033 20417 25067 20451
rect 28273 20417 28307 20451
rect 28733 20417 28767 20451
rect 29929 20417 29963 20451
rect 30113 20417 30147 20451
rect 30849 20417 30883 20451
rect 31033 20417 31067 20451
rect 31401 20417 31435 20451
rect 31585 20417 31619 20451
rect 31677 20417 31711 20451
rect 33701 20417 33735 20451
rect 33885 20417 33919 20451
rect 35089 20417 35123 20451
rect 35265 20417 35299 20451
rect 35541 20417 35575 20451
rect 35725 20417 35759 20451
rect 35820 20417 35854 20451
rect 36093 20417 36127 20451
rect 36185 20417 36219 20451
rect 36333 20417 36367 20451
rect 36461 20417 36495 20451
rect 36553 20417 36587 20451
rect 36691 20417 36725 20451
rect 7941 20349 7975 20383
rect 11989 20349 12023 20383
rect 12541 20349 12575 20383
rect 13645 20349 13679 20383
rect 13737 20349 13771 20383
rect 17233 20349 17267 20383
rect 20177 20349 20211 20383
rect 20637 20349 20671 20383
rect 23213 20349 23247 20383
rect 24133 20349 24167 20383
rect 31861 20349 31895 20383
rect 32689 20349 32723 20383
rect 33977 20349 34011 20383
rect 35633 20349 35667 20383
rect 37289 20349 37323 20383
rect 12173 20281 12207 20315
rect 18153 20281 18187 20315
rect 21373 20281 21407 20315
rect 23949 20281 23983 20315
rect 28641 20281 28675 20315
rect 31033 20281 31067 20315
rect 31493 20281 31527 20315
rect 12725 20213 12759 20247
rect 13277 20213 13311 20247
rect 14105 20213 14139 20247
rect 15209 20213 15243 20247
rect 15577 20213 15611 20247
rect 15761 20213 15795 20247
rect 22477 20213 22511 20247
rect 28549 20213 28583 20247
rect 33517 20213 33551 20247
rect 36093 20213 36127 20247
rect 9597 20009 9631 20043
rect 17049 20009 17083 20043
rect 22477 20009 22511 20043
rect 22569 20009 22603 20043
rect 23029 20009 23063 20043
rect 23765 20009 23799 20043
rect 29101 20009 29135 20043
rect 35265 20009 35299 20043
rect 35541 20009 35575 20043
rect 35909 20009 35943 20043
rect 28917 19941 28951 19975
rect 10609 19873 10643 19907
rect 15301 19873 15335 19907
rect 15577 19873 15611 19907
rect 21833 19873 21867 19907
rect 23857 19873 23891 19907
rect 24685 19873 24719 19907
rect 25237 19873 25271 19907
rect 27537 19873 27571 19907
rect 30113 19873 30147 19907
rect 30297 19873 30331 19907
rect 37197 19873 37231 19907
rect 9505 19805 9539 19839
rect 12633 19805 12667 19839
rect 20545 19805 20579 19839
rect 20729 19805 20763 19839
rect 22201 19805 22235 19839
rect 22293 19805 22327 19839
rect 22753 19805 22787 19839
rect 22845 19805 22879 19839
rect 23121 19805 23155 19839
rect 23581 19805 23615 19839
rect 23765 19805 23799 19839
rect 24041 19805 24075 19839
rect 24225 19805 24259 19839
rect 24409 19805 24443 19839
rect 27804 19805 27838 19839
rect 29285 19805 29319 19839
rect 29377 19805 29411 19839
rect 30481 19805 30515 19839
rect 30573 19805 30607 19839
rect 32045 19805 32079 19839
rect 34345 19805 34379 19839
rect 35081 19805 35115 19839
rect 36553 19805 36587 19839
rect 10885 19737 10919 19771
rect 12817 19737 12851 19771
rect 13001 19737 13035 19771
rect 21971 19737 22005 19771
rect 22109 19737 22143 19771
rect 29101 19737 29135 19771
rect 29561 19737 29595 19771
rect 30665 19737 30699 19771
rect 32312 19737 32346 19771
rect 33701 19737 33735 19771
rect 34713 19737 34747 19771
rect 34989 19737 35023 19771
rect 35725 19737 35759 19771
rect 20637 19669 20671 19703
rect 24593 19669 24627 19703
rect 30849 19669 30883 19703
rect 33425 19669 33459 19703
rect 34897 19669 34931 19703
rect 35357 19669 35391 19703
rect 35525 19669 35559 19703
rect 36645 19669 36679 19703
rect 11713 19465 11747 19499
rect 13093 19465 13127 19499
rect 16405 19465 16439 19499
rect 18521 19465 18555 19499
rect 21373 19465 21407 19499
rect 23213 19465 23247 19499
rect 32781 19465 32815 19499
rect 37013 19465 37047 19499
rect 15393 19397 15427 19431
rect 22078 19397 22112 19431
rect 27077 19397 27111 19431
rect 27629 19397 27663 19431
rect 31697 19397 31731 19431
rect 33057 19397 33091 19431
rect 34957 19397 34991 19431
rect 35173 19397 35207 19431
rect 35265 19397 35299 19431
rect 11621 19329 11655 19363
rect 13461 19329 13495 19363
rect 13553 19329 13587 19363
rect 14473 19329 14507 19363
rect 15669 19329 15703 19363
rect 16313 19329 16347 19363
rect 17316 19329 17350 19363
rect 19645 19329 19679 19363
rect 19901 19329 19935 19363
rect 20269 19329 20303 19363
rect 20545 19329 20579 19363
rect 20821 19329 20855 19363
rect 21005 19329 21039 19363
rect 21097 19329 21131 19363
rect 21189 19329 21223 19363
rect 21465 19329 21499 19363
rect 21649 19329 21683 19363
rect 21833 19329 21867 19363
rect 23489 19329 23523 19363
rect 25062 19329 25096 19363
rect 25329 19329 25363 19363
rect 25421 19329 25455 19363
rect 25688 19329 25722 19363
rect 29745 19329 29779 19363
rect 29929 19329 29963 19363
rect 30205 19329 30239 19363
rect 30481 19329 30515 19363
rect 31953 19329 31987 19363
rect 32597 19329 32631 19363
rect 32873 19329 32907 19363
rect 32965 19329 32999 19363
rect 33241 19329 33275 19363
rect 34069 19329 34103 19363
rect 35541 19329 35575 19363
rect 35633 19329 35667 19363
rect 35889 19329 35923 19363
rect 13737 19261 13771 19295
rect 17049 19261 17083 19295
rect 30113 19261 30147 19295
rect 33885 19261 33919 19295
rect 34621 19261 34655 19295
rect 21649 19193 21683 19227
rect 32597 19193 32631 19227
rect 33241 19193 33275 19227
rect 35449 19193 35483 19227
rect 35541 19193 35575 19227
rect 14381 19125 14415 19159
rect 18429 19125 18463 19159
rect 23581 19125 23615 19159
rect 23949 19125 23983 19159
rect 26801 19125 26835 19159
rect 27169 19125 27203 19159
rect 27721 19125 27755 19159
rect 30573 19125 30607 19159
rect 33333 19125 33367 19159
rect 34805 19125 34839 19159
rect 34989 19125 35023 19159
rect 14933 18921 14967 18955
rect 19993 18921 20027 18955
rect 25973 18921 26007 18955
rect 30481 18921 30515 18955
rect 31953 18921 31987 18955
rect 34345 18921 34379 18955
rect 13737 18853 13771 18887
rect 21649 18853 21683 18887
rect 28733 18853 28767 18887
rect 30665 18853 30699 18887
rect 31585 18853 31619 18887
rect 32781 18853 32815 18887
rect 34989 18853 35023 18887
rect 12725 18785 12759 18819
rect 13093 18785 13127 18819
rect 13553 18785 13587 18819
rect 13645 18785 13679 18819
rect 15577 18785 15611 18819
rect 18889 18785 18923 18819
rect 19901 18785 19935 18819
rect 22109 18785 22143 18819
rect 22293 18785 22327 18819
rect 23581 18785 23615 18819
rect 23765 18785 23799 18819
rect 24133 18785 24167 18819
rect 28365 18785 28399 18819
rect 28549 18785 28583 18819
rect 30757 18785 30791 18819
rect 32597 18785 32631 18819
rect 32965 18785 32999 18819
rect 9597 18717 9631 18751
rect 10609 18717 10643 18751
rect 11069 18717 11103 18751
rect 11529 18717 11563 18751
rect 12909 18717 12943 18751
rect 13369 18717 13403 18751
rect 13737 18717 13771 18751
rect 13921 18717 13955 18751
rect 15301 18717 15335 18751
rect 15393 18717 15427 18751
rect 17417 18717 17451 18751
rect 18061 18717 18095 18751
rect 19257 18717 19291 18751
rect 20177 18717 20211 18751
rect 20269 18717 20303 18751
rect 20361 18717 20395 18751
rect 20637 18717 20671 18751
rect 20729 18717 20763 18751
rect 20913 18717 20947 18751
rect 22017 18717 22051 18751
rect 22937 18717 22971 18751
rect 23121 18717 23155 18751
rect 23213 18717 23247 18751
rect 23397 18717 23431 18751
rect 23673 18717 23707 18751
rect 23949 18717 23983 18751
rect 25789 18717 25823 18751
rect 25973 18717 26007 18751
rect 26065 18717 26099 18751
rect 26617 18717 26651 18751
rect 26893 18717 26927 18751
rect 28641 18717 28675 18751
rect 29009 18717 29043 18751
rect 30113 18717 30147 18751
rect 31401 18717 31435 18751
rect 31493 18717 31527 18751
rect 31769 18717 31803 18751
rect 32873 18717 32907 18751
rect 34805 18717 34839 18751
rect 37197 18717 37231 18751
rect 37473 18717 37507 18751
rect 37657 18717 37691 18751
rect 37933 18717 37967 18751
rect 38485 18717 38519 18751
rect 17172 18649 17206 18683
rect 17509 18649 17543 18683
rect 20479 18649 20513 18683
rect 23029 18649 23063 18683
rect 28365 18649 28399 18683
rect 28733 18649 28767 18683
rect 30297 18649 30331 18683
rect 33210 18649 33244 18683
rect 9505 18581 9539 18615
rect 10425 18581 10459 18615
rect 10977 18581 11011 18615
rect 12173 18581 12207 18615
rect 13185 18581 13219 18615
rect 16037 18581 16071 18615
rect 18337 18581 18371 18615
rect 20821 18581 20855 18615
rect 26985 18581 27019 18615
rect 28917 18581 28951 18615
rect 29561 18581 29595 18615
rect 30497 18581 30531 18615
rect 32873 18581 32907 18615
rect 37013 18581 37047 18615
rect 11345 18377 11379 18411
rect 17509 18377 17543 18411
rect 19533 18377 19567 18411
rect 22661 18377 22695 18411
rect 29193 18377 29227 18411
rect 29561 18377 29595 18411
rect 9873 18309 9907 18343
rect 13461 18309 13495 18343
rect 15209 18309 15243 18343
rect 18245 18309 18279 18343
rect 20085 18309 20119 18343
rect 21189 18309 21223 18343
rect 23305 18309 23339 18343
rect 25053 18309 25087 18343
rect 28080 18309 28114 18343
rect 30696 18309 30730 18343
rect 31033 18309 31067 18343
rect 36645 18309 36679 18343
rect 37534 18309 37568 18343
rect 7757 18241 7791 18275
rect 9597 18241 9631 18275
rect 11529 18241 11563 18275
rect 11713 18241 11747 18275
rect 13185 18241 13219 18275
rect 17693 18241 17727 18275
rect 17785 18241 17819 18275
rect 17877 18241 17911 18275
rect 17995 18241 18029 18275
rect 18153 18241 18187 18275
rect 18429 18241 18463 18275
rect 18521 18241 18555 18275
rect 18705 18241 18739 18275
rect 18797 18241 18831 18275
rect 19993 18241 20027 18275
rect 20453 18241 20487 18275
rect 21465 18241 21499 18275
rect 21925 18241 21959 18275
rect 22569 18241 22603 18275
rect 23029 18241 23063 18275
rect 25513 18241 25547 18275
rect 25789 18241 25823 18275
rect 25881 18241 25915 18275
rect 26065 18241 26099 18275
rect 26985 18241 27019 18275
rect 27813 18241 27847 18275
rect 30941 18241 30975 18275
rect 35081 18241 35115 18275
rect 35173 18241 35207 18275
rect 35357 18241 35391 18275
rect 35449 18241 35483 18275
rect 36369 18241 36403 18275
rect 36462 18241 36496 18275
rect 36737 18241 36771 18275
rect 36873 18241 36907 18275
rect 37289 18241 37323 18275
rect 8033 18173 8067 18207
rect 17233 18173 17267 18207
rect 18981 18173 19015 18207
rect 20177 18173 20211 18207
rect 21557 18173 21591 18207
rect 27629 18173 27663 18207
rect 31585 18173 31619 18207
rect 19625 18105 19659 18139
rect 26065 18105 26099 18139
rect 37013 18105 37047 18139
rect 9505 18037 9539 18071
rect 11621 18037 11655 18071
rect 16681 18037 16715 18071
rect 22201 18037 22235 18071
rect 25329 18037 25363 18071
rect 34897 18037 34931 18071
rect 38669 18037 38703 18071
rect 8953 17833 8987 17867
rect 10517 17833 10551 17867
rect 13139 17833 13173 17867
rect 20729 17833 20763 17867
rect 24501 17833 24535 17867
rect 26525 17833 26559 17867
rect 30849 17833 30883 17867
rect 33701 17833 33735 17867
rect 38117 17833 38151 17867
rect 38301 17833 38335 17867
rect 19901 17765 19935 17799
rect 32873 17765 32907 17799
rect 36093 17765 36127 17799
rect 11161 17697 11195 17731
rect 11345 17697 11379 17731
rect 11713 17697 11747 17731
rect 15117 17697 15151 17731
rect 19441 17697 19475 17731
rect 21373 17697 21407 17731
rect 21833 17697 21867 17731
rect 22937 17697 22971 17731
rect 23581 17697 23615 17731
rect 30389 17697 30423 17731
rect 30573 17697 30607 17731
rect 32965 17697 32999 17731
rect 9137 17629 9171 17663
rect 17969 17629 18003 17663
rect 18245 17629 18279 17663
rect 22017 17629 22051 17663
rect 22477 17629 22511 17663
rect 22845 17629 22879 17663
rect 23673 17629 23707 17663
rect 24409 17629 24443 17663
rect 25145 17629 25179 17663
rect 25412 17629 25446 17663
rect 27997 17629 28031 17663
rect 28273 17629 28307 17663
rect 30757 17629 30791 17663
rect 30849 17629 30883 17663
rect 31217 17629 31251 17663
rect 31401 17629 31435 17663
rect 31493 17629 31527 17663
rect 33885 17629 33919 17663
rect 33977 17629 34011 17663
rect 34713 17629 34747 17663
rect 36277 17629 36311 17663
rect 36829 17629 36863 17663
rect 37105 17629 37139 17663
rect 37197 17629 37231 17663
rect 37841 17629 37875 17663
rect 15384 17561 15418 17595
rect 17724 17561 17758 17595
rect 19349 17561 19383 17595
rect 22569 17561 22603 17595
rect 22661 17561 22695 17595
rect 23949 17561 23983 17595
rect 27752 17561 27786 17595
rect 31309 17561 31343 17595
rect 31738 17561 31772 17595
rect 33701 17561 33735 17595
rect 34958 17561 34992 17595
rect 36553 17561 36587 17595
rect 37933 17561 37967 17595
rect 10885 17493 10919 17527
rect 10977 17493 11011 17527
rect 16497 17493 16531 17527
rect 16589 17493 16623 17527
rect 18061 17493 18095 17527
rect 19441 17493 19475 17527
rect 21097 17493 21131 17527
rect 21189 17493 21223 17527
rect 22201 17493 22235 17527
rect 22293 17493 22327 17527
rect 26617 17493 26651 17527
rect 28089 17493 28123 17527
rect 29837 17493 29871 17527
rect 33609 17493 33643 17527
rect 38133 17493 38167 17527
rect 13185 17289 13219 17323
rect 15301 17289 15335 17323
rect 15662 17289 15696 17323
rect 18981 17289 19015 17323
rect 19073 17289 19107 17323
rect 24593 17289 24627 17323
rect 25789 17289 25823 17323
rect 26801 17289 26835 17323
rect 29745 17289 29779 17323
rect 32413 17289 32447 17323
rect 34713 17289 34747 17323
rect 35909 17289 35943 17323
rect 19257 17255 19291 17289
rect 9873 17221 9907 17255
rect 23121 17221 23155 17255
rect 25605 17221 25639 17255
rect 29929 17221 29963 17255
rect 32229 17221 32263 17255
rect 33885 17221 33919 17255
rect 38025 17221 38059 17255
rect 7481 17153 7515 17187
rect 9781 17153 9815 17187
rect 12357 17153 12391 17187
rect 13277 17153 13311 17187
rect 14861 17153 14895 17187
rect 15117 17153 15151 17187
rect 15209 17153 15243 17187
rect 15393 17153 15427 17187
rect 15485 17153 15519 17187
rect 15577 17153 15611 17187
rect 15761 17153 15795 17187
rect 17233 17153 17267 17187
rect 17868 17153 17902 17187
rect 19254 17153 19288 17187
rect 20545 17153 20579 17187
rect 21833 17153 21867 17187
rect 22385 17153 22419 17187
rect 26617 17153 26651 17187
rect 26985 17153 27019 17187
rect 29653 17153 29687 17187
rect 32137 17153 32171 17187
rect 34897 17153 34931 17187
rect 35173 17153 35207 17187
rect 35357 17153 35391 17187
rect 35817 17153 35851 17187
rect 36093 17153 36127 17187
rect 37289 17153 37323 17187
rect 38209 17153 38243 17187
rect 38301 17153 38335 17187
rect 7757 17085 7791 17119
rect 9965 17085 9999 17119
rect 10793 17085 10827 17119
rect 13001 17085 13035 17119
rect 16405 17085 16439 17119
rect 16681 17085 16715 17119
rect 17601 17085 17635 17119
rect 19717 17085 19751 17119
rect 21281 17085 21315 17119
rect 22109 17085 22143 17119
rect 26433 17085 26467 17119
rect 27905 17085 27939 17119
rect 34161 17085 34195 17119
rect 36185 17085 36219 17119
rect 36829 17085 36863 17119
rect 37933 17085 37967 17119
rect 9413 17017 9447 17051
rect 13737 17017 13771 17051
rect 19993 17017 20027 17051
rect 21925 17017 21959 17051
rect 25237 17017 25271 17051
rect 29929 17017 29963 17051
rect 36093 17017 36127 17051
rect 9229 16949 9263 16983
rect 10241 16949 10275 16983
rect 15853 16949 15887 16983
rect 19625 16949 19659 16983
rect 20729 16949 20763 16983
rect 22017 16949 22051 16983
rect 23029 16949 23063 16983
rect 25605 16949 25639 16983
rect 27629 16949 27663 16983
rect 28549 16949 28583 16983
rect 38117 16949 38151 16983
rect 8585 16745 8619 16779
rect 9597 16745 9631 16779
rect 15209 16745 15243 16779
rect 17969 16745 18003 16779
rect 26341 16745 26375 16779
rect 37565 16745 37599 16779
rect 9505 16677 9539 16711
rect 19349 16677 19383 16711
rect 29929 16677 29963 16711
rect 11253 16609 11287 16643
rect 13921 16609 13955 16643
rect 16589 16609 16623 16643
rect 16773 16609 16807 16643
rect 17877 16609 17911 16643
rect 18981 16609 19015 16643
rect 19717 16609 19751 16643
rect 19809 16609 19843 16643
rect 25145 16609 25179 16643
rect 25329 16609 25363 16643
rect 27997 16609 28031 16643
rect 31401 16609 31435 16643
rect 32321 16609 32355 16643
rect 36185 16609 36219 16643
rect 8493 16541 8527 16575
rect 9229 16541 9263 16575
rect 9781 16541 9815 16575
rect 10149 16541 10183 16575
rect 11437 16541 11471 16575
rect 11713 16541 11747 16575
rect 11890 16541 11924 16575
rect 12265 16541 12299 16575
rect 14105 16541 14139 16575
rect 14749 16541 14783 16575
rect 14933 16541 14967 16575
rect 15025 16541 15059 16575
rect 15209 16541 15243 16575
rect 15301 16541 15335 16575
rect 15945 16541 15979 16575
rect 17417 16541 17451 16575
rect 17509 16541 17543 16575
rect 17693 16541 17727 16575
rect 18153 16541 18187 16575
rect 18889 16541 18923 16575
rect 19073 16541 19107 16575
rect 19533 16541 19567 16575
rect 21373 16541 21407 16575
rect 22845 16541 22879 16575
rect 23112 16541 23146 16575
rect 25237 16541 25271 16575
rect 25789 16541 25823 16575
rect 25881 16541 25915 16575
rect 26065 16541 26099 16575
rect 26157 16541 26191 16575
rect 26985 16541 27019 16575
rect 27813 16541 27847 16575
rect 29653 16541 29687 16575
rect 29837 16541 29871 16575
rect 29929 16541 29963 16575
rect 31134 16541 31168 16575
rect 36452 16541 36486 16575
rect 9505 16473 9539 16507
rect 9873 16473 9907 16507
rect 9965 16473 9999 16507
rect 10241 16473 10275 16507
rect 10425 16473 10459 16507
rect 11805 16473 11839 16507
rect 13676 16473 13710 16507
rect 20054 16473 20088 16507
rect 21640 16473 21674 16507
rect 27261 16473 27295 16507
rect 28264 16473 28298 16507
rect 33149 16473 33183 16507
rect 9321 16405 9355 16439
rect 10609 16405 10643 16439
rect 11621 16405 11655 16439
rect 12449 16405 12483 16439
rect 12541 16405 12575 16439
rect 14197 16405 14231 16439
rect 14841 16405 14875 16439
rect 16037 16405 16071 16439
rect 21189 16405 21223 16439
rect 22753 16405 22787 16439
rect 24225 16405 24259 16439
rect 24961 16405 24995 16439
rect 26433 16405 26467 16439
rect 29377 16405 29411 16439
rect 30021 16405 30055 16439
rect 9689 16201 9723 16235
rect 11989 16201 12023 16235
rect 15117 16201 15151 16235
rect 16497 16201 16531 16235
rect 18981 16201 19015 16235
rect 20637 16201 20671 16235
rect 21833 16201 21867 16235
rect 26985 16201 27019 16235
rect 28549 16201 28583 16235
rect 34805 16201 34839 16235
rect 35357 16201 35391 16235
rect 9841 16133 9875 16167
rect 10057 16133 10091 16167
rect 17969 16133 18003 16167
rect 19165 16133 19199 16167
rect 25114 16133 25148 16167
rect 30297 16133 30331 16167
rect 30573 16133 30607 16167
rect 10793 16065 10827 16099
rect 10885 16065 10919 16099
rect 11069 16065 11103 16099
rect 11161 16065 11195 16099
rect 12265 16065 12299 16099
rect 12357 16065 12391 16099
rect 12541 16065 12575 16099
rect 12725 16065 12759 16099
rect 13185 16065 13219 16099
rect 13277 16065 13311 16099
rect 15117 16065 15151 16099
rect 16313 16065 16347 16099
rect 17601 16065 17635 16099
rect 17877 16065 17911 16099
rect 18061 16065 18095 16099
rect 18889 16065 18923 16099
rect 19257 16065 19291 16099
rect 19513 16065 19547 16099
rect 20729 16065 20763 16099
rect 20913 16065 20947 16099
rect 21557 16065 21591 16099
rect 22385 16065 22419 16099
rect 23121 16065 23155 16099
rect 28109 16065 28143 16099
rect 28365 16065 28399 16099
rect 28457 16065 28491 16099
rect 28641 16065 28675 16099
rect 30389 16065 30423 16099
rect 30665 16065 30699 16099
rect 30757 16065 30791 16099
rect 30941 16065 30975 16099
rect 32321 16065 32355 16099
rect 33425 16065 33459 16099
rect 33692 16065 33726 16099
rect 34897 16065 34931 16099
rect 35416 16065 35450 16099
rect 12081 15997 12115 16031
rect 14841 15997 14875 16031
rect 15761 15997 15795 16031
rect 16129 15997 16163 16031
rect 16681 15997 16715 16031
rect 17785 15997 17819 16031
rect 23949 15997 23983 16031
rect 24869 15997 24903 16031
rect 29745 15997 29779 16031
rect 32597 15997 32631 16031
rect 32689 15997 32723 16031
rect 33333 15997 33367 16031
rect 11989 15929 12023 15963
rect 15025 15929 15059 15963
rect 19165 15929 19199 15963
rect 21005 15929 21039 15963
rect 30389 15929 30423 15963
rect 35541 15929 35575 15963
rect 9873 15861 9907 15895
rect 11345 15861 11379 15895
rect 12173 15861 12207 15895
rect 13737 15861 13771 15895
rect 15209 15861 15243 15895
rect 17325 15861 17359 15895
rect 17417 15861 17451 15895
rect 20729 15861 20763 15895
rect 22569 15861 22603 15895
rect 23397 15861 23431 15895
rect 26249 15861 26283 15895
rect 30757 15861 30791 15895
rect 32137 15861 32171 15895
rect 32505 15861 32539 15895
rect 34989 15861 35023 15895
rect 11621 15657 11655 15691
rect 11989 15657 12023 15691
rect 23213 15657 23247 15691
rect 26893 15657 26927 15691
rect 31493 15657 31527 15691
rect 34161 15657 34195 15691
rect 36369 15657 36403 15691
rect 11161 15589 11195 15623
rect 8769 15521 8803 15555
rect 9597 15521 9631 15555
rect 17601 15521 17635 15555
rect 19257 15521 19291 15555
rect 19901 15521 19935 15555
rect 20361 15521 20395 15555
rect 21189 15521 21223 15555
rect 22017 15521 22051 15555
rect 29929 15521 29963 15555
rect 34989 15521 35023 15555
rect 37013 15521 37047 15555
rect 7021 15453 7055 15487
rect 9965 15453 9999 15487
rect 10149 15453 10183 15487
rect 10977 15453 11011 15487
rect 11069 15453 11103 15487
rect 11253 15453 11287 15487
rect 11345 15453 11379 15487
rect 11621 15453 11655 15487
rect 11805 15453 11839 15487
rect 15218 15453 15252 15487
rect 15485 15453 15519 15487
rect 15853 15453 15887 15487
rect 19073 15453 19107 15487
rect 20177 15453 20211 15487
rect 20269 15453 20303 15487
rect 20453 15453 20487 15487
rect 21558 15453 21592 15487
rect 21741 15453 21775 15487
rect 22109 15453 22143 15487
rect 23029 15453 23063 15487
rect 23213 15453 23247 15487
rect 23305 15453 23339 15487
rect 24133 15453 24167 15487
rect 24409 15453 24443 15487
rect 26341 15453 26375 15487
rect 26709 15453 26743 15487
rect 26985 15453 27019 15487
rect 27813 15453 27847 15487
rect 29745 15453 29779 15487
rect 29837 15453 29871 15487
rect 30021 15453 30055 15487
rect 30297 15453 30331 15487
rect 31033 15453 31067 15487
rect 31309 15453 31343 15487
rect 31769 15453 31803 15487
rect 32036 15453 32070 15487
rect 33793 15453 33827 15487
rect 33977 15453 34011 15487
rect 34161 15453 34195 15487
rect 34253 15453 34287 15487
rect 34713 15453 34747 15487
rect 37381 15453 37415 15487
rect 7297 15385 7331 15419
rect 9413 15385 9447 15419
rect 10057 15385 10091 15419
rect 17356 15385 17390 15419
rect 18828 15385 18862 15419
rect 21649 15385 21683 15419
rect 21879 15385 21913 15419
rect 23397 15385 23431 15419
rect 24654 15385 24688 15419
rect 26525 15385 26559 15419
rect 26617 15385 26651 15419
rect 31125 15385 31159 15419
rect 35256 15385 35290 15419
rect 9045 15317 9079 15351
rect 9505 15317 9539 15351
rect 14105 15317 14139 15351
rect 15761 15317 15795 15351
rect 16221 15317 16255 15351
rect 17693 15317 17727 15351
rect 19993 15317 20027 15351
rect 20637 15317 20671 15351
rect 21373 15317 21407 15351
rect 22753 15317 22787 15351
rect 23581 15317 23615 15351
rect 25789 15317 25823 15351
rect 27629 15317 27663 15351
rect 28457 15317 28491 15351
rect 29561 15317 29595 15351
rect 30941 15317 30975 15351
rect 33149 15317 33183 15351
rect 33241 15317 33275 15351
rect 34345 15317 34379 15351
rect 34805 15317 34839 15351
rect 36461 15317 36495 15351
rect 37289 15317 37323 15351
rect 7941 15113 7975 15147
rect 8585 15113 8619 15147
rect 9689 15113 9723 15147
rect 13277 15113 13311 15147
rect 14197 15113 14231 15147
rect 17693 15113 17727 15147
rect 18705 15113 18739 15147
rect 22017 15113 22051 15147
rect 23489 15113 23523 15147
rect 23765 15113 23799 15147
rect 24409 15113 24443 15147
rect 27629 15113 27663 15147
rect 29469 15113 29503 15147
rect 31861 15113 31895 15147
rect 35357 15113 35391 15147
rect 9857 15045 9891 15079
rect 10057 15045 10091 15079
rect 11529 15045 11563 15079
rect 16497 15045 16531 15079
rect 16865 15045 16899 15079
rect 19993 15045 20027 15079
rect 22354 15045 22388 15079
rect 25145 15045 25179 15079
rect 27813 15045 27847 15079
rect 30481 15045 30515 15079
rect 30686 15045 30720 15079
rect 31033 15045 31067 15079
rect 33250 15045 33284 15079
rect 34345 15045 34379 15079
rect 8125 14977 8159 15011
rect 8677 14977 8711 15011
rect 11713 14977 11747 15011
rect 11805 14977 11839 15011
rect 12081 14977 12115 15011
rect 12541 14977 12575 15011
rect 13093 14977 13127 15011
rect 13553 14977 13587 15011
rect 13737 14977 13771 15011
rect 14289 14977 14323 15011
rect 14565 14977 14599 15011
rect 14657 14977 14691 15011
rect 14841 14977 14875 15011
rect 15025 14977 15059 15011
rect 15853 14977 15887 15011
rect 16681 14977 16715 15011
rect 16957 14977 16991 15011
rect 18521 14977 18555 15011
rect 18981 14977 19015 15011
rect 19165 14977 19199 15011
rect 20269 14977 20303 15011
rect 20453 14977 20487 15011
rect 20545 14977 20579 15011
rect 20729 14977 20763 15011
rect 21833 14977 21867 15011
rect 22109 14977 22143 15011
rect 23706 14977 23740 15011
rect 24133 14977 24167 15011
rect 24225 14977 24259 15011
rect 24317 14977 24351 15011
rect 24501 14977 24535 15011
rect 24777 14977 24811 15011
rect 27261 14977 27295 15011
rect 27537 14977 27571 15011
rect 28089 14977 28123 15011
rect 28345 14977 28379 15011
rect 30941 14977 30975 15011
rect 31125 14977 31159 15011
rect 31217 14977 31251 15011
rect 31401 14977 31435 15011
rect 31493 14977 31527 15011
rect 31585 14977 31619 15011
rect 33517 14977 33551 15011
rect 33609 14977 33643 15011
rect 35541 14977 35575 15011
rect 35633 14977 35667 15011
rect 35817 14977 35851 15011
rect 35909 14977 35943 15011
rect 12817 14909 12851 14943
rect 13461 14909 13495 14943
rect 13645 14909 13679 14943
rect 15669 14909 15703 14943
rect 17049 14909 17083 14943
rect 18797 14909 18831 14943
rect 19257 14909 19291 14943
rect 21465 14909 21499 14943
rect 25053 14909 25087 14943
rect 25697 14909 25731 14943
rect 26709 14909 26743 14943
rect 26985 14909 27019 14943
rect 11989 14841 12023 14875
rect 12633 14841 12667 14875
rect 13001 14841 13035 14875
rect 14749 14841 14783 14875
rect 16681 14841 16715 14875
rect 20177 14841 20211 14875
rect 20821 14841 20855 14875
rect 23581 14841 23615 14875
rect 24593 14841 24627 14875
rect 24961 14841 24995 14875
rect 26157 14841 26191 14875
rect 9873 14773 9907 14807
rect 11805 14773 11839 14807
rect 12265 14773 12299 14807
rect 12909 14773 12943 14807
rect 14381 14773 14415 14807
rect 15117 14773 15151 14807
rect 19901 14773 19935 14807
rect 20085 14773 20119 14807
rect 27077 14773 27111 14807
rect 27445 14773 27479 14807
rect 27813 14773 27847 14807
rect 30665 14773 30699 14807
rect 30849 14773 30883 14807
rect 32137 14773 32171 14807
rect 13277 14569 13311 14603
rect 15945 14569 15979 14603
rect 16681 14569 16715 14603
rect 19257 14569 19291 14603
rect 21189 14569 21223 14603
rect 31769 14569 31803 14603
rect 12817 14501 12851 14535
rect 19533 14501 19567 14535
rect 19625 14501 19659 14535
rect 28181 14501 28215 14535
rect 10057 14433 10091 14467
rect 11529 14433 11563 14467
rect 12081 14433 12115 14467
rect 14197 14433 14231 14467
rect 16865 14433 16899 14467
rect 17141 14433 17175 14467
rect 20821 14433 20855 14467
rect 23765 14433 23799 14467
rect 24685 14433 24719 14467
rect 25329 14433 25363 14467
rect 27261 14433 27295 14467
rect 27813 14433 27847 14467
rect 9137 14365 9171 14399
rect 9413 14365 9447 14399
rect 10425 14365 10459 14399
rect 10701 14365 10735 14399
rect 11345 14365 11379 14399
rect 12357 14365 12391 14399
rect 12449 14365 12483 14399
rect 12541 14365 12575 14399
rect 13829 14365 13863 14399
rect 14105 14365 14139 14399
rect 14289 14365 14323 14399
rect 14565 14365 14599 14399
rect 16957 14365 16991 14399
rect 17049 14365 17083 14399
rect 18153 14365 18187 14399
rect 19441 14365 19475 14399
rect 19717 14365 19751 14399
rect 19901 14365 19935 14399
rect 19993 14365 20027 14399
rect 22569 14365 22603 14399
rect 23489 14365 23523 14399
rect 26985 14365 27019 14399
rect 27077 14365 27111 14399
rect 27997 14365 28031 14399
rect 28181 14365 28215 14399
rect 30021 14365 30055 14399
rect 31585 14365 31619 14399
rect 32873 14365 32907 14399
rect 34529 14365 34563 14399
rect 10241 14297 10275 14331
rect 12239 14297 12273 14331
rect 12725 14297 12759 14331
rect 13001 14297 13035 14331
rect 13185 14297 13219 14331
rect 14832 14297 14866 14331
rect 22324 14297 22358 14331
rect 25574 14297 25608 14331
rect 33701 14297 33735 14331
rect 8953 14229 8987 14263
rect 9321 14229 9355 14263
rect 9505 14229 9539 14263
rect 10609 14229 10643 14263
rect 11161 14229 11195 14263
rect 17601 14229 17635 14263
rect 25237 14229 25271 14263
rect 26709 14229 26743 14263
rect 29837 14229 29871 14263
rect 34437 14229 34471 14263
rect 9321 14025 9355 14059
rect 10149 14025 10183 14059
rect 11069 14025 11103 14059
rect 17699 14025 17733 14059
rect 18889 14025 18923 14059
rect 21833 14025 21867 14059
rect 23765 14025 23799 14059
rect 25237 14025 25271 14059
rect 26249 14025 26283 14059
rect 10680 13957 10714 13991
rect 10885 13957 10919 13991
rect 12909 13957 12943 13991
rect 17785 13957 17819 13991
rect 17969 13957 18003 13991
rect 20002 13957 20036 13991
rect 22201 13957 22235 13991
rect 29469 13957 29503 13991
rect 31861 13957 31895 13991
rect 7573 13889 7607 13923
rect 10057 13889 10091 13923
rect 10241 13889 10275 13923
rect 10977 13889 11011 13923
rect 12633 13889 12667 13923
rect 15025 13889 15059 13923
rect 15209 13889 15243 13923
rect 17049 13889 17083 13923
rect 17233 13889 17267 13923
rect 17601 13889 17635 13923
rect 17877 13889 17911 13923
rect 20545 13889 20579 13923
rect 22293 13889 22327 13923
rect 23213 13889 23247 13923
rect 24889 13889 24923 13923
rect 25145 13889 25179 13923
rect 25421 13889 25455 13923
rect 25697 13889 25731 13923
rect 26157 13889 26191 13923
rect 26341 13889 26375 13923
rect 26709 13889 26743 13923
rect 26985 13889 27019 13923
rect 27252 13889 27286 13923
rect 29193 13889 29227 13923
rect 31953 13889 31987 13923
rect 32597 13889 32631 13923
rect 33057 13889 33091 13923
rect 35081 13889 35115 13923
rect 36001 13889 36035 13923
rect 36185 13889 36219 13923
rect 18521 13821 18555 13855
rect 20269 13821 20303 13855
rect 20637 13821 20671 13855
rect 22385 13821 22419 13855
rect 23489 13821 23523 13855
rect 25605 13821 25639 13855
rect 26617 13821 26651 13855
rect 30941 13821 30975 13855
rect 31585 13821 31619 13855
rect 32689 13821 32723 13855
rect 34805 13821 34839 13855
rect 35265 13821 35299 13855
rect 35909 13821 35943 13855
rect 10517 13753 10551 13787
rect 14381 13753 14415 13787
rect 15209 13753 15243 13787
rect 25513 13753 25547 13787
rect 7836 13685 7870 13719
rect 10701 13685 10735 13719
rect 17233 13685 17267 13719
rect 28365 13685 28399 13719
rect 31033 13685 31067 13719
rect 33149 13685 33183 13719
rect 33333 13685 33367 13719
rect 36001 13685 36035 13719
rect 8585 13481 8619 13515
rect 10885 13481 10919 13515
rect 12081 13481 12115 13515
rect 12541 13481 12575 13515
rect 13829 13481 13863 13515
rect 17969 13481 18003 13515
rect 22477 13481 22511 13515
rect 30389 13481 30423 13515
rect 30849 13481 30883 13515
rect 33977 13481 34011 13515
rect 34345 13481 34379 13515
rect 34713 13481 34747 13515
rect 11529 13413 11563 13447
rect 11897 13413 11931 13447
rect 30573 13413 30607 13447
rect 34529 13413 34563 13447
rect 9597 13345 9631 13379
rect 11345 13345 11379 13379
rect 15117 13345 15151 13379
rect 20085 13345 20119 13379
rect 23029 13345 23063 13379
rect 26985 13345 27019 13379
rect 28733 13345 28767 13379
rect 29837 13345 29871 13379
rect 32229 13345 32263 13379
rect 36093 13345 36127 13379
rect 8493 13277 8527 13311
rect 9689 13277 9723 13311
rect 9965 13277 9999 13311
rect 10149 13277 10183 13311
rect 10701 13277 10735 13311
rect 11069 13277 11103 13311
rect 11253 13277 11287 13311
rect 11621 13277 11655 13311
rect 12725 13277 12759 13311
rect 12909 13277 12943 13311
rect 13001 13277 13035 13311
rect 13921 13277 13955 13311
rect 16589 13277 16623 13311
rect 16856 13277 16890 13311
rect 18061 13277 18095 13311
rect 18245 13277 18279 13311
rect 20453 13277 20487 13311
rect 27813 13277 27847 13311
rect 30021 13277 30055 13311
rect 30481 13277 30515 13311
rect 30665 13287 30699 13321
rect 30941 13277 30975 13311
rect 35357 13277 35391 13311
rect 35449 13277 35483 13311
rect 35633 13277 35667 13311
rect 36645 13277 36679 13311
rect 36829 13277 36863 13311
rect 10057 13209 10091 13243
rect 11345 13209 11379 13243
rect 12265 13209 12299 13243
rect 15384 13209 15418 13243
rect 22937 13209 22971 13243
rect 32505 13209 32539 13243
rect 34161 13209 34195 13243
rect 34377 13209 34411 13243
rect 35725 13209 35759 13243
rect 35817 13209 35851 13243
rect 35955 13209 35989 13243
rect 36185 13209 36219 13243
rect 36369 13209 36403 13243
rect 9413 13141 9447 13175
rect 12065 13141 12099 13175
rect 16497 13141 16531 13175
rect 18153 13141 18187 13175
rect 21879 13141 21913 13175
rect 22845 13141 22879 13175
rect 28181 13141 28215 13175
rect 29929 13141 29963 13175
rect 36553 13141 36587 13175
rect 36737 13141 36771 13175
rect 11989 12937 12023 12971
rect 20453 12937 20487 12971
rect 21465 12937 21499 12971
rect 24593 12937 24627 12971
rect 24961 12937 24995 12971
rect 27307 12937 27341 12971
rect 32781 12937 32815 12971
rect 8677 12869 8711 12903
rect 11253 12869 11287 12903
rect 12633 12869 12667 12903
rect 12843 12869 12877 12903
rect 14841 12869 14875 12903
rect 17693 12869 17727 12903
rect 23765 12869 23799 12903
rect 26525 12869 26559 12903
rect 30297 12869 30331 12903
rect 30481 12869 30515 12903
rect 30665 12869 30699 12903
rect 31033 12869 31067 12903
rect 35633 12869 35667 12903
rect 8401 12801 8435 12835
rect 11161 12801 11195 12835
rect 11897 12801 11931 12835
rect 12541 12801 12575 12835
rect 12725 12801 12759 12835
rect 14013 12801 14047 12835
rect 16957 12801 16991 12835
rect 17877 12801 17911 12835
rect 17969 12801 18003 12835
rect 18153 12801 18187 12835
rect 18409 12801 18443 12835
rect 20361 12801 20395 12835
rect 20545 12801 20579 12835
rect 20637 12801 20671 12835
rect 21373 12801 21407 12835
rect 23857 12801 23891 12835
rect 25421 12801 25455 12835
rect 25605 12801 25639 12835
rect 26433 12801 26467 12835
rect 28733 12801 28767 12835
rect 29929 12801 29963 12835
rect 30113 12801 30147 12835
rect 30389 12801 30423 12835
rect 30941 12801 30975 12835
rect 31125 12801 31159 12835
rect 31217 12801 31251 12835
rect 31401 12801 31435 12835
rect 32965 12801 32999 12835
rect 34437 12801 34471 12835
rect 35265 12801 35299 12835
rect 10149 12733 10183 12767
rect 12173 12733 12207 12767
rect 13001 12733 13035 12767
rect 13277 12733 13311 12767
rect 13829 12733 13863 12767
rect 20177 12733 20211 12767
rect 21189 12733 21223 12767
rect 21833 12733 21867 12767
rect 22109 12733 22143 12767
rect 23581 12733 23615 12767
rect 25053 12733 25087 12767
rect 25237 12733 25271 12767
rect 26617 12733 26651 12767
rect 29101 12733 29135 12767
rect 29745 12733 29779 12767
rect 34529 12733 34563 12767
rect 34713 12733 34747 12767
rect 35173 12733 35207 12767
rect 35357 12733 35391 12767
rect 37841 12733 37875 12767
rect 17693 12665 17727 12699
rect 19533 12665 19567 12699
rect 26065 12665 26099 12699
rect 34069 12665 34103 12699
rect 11529 12597 11563 12631
rect 12357 12597 12391 12631
rect 17601 12597 17635 12631
rect 19625 12597 19659 12631
rect 25421 12597 25455 12631
rect 29193 12597 29227 12631
rect 30665 12597 30699 12631
rect 31585 12597 31619 12631
rect 34897 12597 34931 12631
rect 35081 12597 35115 12631
rect 37105 12597 37139 12631
rect 37289 12597 37323 12631
rect 9413 12393 9447 12427
rect 13737 12393 13771 12427
rect 22293 12393 22327 12427
rect 26801 12393 26835 12427
rect 29009 12393 29043 12427
rect 31401 12393 31435 12427
rect 34161 12393 34195 12427
rect 34713 12393 34747 12427
rect 35909 12393 35943 12427
rect 36369 12393 36403 12427
rect 17325 12325 17359 12359
rect 11989 12257 12023 12291
rect 12265 12257 12299 12291
rect 19441 12257 19475 12291
rect 19533 12257 19567 12291
rect 22017 12257 22051 12291
rect 22661 12257 22695 12291
rect 22753 12257 22787 12291
rect 22937 12257 22971 12291
rect 25053 12257 25087 12291
rect 28457 12257 28491 12291
rect 9321 12189 9355 12223
rect 10885 12189 10919 12223
rect 17417 12189 17451 12223
rect 17509 12189 17543 12223
rect 17693 12189 17727 12223
rect 19625 12189 19659 12223
rect 20637 12189 20671 12223
rect 21649 12189 21683 12223
rect 21833 12189 21867 12223
rect 22477 12189 22511 12223
rect 22845 12189 22879 12223
rect 23029 12189 23063 12223
rect 24685 12189 24719 12223
rect 24777 12189 24811 12223
rect 27721 12189 27755 12223
rect 28917 12189 28951 12223
rect 29101 12189 29135 12223
rect 30849 12189 30883 12223
rect 31033 12189 31067 12223
rect 31309 12189 31343 12223
rect 31585 12189 31619 12223
rect 31677 12189 31711 12223
rect 32505 12189 32539 12223
rect 32689 12189 32723 12223
rect 33793 12189 33827 12223
rect 33885 12189 33919 12223
rect 34253 12189 34287 12223
rect 34713 12189 34747 12223
rect 34897 12189 34931 12223
rect 35357 12189 35391 12223
rect 35633 12189 35667 12223
rect 35725 12189 35759 12223
rect 36277 12189 36311 12223
rect 21373 12121 21407 12155
rect 25329 12121 25363 12155
rect 35541 12121 35575 12155
rect 10701 12053 10735 12087
rect 17693 12053 17727 12087
rect 19993 12053 20027 12087
rect 24961 12053 24995 12087
rect 31217 12053 31251 12087
rect 31861 12053 31895 12087
rect 32597 12053 32631 12087
rect 33609 12053 33643 12087
rect 13093 11849 13127 11883
rect 17785 11849 17819 11883
rect 23259 11849 23293 11883
rect 25329 11849 25363 11883
rect 26801 11849 26835 11883
rect 27813 11849 27847 11883
rect 30757 11849 30791 11883
rect 32229 11849 32263 11883
rect 33149 11849 33183 11883
rect 33333 11849 33367 11883
rect 34713 11849 34747 11883
rect 35265 11849 35299 11883
rect 15761 11781 15795 11815
rect 17693 11781 17727 11815
rect 19441 11781 19475 11815
rect 21097 11781 21131 11815
rect 21833 11781 21867 11815
rect 27905 11781 27939 11815
rect 31401 11781 31435 11815
rect 33977 11781 34011 11815
rect 11713 11713 11747 11747
rect 13001 11713 13035 11747
rect 16313 11713 16347 11747
rect 17141 11713 17175 11747
rect 17325 11713 17359 11747
rect 19165 11713 19199 11747
rect 21189 11713 21223 11747
rect 22017 11713 22051 11747
rect 22385 11713 22419 11747
rect 22845 11713 22879 11747
rect 25064 11713 25098 11747
rect 25513 11713 25547 11747
rect 25697 11713 25731 11747
rect 25789 11713 25823 11747
rect 26617 11713 26651 11747
rect 27169 11713 27203 11747
rect 27353 11713 27387 11747
rect 28273 11713 28307 11747
rect 29009 11713 29043 11747
rect 31217 11713 31251 11747
rect 31309 11713 31343 11747
rect 31519 11713 31553 11747
rect 32413 11713 32447 11747
rect 32781 11713 32815 11747
rect 32965 11713 32999 11747
rect 33178 11713 33212 11747
rect 33517 11713 33551 11747
rect 34897 11713 34931 11747
rect 35357 11713 35391 11747
rect 14933 11645 14967 11679
rect 17601 11645 17635 11679
rect 22201 11645 22235 11679
rect 22569 11645 22603 11679
rect 22661 11645 22695 11679
rect 24685 11645 24719 11679
rect 28089 11645 28123 11679
rect 28825 11645 28859 11679
rect 29285 11645 29319 11679
rect 31677 11645 31711 11679
rect 33609 11645 33643 11679
rect 35081 11645 35115 11679
rect 22753 11577 22787 11611
rect 27261 11577 27295 11611
rect 27445 11577 27479 11611
rect 11621 11509 11655 11543
rect 16405 11509 16439 11543
rect 16957 11509 16991 11543
rect 18153 11509 18187 11543
rect 20913 11509 20947 11543
rect 23029 11509 23063 11543
rect 31033 11509 31067 11543
rect 32505 11509 32539 11543
rect 32873 11509 32907 11543
rect 33609 11509 33643 11543
rect 10596 11305 10630 11339
rect 18705 11305 18739 11339
rect 19441 11305 19475 11339
rect 19717 11305 19751 11339
rect 21005 11305 21039 11339
rect 23949 11305 23983 11339
rect 29009 11305 29043 11339
rect 30113 11305 30147 11339
rect 31217 11305 31251 11339
rect 31769 11305 31803 11339
rect 34069 11305 34103 11339
rect 19257 11237 19291 11271
rect 32505 11237 32539 11271
rect 10333 11169 10367 11203
rect 15669 11169 15703 11203
rect 20453 11169 20487 11203
rect 27261 11169 27295 11203
rect 27537 11169 27571 11203
rect 32597 11169 32631 11203
rect 32965 11169 32999 11203
rect 33425 11169 33459 11203
rect 35265 11169 35299 11203
rect 12357 11101 12391 11135
rect 15393 11101 15427 11135
rect 17417 11101 17451 11135
rect 18061 11101 18095 11135
rect 18153 11101 18187 11135
rect 18580 11101 18614 11135
rect 19901 11101 19935 11135
rect 20269 11101 20303 11135
rect 20821 11101 20855 11135
rect 21649 11101 21683 11135
rect 21741 11101 21775 11135
rect 23857 11101 23891 11135
rect 25513 11101 25547 11135
rect 25697 11101 25731 11135
rect 25881 11101 25915 11135
rect 29285 11101 29319 11135
rect 30021 11101 30055 11135
rect 31401 11101 31435 11135
rect 31677 11101 31711 11135
rect 31861 11101 31895 11135
rect 32229 11101 32263 11135
rect 32413 11101 32447 11135
rect 32688 11101 32722 11135
rect 32873 11101 32907 11135
rect 33333 11101 33367 11135
rect 34253 11101 34287 11135
rect 34529 11101 34563 11135
rect 34713 11101 34747 11135
rect 34989 11101 35023 11135
rect 18455 11033 18489 11067
rect 19625 11033 19659 11067
rect 20085 11033 20119 11067
rect 21465 11033 21499 11067
rect 29193 11033 29227 11067
rect 31585 11033 31619 11067
rect 34805 11033 34839 11067
rect 35173 11033 35207 11067
rect 35541 11033 35575 11067
rect 19420 10965 19454 10999
rect 25513 10965 25547 10999
rect 25973 10965 26007 10999
rect 34437 10965 34471 10999
rect 37013 10965 37047 10999
rect 18061 10761 18095 10795
rect 21833 10761 21867 10795
rect 28365 10761 28399 10795
rect 32965 10761 32999 10795
rect 35005 10761 35039 10795
rect 35173 10761 35207 10795
rect 36001 10761 36035 10795
rect 36829 10761 36863 10795
rect 16865 10693 16899 10727
rect 18337 10693 18371 10727
rect 18429 10693 18463 10727
rect 18567 10693 18601 10727
rect 19165 10693 19199 10727
rect 22477 10693 22511 10727
rect 27077 10693 27111 10727
rect 31493 10693 31527 10727
rect 33425 10693 33459 10727
rect 34805 10693 34839 10727
rect 16505 10625 16539 10659
rect 17049 10625 17083 10659
rect 17325 10625 17359 10659
rect 18246 10647 18280 10681
rect 18797 10625 18831 10659
rect 19257 10625 19291 10659
rect 19717 10625 19751 10659
rect 22017 10625 22051 10659
rect 22753 10625 22787 10659
rect 25789 10625 25823 10659
rect 25881 10625 25915 10659
rect 26157 10625 26191 10659
rect 26617 10625 26651 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 27997 10625 28031 10659
rect 28089 10625 28123 10659
rect 28457 10625 28491 10659
rect 29469 10625 29503 10659
rect 36737 10625 36771 10659
rect 17969 10557 18003 10591
rect 18705 10557 18739 10591
rect 19809 10557 19843 10591
rect 22109 10557 22143 10591
rect 23029 10557 23063 10591
rect 25513 10557 25547 10591
rect 26801 10557 26835 10591
rect 29745 10557 29779 10591
rect 36553 10557 36587 10591
rect 33057 10489 33091 10523
rect 16405 10421 16439 10455
rect 17233 10421 17267 10455
rect 18981 10421 19015 10455
rect 20085 10421 20119 10455
rect 22385 10421 22419 10455
rect 24501 10421 24535 10455
rect 24869 10421 24903 10455
rect 25605 10421 25639 10455
rect 26065 10421 26099 10455
rect 26433 10421 26467 10455
rect 27813 10421 27847 10455
rect 34989 10421 35023 10455
rect 20269 10217 20303 10251
rect 20729 10217 20763 10251
rect 23673 10217 23707 10251
rect 24501 10217 24535 10251
rect 25237 10217 25271 10251
rect 26525 10217 26559 10251
rect 30481 10217 30515 10251
rect 18245 10149 18279 10183
rect 25513 10149 25547 10183
rect 14933 10081 14967 10115
rect 20453 10081 20487 10115
rect 25145 10081 25179 10115
rect 31401 10081 31435 10115
rect 31585 10081 31619 10115
rect 32689 10081 32723 10115
rect 33793 10081 33827 10115
rect 33885 10081 33919 10115
rect 35265 10081 35299 10115
rect 14657 10013 14691 10047
rect 16865 10013 16899 10047
rect 17601 10013 17635 10047
rect 18429 10013 18463 10047
rect 18797 10013 18831 10047
rect 18889 10013 18923 10047
rect 19073 10013 19107 10047
rect 19349 10013 19383 10047
rect 19441 10013 19475 10047
rect 19533 10013 19567 10047
rect 20269 10013 20303 10047
rect 20545 10013 20579 10047
rect 23581 10013 23615 10047
rect 24685 10013 24719 10047
rect 25421 10013 25455 10047
rect 25605 10013 25639 10047
rect 25697 10013 25731 10047
rect 25881 10013 25915 10047
rect 26157 10013 26191 10047
rect 26709 10013 26743 10047
rect 29745 10013 29779 10047
rect 30389 10013 30423 10047
rect 31309 10013 31343 10047
rect 32321 10013 32355 10047
rect 32597 10013 32631 10047
rect 32873 10013 32907 10047
rect 33149 10013 33183 10047
rect 33609 10013 33643 10047
rect 33701 10013 33735 10047
rect 35449 10013 35483 10047
rect 68477 10013 68511 10047
rect 18153 9945 18187 9979
rect 18521 9945 18555 9979
rect 18613 9945 18647 9979
rect 18981 9945 19015 9979
rect 19717 9945 19751 9979
rect 24777 9945 24811 9979
rect 24869 9945 24903 9979
rect 24987 9945 25021 9979
rect 25973 9945 26007 9979
rect 32505 9945 32539 9979
rect 33057 9945 33091 9979
rect 16405 9877 16439 9911
rect 17417 9877 17451 9911
rect 26341 9877 26375 9911
rect 29653 9877 29687 9911
rect 30941 9877 30975 9911
rect 32597 9877 32631 9911
rect 33425 9877 33459 9911
rect 34713 9877 34747 9911
rect 35541 9877 35575 9911
rect 23029 9673 23063 9707
rect 24225 9673 24259 9707
rect 25513 9673 25547 9707
rect 26157 9673 26191 9707
rect 35725 9673 35759 9707
rect 18153 9605 18187 9639
rect 18857 9605 18891 9639
rect 19073 9605 19107 9639
rect 20361 9605 20395 9639
rect 21281 9605 21315 9639
rect 21925 9605 21959 9639
rect 24133 9605 24167 9639
rect 26801 9605 26835 9639
rect 31953 9605 31987 9639
rect 32505 9605 32539 9639
rect 32715 9605 32749 9639
rect 33622 9605 33656 9639
rect 34253 9605 34287 9639
rect 35909 9605 35943 9639
rect 16865 9537 16899 9571
rect 16957 9537 16991 9571
rect 17049 9537 17083 9571
rect 17167 9537 17201 9571
rect 17325 9537 17359 9571
rect 17601 9537 17635 9571
rect 17785 9537 17819 9571
rect 17877 9537 17911 9571
rect 18337 9537 18371 9571
rect 20545 9537 20579 9571
rect 21189 9537 21223 9571
rect 21373 9537 21407 9571
rect 21557 9537 21591 9571
rect 22661 9537 22695 9571
rect 22845 9537 22879 9571
rect 23305 9537 23339 9571
rect 24777 9537 24811 9571
rect 24961 9537 24995 9571
rect 26341 9537 26375 9571
rect 29377 9537 29411 9571
rect 29561 9537 29595 9571
rect 32413 9537 32447 9571
rect 32597 9537 32631 9571
rect 32873 9537 32907 9571
rect 33426 9543 33460 9577
rect 33518 9537 33552 9571
rect 33727 9537 33761 9571
rect 33977 9537 34011 9571
rect 36001 9537 36035 9571
rect 14657 9469 14691 9503
rect 14933 9469 14967 9503
rect 16681 9469 16715 9503
rect 17693 9469 17727 9503
rect 18619 9469 18653 9503
rect 22477 9469 22511 9503
rect 24409 9469 24443 9503
rect 25237 9469 25271 9503
rect 26433 9469 26467 9503
rect 27537 9469 27571 9503
rect 27813 9469 27847 9503
rect 29929 9469 29963 9503
rect 30205 9469 30239 9503
rect 33885 9469 33919 9503
rect 16405 9401 16439 9435
rect 17417 9401 17451 9435
rect 18521 9401 18555 9435
rect 18705 9401 18739 9435
rect 23765 9401 23799 9435
rect 25145 9401 25179 9435
rect 29285 9401 29319 9435
rect 18889 9333 18923 9367
rect 20729 9333 20763 9367
rect 21005 9333 21039 9367
rect 23121 9333 23155 9367
rect 25053 9333 25087 9367
rect 26341 9333 26375 9367
rect 29745 9333 29779 9367
rect 32229 9333 32263 9367
rect 33241 9333 33275 9367
rect 15945 9129 15979 9163
rect 17785 9129 17819 9163
rect 20269 9129 20303 9163
rect 20808 9129 20842 9163
rect 24133 9129 24167 9163
rect 24869 9129 24903 9163
rect 25513 9129 25547 9163
rect 26433 9129 26467 9163
rect 26985 9129 27019 9163
rect 27537 9129 27571 9163
rect 27813 9129 27847 9163
rect 31125 9129 31159 9163
rect 33977 9129 34011 9163
rect 17417 9061 17451 9095
rect 19993 9061 20027 9095
rect 22293 9061 22327 9095
rect 33425 9061 33459 9095
rect 17049 8993 17083 9027
rect 18705 8993 18739 9027
rect 20545 8993 20579 9027
rect 22385 8993 22419 9027
rect 22661 8993 22695 9027
rect 25329 8993 25363 9027
rect 30113 8993 30147 9027
rect 31309 8993 31343 9027
rect 31585 8993 31619 9027
rect 33333 8993 33367 9027
rect 16037 8925 16071 8959
rect 17233 8925 17267 8959
rect 17877 8925 17911 8959
rect 18889 8925 18923 8959
rect 19809 8925 19843 8959
rect 19993 8925 20027 8959
rect 25237 8925 25271 8959
rect 25697 8925 25731 8959
rect 25789 8925 25823 8959
rect 25881 8925 25915 8959
rect 26617 8925 26651 8959
rect 26709 8925 26743 8959
rect 27077 8925 27111 8959
rect 28457 8925 28491 8959
rect 28549 8925 28583 8959
rect 28733 8925 28767 8959
rect 29193 8925 29227 8959
rect 29561 8925 29595 8959
rect 30849 8925 30883 8959
rect 31217 8925 31251 8959
rect 33609 8925 33643 8959
rect 33701 8925 33735 8959
rect 19073 8857 19107 8891
rect 20237 8857 20271 8891
rect 20453 8857 20487 8891
rect 27353 8857 27387 8891
rect 27569 8857 27603 8891
rect 28826 8857 28860 8891
rect 28917 8857 28951 8891
rect 29055 8857 29089 8891
rect 33793 8857 33827 8891
rect 20085 8789 20119 8823
rect 27721 8789 27755 8823
rect 30297 8789 30331 8823
rect 17049 8585 17083 8619
rect 18705 8585 18739 8619
rect 19333 8585 19367 8619
rect 19717 8585 19751 8619
rect 21005 8585 21039 8619
rect 22661 8585 22695 8619
rect 23489 8585 23523 8619
rect 27077 8585 27111 8619
rect 30665 8585 30699 8619
rect 30757 8585 30791 8619
rect 31585 8585 31619 8619
rect 17141 8517 17175 8551
rect 19533 8517 19567 8551
rect 20453 8517 20487 8551
rect 20545 8517 20579 8551
rect 20683 8517 20717 8551
rect 28089 8517 28123 8551
rect 18337 8449 18371 8483
rect 18497 8449 18531 8483
rect 18629 8439 18663 8473
rect 18889 8449 18923 8483
rect 19809 8449 19843 8483
rect 20361 8449 20395 8483
rect 20913 8449 20947 8483
rect 21097 8449 21131 8483
rect 22385 8449 22419 8483
rect 22753 8449 22787 8483
rect 23397 8449 23431 8483
rect 24869 8449 24903 8483
rect 26157 8449 26191 8483
rect 27353 8449 27387 8483
rect 27445 8449 27479 8483
rect 27997 8449 28031 8483
rect 28181 8449 28215 8483
rect 28273 8449 28307 8483
rect 28457 8449 28491 8483
rect 28549 8449 28583 8483
rect 28641 8449 28675 8483
rect 28917 8449 28951 8483
rect 30941 8449 30975 8483
rect 31493 8449 31527 8483
rect 17325 8381 17359 8415
rect 20821 8381 20855 8415
rect 21833 8381 21867 8415
rect 24685 8381 24719 8415
rect 24777 8381 24811 8415
rect 24961 8381 24995 8415
rect 25789 8381 25823 8415
rect 26341 8381 26375 8415
rect 29193 8381 29227 8415
rect 18521 8313 18555 8347
rect 28825 8313 28859 8347
rect 16681 8245 16715 8279
rect 19073 8245 19107 8279
rect 19165 8245 19199 8279
rect 19349 8245 19383 8279
rect 20177 8245 20211 8279
rect 25145 8245 25179 8279
rect 25237 8245 25271 8279
rect 25973 8245 26007 8279
rect 27353 8245 27387 8279
rect 17325 8041 17359 8075
rect 29193 8041 29227 8075
rect 30205 8041 30239 8075
rect 15577 7905 15611 7939
rect 19717 7905 19751 7939
rect 19901 7905 19935 7939
rect 25053 7905 25087 7939
rect 25789 7905 25823 7939
rect 18061 7837 18095 7871
rect 18337 7837 18371 7871
rect 18981 7837 19015 7871
rect 19625 7837 19659 7871
rect 21281 7837 21315 7871
rect 22753 7837 22787 7871
rect 24409 7837 24443 7871
rect 25329 7837 25363 7871
rect 25513 7837 25547 7871
rect 26065 7837 26099 7871
rect 27077 7837 27111 7871
rect 27261 7837 27295 7871
rect 29009 7837 29043 7871
rect 29193 7837 29227 7871
rect 30297 7837 30331 7871
rect 15853 7769 15887 7803
rect 25421 7769 25455 7803
rect 25651 7769 25685 7803
rect 17877 7701 17911 7735
rect 18245 7701 18279 7735
rect 18429 7701 18463 7735
rect 19257 7701 19291 7735
rect 21189 7701 21223 7735
rect 22845 7701 22879 7735
rect 25145 7701 25179 7735
rect 25973 7701 26007 7735
rect 27169 7701 27203 7735
rect 16037 7497 16071 7531
rect 16773 7497 16807 7531
rect 19073 7497 19107 7531
rect 25513 7497 25547 7531
rect 26801 7497 26835 7531
rect 17601 7429 17635 7463
rect 20177 7429 20211 7463
rect 24225 7429 24259 7463
rect 24685 7429 24719 7463
rect 24777 7429 24811 7463
rect 25145 7429 25179 7463
rect 25361 7429 25395 7463
rect 25973 7429 26007 7463
rect 28181 7429 28215 7463
rect 16221 7361 16255 7395
rect 16865 7361 16899 7395
rect 19349 7361 19383 7395
rect 19901 7361 19935 7395
rect 21925 7361 21959 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 24593 7361 24627 7395
rect 24915 7361 24949 7395
rect 25053 7361 25087 7395
rect 25789 7361 25823 7395
rect 26617 7361 26651 7395
rect 27353 7361 27387 7395
rect 27997 7361 28031 7395
rect 17325 7293 17359 7327
rect 22201 7293 22235 7327
rect 25605 7293 25639 7327
rect 26433 7293 26467 7327
rect 27077 7293 27111 7327
rect 27261 7293 27295 7327
rect 27813 7293 27847 7327
rect 21649 7225 21683 7259
rect 23673 7225 23707 7259
rect 19533 7157 19567 7191
rect 24409 7157 24443 7191
rect 25329 7157 25363 7191
rect 27721 7157 27755 7191
rect 18429 6953 18463 6987
rect 20066 6953 20100 6987
rect 22464 6953 22498 6987
rect 27353 6953 27387 6987
rect 21557 6817 21591 6851
rect 22201 6817 22235 6851
rect 24225 6817 24259 6851
rect 26525 6817 26559 6851
rect 26801 6817 26835 6851
rect 27445 6817 27479 6851
rect 29193 6817 29227 6851
rect 18337 6749 18371 6783
rect 19809 6749 19843 6783
rect 21833 6749 21867 6783
rect 26985 6749 27019 6783
rect 27169 6749 27203 6783
rect 29745 6749 29779 6783
rect 21741 6681 21775 6715
rect 27721 6681 27755 6715
rect 29653 6681 29687 6715
rect 25053 6613 25087 6647
rect 23581 6409 23615 6443
rect 26157 6409 26191 6443
rect 28365 6409 28399 6443
rect 27905 6341 27939 6375
rect 27997 6341 28031 6375
rect 23673 6273 23707 6307
rect 26065 6273 26099 6307
rect 26985 6273 27019 6307
rect 27629 6273 27663 6307
rect 27721 6273 27755 6307
rect 28089 6273 28123 6307
rect 28549 6273 28583 6307
rect 28273 6137 28307 6171
rect 43085 3009 43119 3043
rect 43269 2805 43303 2839
rect 26525 2397 26559 2431
rect 44005 2397 44039 2431
rect 67649 2397 67683 2431
rect 44281 2261 44315 2295
rect 67925 2261 67959 2295
<< metal1 >>
rect 1104 67482 68816 67504
rect 1104 67430 19574 67482
rect 19626 67430 19638 67482
rect 19690 67430 19702 67482
rect 19754 67430 19766 67482
rect 19818 67430 19830 67482
rect 19882 67430 50294 67482
rect 50346 67430 50358 67482
rect 50410 67430 50422 67482
rect 50474 67430 50486 67482
rect 50538 67430 50550 67482
rect 50602 67430 68816 67482
rect 1104 67408 68816 67430
rect 12986 67192 12992 67244
rect 13044 67192 13050 67244
rect 30374 67192 30380 67244
rect 30432 67192 30438 67244
rect 39390 67192 39396 67244
rect 39448 67192 39454 67244
rect 1104 66938 68816 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 68816 66938
rect 1104 66864 68816 66886
rect 1104 66394 68816 66416
rect 1104 66342 19574 66394
rect 19626 66342 19638 66394
rect 19690 66342 19702 66394
rect 19754 66342 19766 66394
rect 19818 66342 19830 66394
rect 19882 66342 50294 66394
rect 50346 66342 50358 66394
rect 50410 66342 50422 66394
rect 50474 66342 50486 66394
rect 50538 66342 50550 66394
rect 50602 66342 68816 66394
rect 1104 66320 68816 66342
rect 1104 65850 68816 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 68816 65850
rect 1104 65776 68816 65798
rect 1104 65306 68816 65328
rect 1104 65254 19574 65306
rect 19626 65254 19638 65306
rect 19690 65254 19702 65306
rect 19754 65254 19766 65306
rect 19818 65254 19830 65306
rect 19882 65254 50294 65306
rect 50346 65254 50358 65306
rect 50410 65254 50422 65306
rect 50474 65254 50486 65306
rect 50538 65254 50550 65306
rect 50602 65254 68816 65306
rect 1104 65232 68816 65254
rect 1394 64948 1400 65000
rect 1452 64948 1458 65000
rect 1104 64762 68816 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 34934 64762
rect 34986 64710 34998 64762
rect 35050 64710 35062 64762
rect 35114 64710 35126 64762
rect 35178 64710 35190 64762
rect 35242 64710 65654 64762
rect 65706 64710 65718 64762
rect 65770 64710 65782 64762
rect 65834 64710 65846 64762
rect 65898 64710 65910 64762
rect 65962 64710 68816 64762
rect 1104 64688 68816 64710
rect 1104 64218 68816 64240
rect 1104 64166 19574 64218
rect 19626 64166 19638 64218
rect 19690 64166 19702 64218
rect 19754 64166 19766 64218
rect 19818 64166 19830 64218
rect 19882 64166 50294 64218
rect 50346 64166 50358 64218
rect 50410 64166 50422 64218
rect 50474 64166 50486 64218
rect 50538 64166 50550 64218
rect 50602 64166 68816 64218
rect 1104 64144 68816 64166
rect 1104 63674 68816 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 34934 63674
rect 34986 63622 34998 63674
rect 35050 63622 35062 63674
rect 35114 63622 35126 63674
rect 35178 63622 35190 63674
rect 35242 63622 65654 63674
rect 65706 63622 65718 63674
rect 65770 63622 65782 63674
rect 65834 63622 65846 63674
rect 65898 63622 65910 63674
rect 65962 63622 68816 63674
rect 1104 63600 68816 63622
rect 1104 63130 68816 63152
rect 1104 63078 19574 63130
rect 19626 63078 19638 63130
rect 19690 63078 19702 63130
rect 19754 63078 19766 63130
rect 19818 63078 19830 63130
rect 19882 63078 50294 63130
rect 50346 63078 50358 63130
rect 50410 63078 50422 63130
rect 50474 63078 50486 63130
rect 50538 63078 50550 63130
rect 50602 63078 68816 63130
rect 1104 63056 68816 63078
rect 1104 62586 68816 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 34934 62586
rect 34986 62534 34998 62586
rect 35050 62534 35062 62586
rect 35114 62534 35126 62586
rect 35178 62534 35190 62586
rect 35242 62534 65654 62586
rect 65706 62534 65718 62586
rect 65770 62534 65782 62586
rect 65834 62534 65846 62586
rect 65898 62534 65910 62586
rect 65962 62534 68816 62586
rect 1104 62512 68816 62534
rect 1104 62042 68816 62064
rect 1104 61990 19574 62042
rect 19626 61990 19638 62042
rect 19690 61990 19702 62042
rect 19754 61990 19766 62042
rect 19818 61990 19830 62042
rect 19882 61990 50294 62042
rect 50346 61990 50358 62042
rect 50410 61990 50422 62042
rect 50474 61990 50486 62042
rect 50538 61990 50550 62042
rect 50602 61990 68816 62042
rect 1104 61968 68816 61990
rect 1104 61498 68816 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 65654 61498
rect 65706 61446 65718 61498
rect 65770 61446 65782 61498
rect 65834 61446 65846 61498
rect 65898 61446 65910 61498
rect 65962 61446 68816 61498
rect 1104 61424 68816 61446
rect 1104 60954 68816 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 68816 60954
rect 1104 60880 68816 60902
rect 1104 60410 68816 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 65654 60410
rect 65706 60358 65718 60410
rect 65770 60358 65782 60410
rect 65834 60358 65846 60410
rect 65898 60358 65910 60410
rect 65962 60358 68816 60410
rect 1104 60336 68816 60358
rect 1104 59866 68816 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 68816 59866
rect 1104 59792 68816 59814
rect 1104 59322 68816 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 65654 59322
rect 65706 59270 65718 59322
rect 65770 59270 65782 59322
rect 65834 59270 65846 59322
rect 65898 59270 65910 59322
rect 65962 59270 68816 59322
rect 1104 59248 68816 59270
rect 1104 58778 68816 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 68816 58778
rect 1104 58704 68816 58726
rect 1104 58234 68816 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 65654 58234
rect 65706 58182 65718 58234
rect 65770 58182 65782 58234
rect 65834 58182 65846 58234
rect 65898 58182 65910 58234
rect 65962 58182 68816 58234
rect 1104 58160 68816 58182
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 68462 56108 68468 56160
rect 68520 56108 68526 56160
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 1762 46520 1768 46572
rect 1820 46520 1826 46572
rect 934 46316 940 46368
rect 992 46356 998 46368
rect 1489 46359 1547 46365
rect 1489 46356 1501 46359
rect 992 46328 1501 46356
rect 992 46316 998 46328
rect 1489 46325 1501 46328
rect 1535 46325 1547 46359
rect 1489 46319 1547 46325
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 1765 37315 1823 37321
rect 1765 37281 1777 37315
rect 1811 37312 1823 37315
rect 18230 37312 18236 37324
rect 1811 37284 18236 37312
rect 1811 37281 1823 37284
rect 1765 37275 1823 37281
rect 18230 37272 18236 37284
rect 18288 37272 18294 37324
rect 934 37136 940 37188
rect 992 37176 998 37188
rect 1489 37179 1547 37185
rect 1489 37176 1501 37179
rect 992 37148 1501 37176
rect 992 37136 998 37148
rect 1489 37145 1501 37148
rect 1535 37145 1547 37179
rect 1489 37139 1547 37145
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 20993 29155 21051 29161
rect 20993 29121 21005 29155
rect 21039 29152 21051 29155
rect 21726 29152 21732 29164
rect 21039 29124 21732 29152
rect 21039 29121 21051 29124
rect 20993 29115 21051 29121
rect 21726 29112 21732 29124
rect 21784 29152 21790 29164
rect 22649 29155 22707 29161
rect 22649 29152 22661 29155
rect 21784 29124 22661 29152
rect 21784 29112 21790 29124
rect 22649 29121 22661 29124
rect 22695 29152 22707 29155
rect 24029 29155 24087 29161
rect 24029 29152 24041 29155
rect 22695 29124 24041 29152
rect 22695 29121 22707 29124
rect 22649 29115 22707 29121
rect 24029 29121 24041 29124
rect 24075 29152 24087 29155
rect 24765 29155 24823 29161
rect 24765 29152 24777 29155
rect 24075 29124 24777 29152
rect 24075 29121 24087 29124
rect 24029 29115 24087 29121
rect 24765 29121 24777 29124
rect 24811 29121 24823 29155
rect 24765 29115 24823 29121
rect 23934 29044 23940 29096
rect 23992 29044 23998 29096
rect 22741 29019 22799 29025
rect 22741 28985 22753 29019
rect 22787 29016 22799 29019
rect 24121 29019 24179 29025
rect 22787 28988 23520 29016
rect 22787 28985 22799 28988
rect 22741 28979 22799 28985
rect 23492 28960 23520 28988
rect 24121 28985 24133 29019
rect 24167 29016 24179 29019
rect 24167 28988 25176 29016
rect 24167 28985 24179 28988
rect 24121 28979 24179 28985
rect 25148 28960 25176 28988
rect 21082 28908 21088 28960
rect 21140 28908 21146 28960
rect 23290 28908 23296 28960
rect 23348 28908 23354 28960
rect 23474 28908 23480 28960
rect 23532 28908 23538 28960
rect 24854 28908 24860 28960
rect 24912 28908 24918 28960
rect 25130 28908 25136 28960
rect 25188 28908 25194 28960
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 24397 28611 24455 28617
rect 24397 28577 24409 28611
rect 24443 28608 24455 28611
rect 25406 28608 25412 28620
rect 24443 28580 25412 28608
rect 24443 28577 24455 28580
rect 24397 28571 24455 28577
rect 25406 28568 25412 28580
rect 25464 28568 25470 28620
rect 20073 28543 20131 28549
rect 20073 28509 20085 28543
rect 20119 28509 20131 28543
rect 20073 28503 20131 28509
rect 22189 28543 22247 28549
rect 22189 28509 22201 28543
rect 22235 28509 22247 28543
rect 22189 28503 22247 28509
rect 17954 28364 17960 28416
rect 18012 28404 18018 28416
rect 20088 28404 20116 28503
rect 20346 28432 20352 28484
rect 20404 28432 20410 28484
rect 21082 28432 21088 28484
rect 21140 28432 21146 28484
rect 22094 28432 22100 28484
rect 22152 28432 22158 28484
rect 22204 28404 22232 28503
rect 22462 28432 22468 28484
rect 22520 28432 22526 28484
rect 23474 28432 23480 28484
rect 23532 28432 23538 28484
rect 24670 28432 24676 28484
rect 24728 28432 24734 28484
rect 25130 28432 25136 28484
rect 25188 28432 25194 28484
rect 25958 28432 25964 28484
rect 26016 28472 26022 28484
rect 26421 28475 26479 28481
rect 26421 28472 26433 28475
rect 26016 28444 26433 28472
rect 26016 28432 26022 28444
rect 26421 28441 26433 28444
rect 26467 28441 26479 28475
rect 26421 28435 26479 28441
rect 18012 28376 22232 28404
rect 18012 28364 18018 28376
rect 23934 28364 23940 28416
rect 23992 28364 23998 28416
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 20346 28160 20352 28212
rect 20404 28200 20410 28212
rect 20441 28203 20499 28209
rect 20441 28200 20453 28203
rect 20404 28172 20453 28200
rect 20404 28160 20410 28172
rect 20441 28169 20453 28172
rect 20487 28169 20499 28203
rect 20441 28163 20499 28169
rect 20717 28203 20775 28209
rect 20717 28169 20729 28203
rect 20763 28169 20775 28203
rect 20717 28163 20775 28169
rect 22189 28203 22247 28209
rect 22189 28169 22201 28203
rect 22235 28200 22247 28203
rect 22462 28200 22468 28212
rect 22235 28172 22468 28200
rect 22235 28169 22247 28172
rect 22189 28163 22247 28169
rect 20625 28067 20683 28073
rect 20625 28033 20637 28067
rect 20671 28064 20683 28067
rect 20732 28064 20760 28163
rect 22462 28160 22468 28172
rect 22520 28160 22526 28212
rect 21085 28135 21143 28141
rect 21085 28101 21097 28135
rect 21131 28132 21143 28135
rect 22675 28135 22733 28141
rect 21131 28104 22600 28132
rect 21131 28101 21143 28104
rect 21085 28095 21143 28101
rect 22572 28076 22600 28104
rect 22675 28101 22687 28135
rect 22721 28101 22733 28135
rect 22675 28095 22733 28101
rect 20671 28036 20760 28064
rect 20671 28033 20683 28036
rect 20625 28027 20683 28033
rect 21174 28024 21180 28076
rect 21232 28064 21238 28076
rect 21232 28036 22324 28064
rect 21232 28024 21238 28036
rect 21361 27999 21419 28005
rect 21361 27965 21373 27999
rect 21407 27996 21419 27999
rect 22094 27996 22100 28008
rect 21407 27968 22100 27996
rect 21407 27965 21419 27968
rect 21361 27959 21419 27965
rect 22094 27956 22100 27968
rect 22152 27956 22158 28008
rect 22296 27996 22324 28036
rect 22370 28024 22376 28076
rect 22428 28024 22434 28076
rect 22462 28024 22468 28076
rect 22520 28024 22526 28076
rect 22554 28024 22560 28076
rect 22612 28024 22618 28076
rect 22690 28064 22718 28095
rect 24854 28092 24860 28144
rect 24912 28092 24918 28144
rect 25406 28092 25412 28144
rect 25464 28132 25470 28144
rect 25464 28104 25728 28132
rect 25464 28092 25470 28104
rect 22664 28036 22718 28064
rect 22833 28067 22891 28073
rect 22664 28008 22692 28036
rect 22833 28033 22845 28067
rect 22879 28064 22891 28067
rect 23290 28064 23296 28076
rect 22879 28036 23296 28064
rect 22879 28033 22891 28036
rect 22833 28027 22891 28033
rect 23290 28024 23296 28036
rect 23348 28024 23354 28076
rect 25700 28073 25728 28104
rect 25685 28067 25743 28073
rect 25685 28033 25697 28067
rect 25731 28033 25743 28067
rect 25685 28027 25743 28033
rect 68373 28067 68431 28073
rect 68373 28033 68385 28067
rect 68419 28064 68431 28067
rect 68830 28064 68836 28076
rect 68419 28036 68836 28064
rect 68419 28033 68431 28036
rect 68373 28027 68431 28033
rect 68830 28024 68836 28036
rect 68888 28024 68894 28076
rect 22646 27996 22652 28008
rect 22296 27968 22652 27996
rect 22646 27956 22652 27968
rect 22704 27956 22710 28008
rect 23201 27999 23259 28005
rect 23201 27965 23213 27999
rect 23247 27996 23259 27999
rect 23247 27968 23612 27996
rect 23247 27965 23259 27968
rect 23201 27959 23259 27965
rect 23584 27928 23612 27968
rect 25038 27956 25044 28008
rect 25096 27996 25102 28008
rect 25409 27999 25467 28005
rect 25409 27996 25421 27999
rect 25096 27968 25421 27996
rect 25096 27956 25102 27968
rect 25409 27965 25421 27968
rect 25455 27965 25467 27999
rect 25409 27959 25467 27965
rect 23937 27931 23995 27937
rect 23937 27928 23949 27931
rect 23584 27900 23949 27928
rect 23584 27872 23612 27900
rect 23937 27897 23949 27900
rect 23983 27897 23995 27931
rect 23937 27891 23995 27897
rect 23566 27820 23572 27872
rect 23624 27820 23630 27872
rect 23750 27820 23756 27872
rect 23808 27820 23814 27872
rect 68278 27820 68284 27872
rect 68336 27820 68342 27872
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 22370 27616 22376 27668
rect 22428 27656 22434 27668
rect 22925 27659 22983 27665
rect 22925 27656 22937 27659
rect 22428 27628 22937 27656
rect 22428 27616 22434 27628
rect 22925 27625 22937 27628
rect 22971 27625 22983 27659
rect 22925 27619 22983 27625
rect 25038 27616 25044 27668
rect 25096 27616 25102 27668
rect 22646 27548 22652 27600
rect 22704 27588 22710 27600
rect 24210 27588 24216 27600
rect 22704 27560 24216 27588
rect 22704 27548 22710 27560
rect 24210 27548 24216 27560
rect 24268 27588 24274 27600
rect 24268 27560 24532 27588
rect 24268 27548 24274 27560
rect 22094 27480 22100 27532
rect 22152 27520 22158 27532
rect 22922 27520 22928 27532
rect 22152 27492 22928 27520
rect 22152 27480 22158 27492
rect 22922 27480 22928 27492
rect 22980 27520 22986 27532
rect 23109 27523 23167 27529
rect 23109 27520 23121 27523
rect 22980 27492 23121 27520
rect 22980 27480 22986 27492
rect 23109 27489 23121 27492
rect 23155 27489 23167 27523
rect 23109 27483 23167 27489
rect 23293 27523 23351 27529
rect 23293 27489 23305 27523
rect 23339 27520 23351 27523
rect 23339 27492 23612 27520
rect 23339 27489 23351 27492
rect 23293 27483 23351 27489
rect 23584 27464 23612 27492
rect 23750 27480 23756 27532
rect 23808 27520 23814 27532
rect 24397 27523 24455 27529
rect 24397 27520 24409 27523
rect 23808 27492 24409 27520
rect 23808 27480 23814 27492
rect 24397 27489 24409 27492
rect 24443 27489 24455 27523
rect 24504 27520 24532 27560
rect 25406 27548 25412 27600
rect 25464 27588 25470 27600
rect 25464 27560 26188 27588
rect 25464 27548 25470 27560
rect 26160 27529 26188 27560
rect 25225 27523 25283 27529
rect 25225 27520 25237 27523
rect 24504 27492 24578 27520
rect 24397 27483 24455 27489
rect 20809 27455 20867 27461
rect 20809 27452 20821 27455
rect 20640 27424 20821 27452
rect 20640 27328 20668 27424
rect 20809 27421 20821 27424
rect 20855 27421 20867 27455
rect 20809 27415 20867 27421
rect 20990 27412 20996 27464
rect 21048 27412 21054 27464
rect 23201 27455 23259 27461
rect 23201 27421 23213 27455
rect 23247 27452 23259 27455
rect 23247 27424 23336 27452
rect 23247 27421 23259 27424
rect 23201 27415 23259 27421
rect 23308 27396 23336 27424
rect 23382 27412 23388 27464
rect 23440 27412 23446 27464
rect 23566 27412 23572 27464
rect 23624 27412 23630 27464
rect 24550 27461 24578 27492
rect 24872 27492 25237 27520
rect 24872 27461 24900 27492
rect 25225 27489 25237 27492
rect 25271 27489 25283 27523
rect 25225 27483 25283 27489
rect 26145 27523 26203 27529
rect 26145 27489 26157 27523
rect 26191 27489 26203 27523
rect 26145 27483 26203 27489
rect 24535 27455 24593 27461
rect 24535 27421 24547 27455
rect 24581 27421 24593 27455
rect 24535 27415 24593 27421
rect 24857 27455 24915 27461
rect 24857 27421 24869 27455
rect 24903 27421 24915 27455
rect 24857 27415 24915 27421
rect 25133 27455 25191 27461
rect 25133 27421 25145 27455
rect 25179 27421 25191 27455
rect 25133 27415 25191 27421
rect 23290 27344 23296 27396
rect 23348 27344 23354 27396
rect 23400 27384 23428 27412
rect 23934 27384 23940 27396
rect 23400 27356 23940 27384
rect 23934 27344 23940 27356
rect 23992 27344 23998 27396
rect 24673 27387 24731 27393
rect 24673 27353 24685 27387
rect 24719 27353 24731 27387
rect 24673 27347 24731 27353
rect 20622 27276 20628 27328
rect 20680 27276 20686 27328
rect 20901 27319 20959 27325
rect 20901 27285 20913 27319
rect 20947 27316 20959 27319
rect 21266 27316 21272 27328
rect 20947 27288 21272 27316
rect 20947 27285 20959 27288
rect 20901 27279 20959 27285
rect 21266 27276 21272 27288
rect 21324 27276 21330 27328
rect 21634 27276 21640 27328
rect 21692 27316 21698 27328
rect 22554 27316 22560 27328
rect 21692 27288 22560 27316
rect 21692 27276 21698 27288
rect 22554 27276 22560 27288
rect 22612 27316 22618 27328
rect 23014 27316 23020 27328
rect 22612 27288 23020 27316
rect 22612 27276 22618 27288
rect 23014 27276 23020 27288
rect 23072 27316 23078 27328
rect 24688 27316 24716 27347
rect 24762 27344 24768 27396
rect 24820 27344 24826 27396
rect 25038 27344 25044 27396
rect 25096 27384 25102 27396
rect 25148 27384 25176 27415
rect 25314 27412 25320 27464
rect 25372 27412 25378 27464
rect 25406 27412 25412 27464
rect 25464 27412 25470 27464
rect 26050 27412 26056 27464
rect 26108 27452 26114 27464
rect 26160 27452 26188 27483
rect 27985 27455 28043 27461
rect 27985 27452 27997 27455
rect 26108 27424 27997 27452
rect 26108 27412 26114 27424
rect 27985 27421 27997 27424
rect 28031 27421 28043 27455
rect 30101 27455 30159 27461
rect 30101 27452 30113 27455
rect 27985 27415 28043 27421
rect 29380 27424 30113 27452
rect 26412 27387 26470 27393
rect 25096 27356 25544 27384
rect 25096 27344 25102 27356
rect 25516 27325 25544 27356
rect 26412 27353 26424 27387
rect 26458 27384 26470 27387
rect 26602 27384 26608 27396
rect 26458 27356 26608 27384
rect 26458 27353 26470 27356
rect 26412 27347 26470 27353
rect 26602 27344 26608 27356
rect 26660 27344 26666 27396
rect 28252 27387 28310 27393
rect 28252 27353 28264 27387
rect 28298 27384 28310 27387
rect 28626 27384 28632 27396
rect 28298 27356 28632 27384
rect 28298 27353 28310 27356
rect 28252 27347 28310 27353
rect 28626 27344 28632 27356
rect 28684 27344 28690 27396
rect 29380 27328 29408 27424
rect 30101 27421 30113 27424
rect 30147 27421 30159 27455
rect 30101 27415 30159 27421
rect 30469 27455 30527 27461
rect 30469 27421 30481 27455
rect 30515 27452 30527 27455
rect 30558 27452 30564 27464
rect 30515 27424 30564 27452
rect 30515 27421 30527 27424
rect 30469 27415 30527 27421
rect 30558 27412 30564 27424
rect 30616 27412 30622 27464
rect 23072 27288 24716 27316
rect 25501 27319 25559 27325
rect 23072 27276 23078 27288
rect 25501 27285 25513 27319
rect 25547 27316 25559 27319
rect 25774 27316 25780 27328
rect 25547 27288 25780 27316
rect 25547 27285 25559 27288
rect 25501 27279 25559 27285
rect 25774 27276 25780 27288
rect 25832 27276 25838 27328
rect 27525 27319 27583 27325
rect 27525 27285 27537 27319
rect 27571 27316 27583 27319
rect 27706 27316 27712 27328
rect 27571 27288 27712 27316
rect 27571 27285 27583 27288
rect 27525 27279 27583 27285
rect 27706 27276 27712 27288
rect 27764 27276 27770 27328
rect 29362 27276 29368 27328
rect 29420 27276 29426 27328
rect 29546 27276 29552 27328
rect 29604 27276 29610 27328
rect 30282 27276 30288 27328
rect 30340 27276 30346 27328
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 19613 27115 19671 27121
rect 19613 27081 19625 27115
rect 19659 27112 19671 27115
rect 20622 27112 20628 27124
rect 19659 27084 20628 27112
rect 19659 27081 19671 27084
rect 19613 27075 19671 27081
rect 20622 27072 20628 27084
rect 20680 27112 20686 27124
rect 20680 27084 20944 27112
rect 20680 27072 20686 27084
rect 18782 27004 18788 27056
rect 18840 27004 18846 27056
rect 17862 26936 17868 26988
rect 17920 26936 17926 26988
rect 20073 26979 20131 26985
rect 20073 26945 20085 26979
rect 20119 26976 20131 26979
rect 20806 26976 20812 26988
rect 20119 26948 20812 26976
rect 20119 26945 20131 26948
rect 20073 26939 20131 26945
rect 20806 26936 20812 26948
rect 20864 26936 20870 26988
rect 18141 26911 18199 26917
rect 18141 26877 18153 26911
rect 18187 26908 18199 26911
rect 19794 26908 19800 26920
rect 18187 26880 19800 26908
rect 18187 26877 18199 26880
rect 18141 26871 18199 26877
rect 19794 26868 19800 26880
rect 19852 26868 19858 26920
rect 20165 26911 20223 26917
rect 20165 26877 20177 26911
rect 20211 26877 20223 26911
rect 20165 26871 20223 26877
rect 19702 26732 19708 26784
rect 19760 26732 19766 26784
rect 20180 26772 20208 26871
rect 20346 26868 20352 26920
rect 20404 26868 20410 26920
rect 20916 26908 20944 27084
rect 20990 27072 20996 27124
rect 21048 27072 21054 27124
rect 21266 27072 21272 27124
rect 21324 27112 21330 27124
rect 21427 27115 21485 27121
rect 21427 27112 21439 27115
rect 21324 27084 21439 27112
rect 21324 27072 21330 27084
rect 21427 27081 21439 27084
rect 21473 27081 21485 27115
rect 21427 27075 21485 27081
rect 22462 27072 22468 27124
rect 22520 27112 22526 27124
rect 22649 27115 22707 27121
rect 22649 27112 22661 27115
rect 22520 27084 22661 27112
rect 22520 27072 22526 27084
rect 22649 27081 22661 27084
rect 22695 27081 22707 27115
rect 22649 27075 22707 27081
rect 22738 27072 22744 27124
rect 22796 27112 22802 27124
rect 22922 27112 22928 27124
rect 22796 27084 22928 27112
rect 22796 27072 22802 27084
rect 22922 27072 22928 27084
rect 22980 27112 22986 27124
rect 23017 27115 23075 27121
rect 23017 27112 23029 27115
rect 22980 27084 23029 27112
rect 22980 27072 22986 27084
rect 23017 27081 23029 27084
rect 23063 27081 23075 27115
rect 23017 27075 23075 27081
rect 23109 27115 23167 27121
rect 23109 27081 23121 27115
rect 23155 27112 23167 27115
rect 23290 27112 23296 27124
rect 23155 27084 23296 27112
rect 23155 27081 23167 27084
rect 23109 27075 23167 27081
rect 23290 27072 23296 27084
rect 23348 27112 23354 27124
rect 23348 27084 24072 27112
rect 23348 27072 23354 27084
rect 21008 26976 21036 27072
rect 21634 27004 21640 27056
rect 21692 27004 21698 27056
rect 22480 27044 22508 27072
rect 22296 27016 22508 27044
rect 23201 27047 23259 27053
rect 22296 26985 22324 27016
rect 23201 27013 23213 27047
rect 23247 27044 23259 27047
rect 23566 27044 23572 27056
rect 23247 27016 23572 27044
rect 23247 27013 23259 27016
rect 23201 27007 23259 27013
rect 23566 27004 23572 27016
rect 23624 27004 23630 27056
rect 22281 26979 22339 26985
rect 21008 26948 21404 26976
rect 21085 26911 21143 26917
rect 21085 26908 21097 26911
rect 20916 26880 21097 26908
rect 21085 26877 21097 26880
rect 21131 26877 21143 26911
rect 21085 26871 21143 26877
rect 20438 26800 20444 26852
rect 20496 26840 20502 26852
rect 21269 26843 21327 26849
rect 21269 26840 21281 26843
rect 20496 26812 21281 26840
rect 20496 26800 20502 26812
rect 21269 26809 21281 26812
rect 21315 26809 21327 26843
rect 21269 26803 21327 26809
rect 20254 26772 20260 26784
rect 20180 26744 20260 26772
rect 20254 26732 20260 26744
rect 20312 26732 20318 26784
rect 20530 26732 20536 26784
rect 20588 26732 20594 26784
rect 21376 26772 21404 26948
rect 22281 26945 22293 26979
rect 22327 26945 22339 26979
rect 22281 26939 22339 26945
rect 22465 26979 22523 26985
rect 22465 26945 22477 26979
rect 22511 26945 22523 26979
rect 22465 26939 22523 26945
rect 22741 26979 22799 26985
rect 22741 26945 22753 26979
rect 22787 26976 22799 26979
rect 22830 26976 22836 26988
rect 22787 26948 22836 26976
rect 22787 26945 22799 26948
rect 22741 26939 22799 26945
rect 22480 26908 22508 26939
rect 22830 26936 22836 26948
rect 22888 26936 22894 26988
rect 23474 26936 23480 26988
rect 23532 26936 23538 26988
rect 22646 26908 22652 26920
rect 22480 26880 22652 26908
rect 22646 26868 22652 26880
rect 22704 26908 22710 26920
rect 23584 26917 23612 27004
rect 23569 26911 23627 26917
rect 22704 26880 23520 26908
rect 22704 26868 22710 26880
rect 22922 26800 22928 26852
rect 22980 26840 22986 26852
rect 23382 26840 23388 26852
rect 22980 26812 23388 26840
rect 22980 26800 22986 26812
rect 23382 26800 23388 26812
rect 23440 26800 23446 26852
rect 21453 26775 21511 26781
rect 21453 26772 21465 26775
rect 21376 26744 21465 26772
rect 21453 26741 21465 26744
rect 21499 26772 21511 26775
rect 22281 26775 22339 26781
rect 22281 26772 22293 26775
rect 21499 26744 22293 26772
rect 21499 26741 21511 26744
rect 21453 26735 21511 26741
rect 22281 26741 22293 26744
rect 22327 26741 22339 26775
rect 22281 26735 22339 26741
rect 22830 26732 22836 26784
rect 22888 26732 22894 26784
rect 23492 26781 23520 26880
rect 23569 26877 23581 26911
rect 23615 26908 23627 26911
rect 23658 26908 23664 26920
rect 23615 26880 23664 26908
rect 23615 26877 23627 26880
rect 23569 26871 23627 26877
rect 23658 26868 23664 26880
rect 23716 26868 23722 26920
rect 24044 26917 24072 27084
rect 24670 27072 24676 27124
rect 24728 27072 24734 27124
rect 24762 27072 24768 27124
rect 24820 27072 24826 27124
rect 26602 27072 26608 27124
rect 26660 27112 26666 27124
rect 26697 27115 26755 27121
rect 26697 27112 26709 27115
rect 26660 27084 26709 27112
rect 26660 27072 26666 27084
rect 26697 27081 26709 27084
rect 26743 27081 26755 27115
rect 26697 27075 26755 27081
rect 28626 27072 28632 27124
rect 28684 27072 28690 27124
rect 29546 27072 29552 27124
rect 29604 27072 29610 27124
rect 30282 27072 30288 27124
rect 30340 27072 30346 27124
rect 24210 27053 24216 27056
rect 24187 27047 24216 27053
rect 24187 27013 24199 27047
rect 24187 27007 24216 27013
rect 24210 27004 24216 27007
rect 24268 27004 24274 27056
rect 24397 27047 24455 27053
rect 24397 27013 24409 27047
rect 24443 27044 24455 27047
rect 25225 27047 25283 27053
rect 25225 27044 25237 27047
rect 24443 27016 25237 27044
rect 24443 27013 24455 27016
rect 24397 27007 24455 27013
rect 25225 27013 25237 27016
rect 25271 27013 25283 27047
rect 25225 27007 25283 27013
rect 25409 27047 25467 27053
rect 25409 27013 25421 27047
rect 25455 27044 25467 27047
rect 25498 27044 25504 27056
rect 25455 27016 25504 27044
rect 25455 27013 25467 27016
rect 25409 27007 25467 27013
rect 25498 27004 25504 27016
rect 25556 27044 25562 27056
rect 25958 27044 25964 27056
rect 25556 27016 25964 27044
rect 25556 27004 25562 27016
rect 25958 27004 25964 27016
rect 26016 27004 26022 27056
rect 27065 27047 27123 27053
rect 27065 27044 27077 27047
rect 26620 27016 27077 27044
rect 24302 26936 24308 26988
rect 24360 26936 24366 26988
rect 24489 26979 24547 26985
rect 24489 26945 24501 26979
rect 24535 26945 24547 26979
rect 24489 26939 24547 26945
rect 24949 26979 25007 26985
rect 24949 26945 24961 26979
rect 24995 26976 25007 26979
rect 25038 26976 25044 26988
rect 24995 26948 25044 26976
rect 24995 26945 25007 26948
rect 24949 26939 25007 26945
rect 24029 26911 24087 26917
rect 24029 26877 24041 26911
rect 24075 26877 24087 26911
rect 24504 26908 24532 26939
rect 25038 26936 25044 26948
rect 25096 26936 25102 26988
rect 25133 26979 25191 26985
rect 25133 26945 25145 26979
rect 25179 26945 25191 26979
rect 25133 26939 25191 26945
rect 25148 26908 25176 26939
rect 25590 26936 25596 26988
rect 25648 26976 25654 26988
rect 25685 26979 25743 26985
rect 25685 26976 25697 26979
rect 25648 26948 25697 26976
rect 25648 26936 25654 26948
rect 25685 26945 25697 26948
rect 25731 26945 25743 26979
rect 25685 26939 25743 26945
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26976 25927 26979
rect 25976 26976 26004 27004
rect 26620 26985 26648 27016
rect 27065 27013 27077 27016
rect 27111 27013 27123 27047
rect 27893 27047 27951 27053
rect 27893 27044 27905 27047
rect 27065 27007 27123 27013
rect 27356 27016 27905 27044
rect 27356 26985 27384 27016
rect 27893 27013 27905 27016
rect 27939 27013 27951 27047
rect 27893 27007 27951 27013
rect 25915 26948 26004 26976
rect 26605 26979 26663 26985
rect 25915 26945 25927 26948
rect 25869 26939 25927 26945
rect 26605 26945 26617 26979
rect 26651 26945 26663 26979
rect 26605 26939 26663 26945
rect 26789 26979 26847 26985
rect 26789 26945 26801 26979
rect 26835 26945 26847 26979
rect 26789 26939 26847 26945
rect 27341 26979 27399 26985
rect 27341 26945 27353 26979
rect 27387 26945 27399 26979
rect 27341 26939 27399 26945
rect 27617 26979 27675 26985
rect 27617 26945 27629 26979
rect 27663 26945 27675 26979
rect 27617 26939 27675 26945
rect 25314 26908 25320 26920
rect 24504 26880 25320 26908
rect 24029 26871 24087 26877
rect 23477 26775 23535 26781
rect 23477 26741 23489 26775
rect 23523 26741 23535 26775
rect 23477 26735 23535 26741
rect 23842 26732 23848 26784
rect 23900 26732 23906 26784
rect 24044 26772 24072 26871
rect 25314 26868 25320 26880
rect 25372 26908 25378 26920
rect 25777 26911 25835 26917
rect 25777 26908 25789 26911
rect 25372 26880 25789 26908
rect 25372 26868 25378 26880
rect 25777 26877 25789 26880
rect 25823 26877 25835 26911
rect 25777 26871 25835 26877
rect 25498 26800 25504 26852
rect 25556 26800 25562 26852
rect 26804 26840 26832 26939
rect 27065 26911 27123 26917
rect 27065 26877 27077 26911
rect 27111 26908 27123 26911
rect 27154 26908 27160 26920
rect 27111 26880 27160 26908
rect 27111 26877 27123 26880
rect 27065 26871 27123 26877
rect 27154 26868 27160 26880
rect 27212 26868 27218 26920
rect 27249 26911 27307 26917
rect 27249 26877 27261 26911
rect 27295 26908 27307 26911
rect 27430 26908 27436 26920
rect 27295 26880 27436 26908
rect 27295 26877 27307 26880
rect 27249 26871 27307 26877
rect 27430 26868 27436 26880
rect 27488 26908 27494 26920
rect 27632 26908 27660 26939
rect 27706 26936 27712 26988
rect 27764 26976 27770 26988
rect 28445 26979 28503 26985
rect 28445 26976 28457 26979
rect 27764 26948 28457 26976
rect 27764 26936 27770 26948
rect 28445 26945 28457 26948
rect 28491 26945 28503 26979
rect 28445 26939 28503 26945
rect 28810 26936 28816 26988
rect 28868 26936 28874 26988
rect 29089 26979 29147 26985
rect 29089 26945 29101 26979
rect 29135 26945 29147 26979
rect 29089 26939 29147 26945
rect 29273 26979 29331 26985
rect 29273 26945 29285 26979
rect 29319 26976 29331 26979
rect 29564 26976 29592 27072
rect 30184 27047 30242 27053
rect 30184 27013 30196 27047
rect 30230 27044 30242 27047
rect 30300 27044 30328 27072
rect 30230 27016 30328 27044
rect 30230 27013 30242 27016
rect 30184 27007 30242 27013
rect 32950 27004 32956 27056
rect 33008 27044 33014 27056
rect 33008 27016 34008 27044
rect 33008 27004 33014 27016
rect 29319 26948 29592 26976
rect 29319 26945 29331 26948
rect 29273 26939 29331 26945
rect 27488 26880 27660 26908
rect 29104 26908 29132 26939
rect 32398 26936 32404 26988
rect 32456 26976 32462 26988
rect 32841 26979 32899 26985
rect 32841 26976 32853 26979
rect 32456 26948 32853 26976
rect 32456 26936 32462 26948
rect 32841 26945 32853 26948
rect 32887 26945 32899 26979
rect 32841 26939 32899 26945
rect 29917 26911 29975 26917
rect 29104 26880 29776 26908
rect 27488 26868 27494 26880
rect 26804 26812 27476 26840
rect 25516 26772 25544 26800
rect 27448 26781 27476 26812
rect 24044 26744 25544 26772
rect 27433 26775 27491 26781
rect 27433 26741 27445 26775
rect 27479 26772 27491 26775
rect 29104 26772 29132 26880
rect 29748 26784 29776 26880
rect 29917 26877 29929 26911
rect 29963 26877 29975 26911
rect 32585 26911 32643 26917
rect 32585 26908 32597 26911
rect 29917 26871 29975 26877
rect 30944 26880 32597 26908
rect 27479 26744 29132 26772
rect 27479 26741 27491 26744
rect 27433 26735 27491 26741
rect 29730 26732 29736 26784
rect 29788 26732 29794 26784
rect 29932 26772 29960 26871
rect 30282 26772 30288 26784
rect 29932 26744 30288 26772
rect 30282 26732 30288 26744
rect 30340 26772 30346 26784
rect 30944 26772 30972 26880
rect 32585 26877 32597 26880
rect 32631 26877 32643 26911
rect 32585 26871 32643 26877
rect 30340 26744 30972 26772
rect 31297 26775 31355 26781
rect 30340 26732 30346 26744
rect 31297 26741 31309 26775
rect 31343 26772 31355 26775
rect 31478 26772 31484 26784
rect 31343 26744 31484 26772
rect 31343 26741 31355 26744
rect 31297 26735 31355 26741
rect 31478 26732 31484 26744
rect 31536 26732 31542 26784
rect 32600 26772 32628 26871
rect 33980 26849 34008 27016
rect 34609 26911 34667 26917
rect 34609 26877 34621 26911
rect 34655 26877 34667 26911
rect 34609 26871 34667 26877
rect 33965 26843 34023 26849
rect 33965 26809 33977 26843
rect 34011 26840 34023 26843
rect 34624 26840 34652 26871
rect 34011 26812 34652 26840
rect 34011 26809 34023 26812
rect 33965 26803 34023 26809
rect 33778 26772 33784 26784
rect 32600 26744 33784 26772
rect 33778 26732 33784 26744
rect 33836 26732 33842 26784
rect 34054 26732 34060 26784
rect 34112 26732 34118 26784
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 18141 26571 18199 26577
rect 18141 26537 18153 26571
rect 18187 26568 18199 26571
rect 18322 26568 18328 26580
rect 18187 26540 18328 26568
rect 18187 26537 18199 26540
rect 18141 26531 18199 26537
rect 18322 26528 18328 26540
rect 18380 26528 18386 26580
rect 18782 26528 18788 26580
rect 18840 26528 18846 26580
rect 19702 26528 19708 26580
rect 19760 26528 19766 26580
rect 19794 26528 19800 26580
rect 19852 26528 19858 26580
rect 20438 26568 20444 26580
rect 19996 26540 20444 26568
rect 19334 26460 19340 26512
rect 19392 26500 19398 26512
rect 19521 26503 19579 26509
rect 19521 26500 19533 26503
rect 19392 26472 19533 26500
rect 19392 26460 19398 26472
rect 19521 26469 19533 26472
rect 19567 26469 19579 26503
rect 19521 26463 19579 26469
rect 12161 26367 12219 26373
rect 12161 26333 12173 26367
rect 12207 26333 12219 26367
rect 12161 26327 12219 26333
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26364 14335 26367
rect 14323 26336 16252 26364
rect 14323 26333 14335 26336
rect 14277 26327 14335 26333
rect 10410 26256 10416 26308
rect 10468 26296 10474 26308
rect 12176 26296 12204 26327
rect 10468 26268 12388 26296
rect 10468 26256 10474 26268
rect 12360 26228 12388 26268
rect 12434 26256 12440 26308
rect 12492 26256 12498 26308
rect 14185 26299 14243 26305
rect 14185 26296 14197 26299
rect 13662 26268 14197 26296
rect 14185 26265 14197 26268
rect 14231 26265 14243 26299
rect 14185 26259 14243 26265
rect 16224 26240 16252 26336
rect 18230 26324 18236 26376
rect 18288 26324 18294 26376
rect 19720 26373 19748 26528
rect 19996 26373 20024 26540
rect 20438 26528 20444 26540
rect 20496 26528 20502 26580
rect 20530 26528 20536 26580
rect 20588 26528 20594 26580
rect 20806 26528 20812 26580
rect 20864 26528 20870 26580
rect 21361 26571 21419 26577
rect 21361 26537 21373 26571
rect 21407 26568 21419 26571
rect 21634 26568 21640 26580
rect 21407 26540 21640 26568
rect 21407 26537 21419 26540
rect 21361 26531 21419 26537
rect 21634 26528 21640 26540
rect 21692 26528 21698 26580
rect 22738 26528 22744 26580
rect 22796 26528 22802 26580
rect 23109 26571 23167 26577
rect 23109 26537 23121 26571
rect 23155 26568 23167 26571
rect 23474 26568 23480 26580
rect 23155 26540 23480 26568
rect 23155 26537 23167 26540
rect 23109 26531 23167 26537
rect 23474 26528 23480 26540
rect 23532 26528 23538 26580
rect 25317 26571 25375 26577
rect 25317 26537 25329 26571
rect 25363 26568 25375 26571
rect 25498 26568 25504 26580
rect 25363 26540 25504 26568
rect 25363 26537 25375 26540
rect 25317 26531 25375 26537
rect 25498 26528 25504 26540
rect 25556 26528 25562 26580
rect 27430 26528 27436 26580
rect 27488 26528 27494 26580
rect 27706 26528 27712 26580
rect 27764 26528 27770 26580
rect 28534 26528 28540 26580
rect 28592 26528 28598 26580
rect 28810 26528 28816 26580
rect 28868 26568 28874 26580
rect 29549 26571 29607 26577
rect 29549 26568 29561 26571
rect 28868 26540 29561 26568
rect 28868 26528 28874 26540
rect 29549 26537 29561 26540
rect 29595 26537 29607 26571
rect 33505 26571 33563 26577
rect 33505 26568 33517 26571
rect 29549 26531 29607 26537
rect 33152 26540 33517 26568
rect 20548 26432 20576 26528
rect 20824 26500 20852 26528
rect 21821 26503 21879 26509
rect 21821 26500 21833 26503
rect 20824 26472 21833 26500
rect 21821 26469 21833 26472
rect 21867 26469 21879 26503
rect 21821 26463 21879 26469
rect 23290 26460 23296 26512
rect 23348 26460 23354 26512
rect 27724 26500 27752 26528
rect 28169 26503 28227 26509
rect 28169 26500 28181 26503
rect 27724 26472 28181 26500
rect 28169 26469 28181 26472
rect 28215 26469 28227 26503
rect 31849 26503 31907 26509
rect 31849 26500 31861 26503
rect 28169 26463 28227 26469
rect 30576 26472 31861 26500
rect 21174 26432 21180 26444
rect 20180 26404 20576 26432
rect 20824 26404 21180 26432
rect 20180 26373 20208 26404
rect 18693 26367 18751 26373
rect 18693 26333 18705 26367
rect 18739 26364 18751 26367
rect 19429 26367 19487 26373
rect 19429 26364 19441 26367
rect 18739 26336 19441 26364
rect 18739 26333 18751 26336
rect 18693 26327 18751 26333
rect 19429 26333 19441 26336
rect 19475 26364 19487 26367
rect 19705 26367 19763 26373
rect 19475 26336 19564 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 19337 26299 19395 26305
rect 19337 26265 19349 26299
rect 19383 26296 19395 26299
rect 19536 26296 19564 26336
rect 19705 26333 19717 26367
rect 19751 26333 19763 26367
rect 19705 26327 19763 26333
rect 19981 26367 20039 26373
rect 19981 26333 19993 26367
rect 20027 26333 20039 26367
rect 19981 26327 20039 26333
rect 20165 26367 20223 26373
rect 20165 26333 20177 26367
rect 20211 26333 20223 26367
rect 20165 26327 20223 26333
rect 20254 26324 20260 26376
rect 20312 26364 20318 26376
rect 20824 26373 20852 26404
rect 21174 26392 21180 26404
rect 21232 26392 21238 26444
rect 21266 26392 21272 26444
rect 21324 26432 21330 26444
rect 21324 26404 21864 26432
rect 21324 26392 21330 26404
rect 20625 26367 20683 26373
rect 20625 26364 20637 26367
rect 20312 26336 20637 26364
rect 20312 26324 20318 26336
rect 20625 26333 20637 26336
rect 20671 26333 20683 26367
rect 20625 26327 20683 26333
rect 20809 26367 20867 26373
rect 20809 26333 20821 26367
rect 20855 26333 20867 26367
rect 20809 26327 20867 26333
rect 21085 26367 21143 26373
rect 21085 26333 21097 26367
rect 21131 26364 21143 26367
rect 21284 26364 21312 26392
rect 21131 26336 21312 26364
rect 21131 26333 21143 26336
rect 21085 26327 21143 26333
rect 21542 26324 21548 26376
rect 21600 26324 21606 26376
rect 21634 26324 21640 26376
rect 21692 26324 21698 26376
rect 21836 26373 21864 26404
rect 21729 26367 21787 26373
rect 21729 26333 21741 26367
rect 21775 26333 21787 26367
rect 21729 26327 21787 26333
rect 21821 26367 21879 26373
rect 21821 26333 21833 26367
rect 21867 26333 21879 26367
rect 21821 26327 21879 26333
rect 20070 26296 20076 26308
rect 19383 26268 19472 26296
rect 19536 26268 20076 26296
rect 19383 26265 19395 26268
rect 19337 26259 19395 26265
rect 19444 26240 19472 26268
rect 20070 26256 20076 26268
rect 20128 26256 20134 26308
rect 20993 26299 21051 26305
rect 20993 26265 21005 26299
rect 21039 26296 21051 26299
rect 21652 26296 21680 26324
rect 21039 26268 21680 26296
rect 21039 26265 21051 26268
rect 20993 26259 21051 26265
rect 13814 26228 13820 26240
rect 12360 26200 13820 26228
rect 13814 26188 13820 26200
rect 13872 26188 13878 26240
rect 13906 26188 13912 26240
rect 13964 26188 13970 26240
rect 16206 26188 16212 26240
rect 16264 26188 16270 26240
rect 19426 26188 19432 26240
rect 19484 26188 19490 26240
rect 21744 26228 21772 26327
rect 22002 26324 22008 26376
rect 22060 26324 22066 26376
rect 22186 26324 22192 26376
rect 22244 26364 22250 26376
rect 22833 26367 22891 26373
rect 22833 26364 22845 26367
rect 22244 26336 22845 26364
rect 22244 26324 22250 26336
rect 22833 26333 22845 26336
rect 22879 26333 22891 26367
rect 22833 26327 22891 26333
rect 22925 26367 22983 26373
rect 22925 26333 22937 26367
rect 22971 26364 22983 26367
rect 23308 26364 23336 26460
rect 23658 26392 23664 26444
rect 23716 26432 23722 26444
rect 25406 26432 25412 26444
rect 23716 26404 25412 26432
rect 23716 26392 23722 26404
rect 25406 26392 25412 26404
rect 25464 26392 25470 26444
rect 27080 26404 30144 26432
rect 27080 26376 27108 26404
rect 22971 26336 23336 26364
rect 25133 26367 25191 26373
rect 22971 26333 22983 26336
rect 22925 26327 22983 26333
rect 25133 26333 25145 26367
rect 25179 26364 25191 26367
rect 25314 26364 25320 26376
rect 25179 26336 25320 26364
rect 25179 26333 25191 26336
rect 25133 26327 25191 26333
rect 22462 26256 22468 26308
rect 22520 26296 22526 26308
rect 22649 26299 22707 26305
rect 22649 26296 22661 26299
rect 22520 26268 22661 26296
rect 22520 26256 22526 26268
rect 22649 26265 22661 26268
rect 22695 26265 22707 26299
rect 22649 26259 22707 26265
rect 22738 26256 22744 26308
rect 22796 26296 22802 26308
rect 25148 26296 25176 26327
rect 25314 26324 25320 26336
rect 25372 26364 25378 26376
rect 25590 26364 25596 26376
rect 25372 26336 25596 26364
rect 25372 26324 25378 26336
rect 25590 26324 25596 26336
rect 25648 26324 25654 26376
rect 27062 26324 27068 26376
rect 27120 26324 27126 26376
rect 27709 26367 27767 26373
rect 27709 26333 27721 26367
rect 27755 26364 27767 26367
rect 27798 26364 27804 26376
rect 27755 26336 27804 26364
rect 27755 26333 27767 26336
rect 27709 26327 27767 26333
rect 27798 26324 27804 26336
rect 27856 26324 27862 26376
rect 29730 26324 29736 26376
rect 29788 26324 29794 26376
rect 30116 26373 30144 26404
rect 30466 26392 30472 26444
rect 30524 26392 30530 26444
rect 29825 26367 29883 26373
rect 29825 26333 29837 26367
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 30009 26367 30067 26373
rect 30009 26333 30021 26367
rect 30055 26333 30067 26367
rect 30009 26327 30067 26333
rect 30101 26367 30159 26373
rect 30101 26333 30113 26367
rect 30147 26364 30159 26367
rect 30484 26364 30512 26392
rect 30576 26373 30604 26472
rect 31849 26469 31861 26472
rect 31895 26469 31907 26503
rect 33152 26500 33180 26540
rect 33505 26537 33517 26540
rect 33551 26537 33563 26571
rect 33505 26531 33563 26537
rect 34054 26528 34060 26580
rect 34112 26528 34118 26580
rect 31849 26463 31907 26469
rect 32324 26472 33180 26500
rect 31297 26435 31355 26441
rect 31297 26432 31309 26435
rect 30668 26404 31309 26432
rect 30668 26373 30696 26404
rect 31297 26401 31309 26404
rect 31343 26401 31355 26435
rect 31297 26395 31355 26401
rect 31496 26404 31892 26432
rect 31496 26376 31524 26404
rect 30147 26336 30512 26364
rect 30561 26367 30619 26373
rect 30147 26333 30159 26336
rect 30101 26327 30159 26333
rect 30561 26333 30573 26367
rect 30607 26333 30619 26367
rect 30561 26327 30619 26333
rect 30653 26367 30711 26373
rect 30653 26333 30665 26367
rect 30699 26333 30711 26367
rect 30653 26327 30711 26333
rect 31021 26367 31079 26373
rect 31021 26333 31033 26367
rect 31067 26364 31079 26367
rect 31478 26364 31484 26376
rect 31067 26336 31484 26364
rect 31067 26333 31079 26336
rect 31021 26327 31079 26333
rect 22796 26268 25176 26296
rect 27985 26299 28043 26305
rect 22796 26256 22802 26268
rect 27985 26265 27997 26299
rect 28031 26296 28043 26299
rect 28074 26296 28080 26308
rect 28031 26268 28080 26296
rect 28031 26265 28043 26268
rect 27985 26259 28043 26265
rect 28074 26256 28080 26268
rect 28132 26256 28138 26308
rect 28537 26299 28595 26305
rect 28537 26265 28549 26299
rect 28583 26296 28595 26299
rect 29362 26296 29368 26308
rect 28583 26268 29368 26296
rect 28583 26265 28595 26268
rect 28537 26259 28595 26265
rect 29362 26256 29368 26268
rect 29420 26296 29426 26308
rect 29840 26296 29868 26327
rect 29420 26268 29868 26296
rect 29420 26256 29426 26268
rect 21818 26228 21824 26240
rect 21744 26200 21824 26228
rect 21818 26188 21824 26200
rect 21876 26228 21882 26240
rect 23106 26228 23112 26240
rect 21876 26200 23112 26228
rect 21876 26188 21882 26200
rect 23106 26188 23112 26200
rect 23164 26188 23170 26240
rect 24946 26188 24952 26240
rect 25004 26188 25010 26240
rect 27617 26231 27675 26237
rect 27617 26197 27629 26231
rect 27663 26228 27675 26231
rect 27706 26228 27712 26240
rect 27663 26200 27712 26228
rect 27663 26197 27675 26200
rect 27617 26191 27675 26197
rect 27706 26188 27712 26200
rect 27764 26188 27770 26240
rect 27801 26231 27859 26237
rect 27801 26197 27813 26231
rect 27847 26228 27859 26231
rect 27890 26228 27896 26240
rect 27847 26200 27896 26228
rect 27847 26197 27859 26200
rect 27801 26191 27859 26197
rect 27890 26188 27896 26200
rect 27948 26188 27954 26240
rect 28718 26188 28724 26240
rect 28776 26188 28782 26240
rect 29270 26188 29276 26240
rect 29328 26228 29334 26240
rect 30024 26228 30052 26327
rect 31478 26324 31484 26336
rect 31536 26324 31542 26376
rect 31754 26324 31760 26376
rect 31812 26324 31818 26376
rect 31864 26373 31892 26404
rect 32324 26373 32352 26472
rect 32398 26392 32404 26444
rect 32456 26392 32462 26444
rect 32585 26435 32643 26441
rect 32585 26432 32597 26435
rect 32508 26404 32597 26432
rect 32508 26373 32536 26404
rect 32585 26401 32597 26404
rect 32631 26401 32643 26435
rect 32585 26395 32643 26401
rect 32950 26392 32956 26444
rect 33008 26392 33014 26444
rect 33042 26392 33048 26444
rect 33100 26432 33106 26444
rect 33870 26432 33876 26444
rect 33100 26404 33876 26432
rect 33100 26392 33106 26404
rect 33870 26392 33876 26404
rect 33928 26392 33934 26444
rect 31849 26367 31907 26373
rect 31849 26333 31861 26367
rect 31895 26333 31907 26367
rect 31849 26327 31907 26333
rect 31941 26367 31999 26373
rect 31941 26333 31953 26367
rect 31987 26364 31999 26367
rect 32309 26367 32367 26373
rect 31987 26336 32260 26364
rect 31987 26333 31999 26336
rect 31941 26327 31999 26333
rect 30742 26256 30748 26308
rect 30800 26256 30806 26308
rect 30926 26305 30932 26308
rect 30883 26299 30932 26305
rect 30883 26265 30895 26299
rect 30929 26265 30932 26299
rect 30883 26259 30932 26265
rect 30926 26256 30932 26259
rect 30984 26256 30990 26308
rect 31956 26296 31984 26327
rect 31680 26268 31984 26296
rect 32125 26299 32183 26305
rect 29328 26200 30052 26228
rect 30377 26231 30435 26237
rect 29328 26188 29334 26200
rect 30377 26197 30389 26231
rect 30423 26228 30435 26231
rect 30466 26228 30472 26240
rect 30423 26200 30472 26228
rect 30423 26197 30435 26200
rect 30377 26191 30435 26197
rect 30466 26188 30472 26200
rect 30524 26188 30530 26240
rect 31202 26188 31208 26240
rect 31260 26228 31266 26240
rect 31680 26237 31708 26268
rect 32125 26265 32137 26299
rect 32171 26265 32183 26299
rect 32232 26296 32260 26336
rect 32309 26333 32321 26367
rect 32355 26333 32367 26367
rect 32309 26327 32367 26333
rect 32493 26367 32551 26373
rect 32493 26333 32505 26367
rect 32539 26333 32551 26367
rect 32493 26327 32551 26333
rect 32674 26324 32680 26376
rect 32732 26364 32738 26376
rect 32769 26367 32827 26373
rect 32769 26364 32781 26367
rect 32732 26336 32781 26364
rect 32732 26324 32738 26336
rect 32769 26333 32781 26336
rect 32815 26333 32827 26367
rect 32769 26327 32827 26333
rect 32858 26324 32864 26376
rect 32916 26324 32922 26376
rect 32968 26296 32996 26392
rect 33229 26367 33287 26373
rect 33229 26364 33241 26367
rect 32232 26268 32996 26296
rect 33060 26336 33241 26364
rect 32125 26259 32183 26265
rect 31665 26231 31723 26237
rect 31665 26228 31677 26231
rect 31260 26200 31677 26228
rect 31260 26188 31266 26200
rect 31665 26197 31677 26200
rect 31711 26197 31723 26231
rect 31665 26191 31723 26197
rect 31754 26188 31760 26240
rect 31812 26228 31818 26240
rect 32140 26228 32168 26259
rect 32214 26228 32220 26240
rect 31812 26200 32220 26228
rect 31812 26188 31818 26200
rect 32214 26188 32220 26200
rect 32272 26228 32278 26240
rect 32674 26228 32680 26240
rect 32272 26200 32680 26228
rect 32272 26188 32278 26200
rect 32674 26188 32680 26200
rect 32732 26228 32738 26240
rect 33060 26228 33088 26336
rect 33229 26333 33241 26336
rect 33275 26333 33287 26367
rect 33229 26327 33287 26333
rect 33505 26367 33563 26373
rect 33505 26333 33517 26367
rect 33551 26364 33563 26367
rect 34072 26364 34100 26528
rect 33551 26336 34100 26364
rect 33551 26333 33563 26336
rect 33505 26327 33563 26333
rect 33318 26256 33324 26308
rect 33376 26256 33382 26308
rect 32732 26200 33088 26228
rect 32732 26188 32738 26200
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 12345 26027 12403 26033
rect 12345 25993 12357 26027
rect 12391 25993 12403 26027
rect 19334 26024 19340 26036
rect 12345 25987 12403 25993
rect 18432 25996 19340 26024
rect 11977 25891 12035 25897
rect 11977 25857 11989 25891
rect 12023 25888 12035 25891
rect 12360 25888 12388 25987
rect 16298 25956 16304 25968
rect 15502 25928 16304 25956
rect 16298 25916 16304 25928
rect 16356 25916 16362 25968
rect 18432 25965 18460 25996
rect 19334 25984 19340 25996
rect 19392 25984 19398 26036
rect 19889 26027 19947 26033
rect 19889 25993 19901 26027
rect 19935 25993 19947 26027
rect 19889 25987 19947 25993
rect 18417 25959 18475 25965
rect 18417 25925 18429 25959
rect 18463 25925 18475 25959
rect 18417 25919 18475 25925
rect 19426 25916 19432 25968
rect 19484 25916 19490 25968
rect 19904 25956 19932 25987
rect 21174 25984 21180 26036
rect 21232 25984 21238 26036
rect 21542 25984 21548 26036
rect 21600 25984 21606 26036
rect 21913 26027 21971 26033
rect 21913 25993 21925 26027
rect 21959 26024 21971 26027
rect 22002 26024 22008 26036
rect 21959 25996 22008 26024
rect 21959 25993 21971 25996
rect 21913 25987 21971 25993
rect 22002 25984 22008 25996
rect 22060 25984 22066 26036
rect 22646 25984 22652 26036
rect 22704 25984 22710 26036
rect 25498 25984 25504 26036
rect 25556 25984 25562 26036
rect 28261 26027 28319 26033
rect 28261 25993 28273 26027
rect 28307 26024 28319 26027
rect 28534 26024 28540 26036
rect 28307 25996 28540 26024
rect 28307 25993 28319 25996
rect 28261 25987 28319 25993
rect 28534 25984 28540 25996
rect 28592 25984 28598 26036
rect 30466 25984 30472 26036
rect 30524 25984 30530 26036
rect 20346 25956 20352 25968
rect 19904 25928 20352 25956
rect 20346 25916 20352 25928
rect 20404 25956 20410 25968
rect 20809 25959 20867 25965
rect 20809 25956 20821 25959
rect 20404 25928 20821 25956
rect 20404 25916 20410 25928
rect 20809 25925 20821 25928
rect 20855 25925 20867 25959
rect 21560 25956 21588 25984
rect 21560 25928 22048 25956
rect 20809 25919 20867 25925
rect 12023 25860 12388 25888
rect 12023 25857 12035 25860
rect 11977 25851 12035 25857
rect 12710 25848 12716 25900
rect 12768 25848 12774 25900
rect 13814 25848 13820 25900
rect 13872 25888 13878 25900
rect 14001 25891 14059 25897
rect 14001 25888 14013 25891
rect 13872 25860 14013 25888
rect 13872 25848 13878 25860
rect 14001 25857 14013 25860
rect 14047 25857 14059 25891
rect 14001 25851 14059 25857
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18141 25891 18199 25897
rect 18141 25888 18153 25891
rect 18012 25860 18153 25888
rect 18012 25848 18018 25860
rect 18141 25857 18153 25860
rect 18187 25857 18199 25891
rect 18141 25851 18199 25857
rect 20622 25848 20628 25900
rect 20680 25848 20686 25900
rect 21361 25891 21419 25897
rect 21361 25857 21373 25891
rect 21407 25857 21419 25891
rect 21361 25851 21419 25857
rect 12802 25780 12808 25832
rect 12860 25780 12866 25832
rect 12989 25823 13047 25829
rect 12989 25789 13001 25823
rect 13035 25820 13047 25823
rect 13906 25820 13912 25832
rect 13035 25792 13912 25820
rect 13035 25789 13047 25792
rect 12989 25783 13047 25789
rect 13906 25780 13912 25792
rect 13964 25780 13970 25832
rect 14274 25780 14280 25832
rect 14332 25780 14338 25832
rect 21376 25820 21404 25851
rect 21542 25848 21548 25900
rect 21600 25848 21606 25900
rect 21818 25848 21824 25900
rect 21876 25848 21882 25900
rect 21910 25848 21916 25900
rect 21968 25848 21974 25900
rect 22020 25897 22048 25928
rect 22005 25891 22063 25897
rect 22005 25857 22017 25891
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 21928 25820 21956 25848
rect 21376 25792 21956 25820
rect 12161 25755 12219 25761
rect 12161 25721 12173 25755
rect 12207 25752 12219 25755
rect 12434 25752 12440 25764
rect 12207 25724 12440 25752
rect 12207 25721 12219 25724
rect 12161 25715 12219 25721
rect 12434 25712 12440 25724
rect 12492 25712 12498 25764
rect 22020 25752 22048 25851
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22557 25891 22615 25897
rect 22557 25888 22569 25891
rect 22152 25860 22569 25888
rect 22152 25848 22158 25860
rect 22557 25857 22569 25860
rect 22603 25857 22615 25891
rect 22557 25851 22615 25857
rect 22738 25848 22744 25900
rect 22796 25848 22802 25900
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25888 23351 25891
rect 23842 25888 23848 25900
rect 23339 25860 23848 25888
rect 23339 25857 23351 25860
rect 23293 25851 23351 25857
rect 23842 25848 23848 25860
rect 23900 25848 23906 25900
rect 24762 25848 24768 25900
rect 24820 25848 24826 25900
rect 24946 25848 24952 25900
rect 25004 25848 25010 25900
rect 25130 25848 25136 25900
rect 25188 25848 25194 25900
rect 25516 25888 25544 25984
rect 27062 25956 27068 25968
rect 26252 25928 27068 25956
rect 26252 25900 26280 25928
rect 27062 25916 27068 25928
rect 27120 25956 27126 25968
rect 28077 25959 28135 25965
rect 28077 25956 28089 25959
rect 27120 25928 27200 25956
rect 27120 25916 27126 25928
rect 25685 25891 25743 25897
rect 25685 25888 25697 25891
rect 25516 25860 25697 25888
rect 25685 25857 25697 25860
rect 25731 25857 25743 25891
rect 25685 25851 25743 25857
rect 26234 25848 26240 25900
rect 26292 25848 26298 25900
rect 27172 25897 27200 25928
rect 27908 25928 28089 25956
rect 27908 25900 27936 25928
rect 28077 25925 28089 25928
rect 28123 25925 28135 25959
rect 28077 25919 28135 25925
rect 26789 25891 26847 25897
rect 26789 25857 26801 25891
rect 26835 25888 26847 25891
rect 27157 25891 27215 25897
rect 26835 25860 27016 25888
rect 26835 25857 26847 25860
rect 26789 25851 26847 25857
rect 25038 25780 25044 25832
rect 25096 25780 25102 25832
rect 25314 25780 25320 25832
rect 25372 25820 25378 25832
rect 25409 25823 25467 25829
rect 25409 25820 25421 25823
rect 25372 25792 25421 25820
rect 25372 25780 25378 25792
rect 25409 25789 25421 25792
rect 25455 25789 25467 25823
rect 25409 25783 25467 25789
rect 25225 25755 25283 25761
rect 22020 25724 23152 25752
rect 15746 25644 15752 25696
rect 15804 25644 15810 25696
rect 20993 25687 21051 25693
rect 20993 25653 21005 25687
rect 21039 25684 21051 25687
rect 22186 25684 22192 25696
rect 21039 25656 22192 25684
rect 21039 25653 21051 25656
rect 20993 25647 21051 25653
rect 22186 25644 22192 25656
rect 22244 25644 22250 25696
rect 23124 25693 23152 25724
rect 25225 25721 25237 25755
rect 25271 25752 25283 25755
rect 25590 25752 25596 25764
rect 25271 25724 25596 25752
rect 25271 25721 25283 25724
rect 25225 25715 25283 25721
rect 25590 25712 25596 25724
rect 25648 25712 25654 25764
rect 26988 25761 27016 25860
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 27341 25891 27399 25897
rect 27341 25857 27353 25891
rect 27387 25888 27399 25891
rect 27430 25888 27436 25900
rect 27387 25860 27436 25888
rect 27387 25857 27399 25860
rect 27341 25851 27399 25857
rect 27430 25848 27436 25860
rect 27488 25848 27494 25900
rect 27614 25848 27620 25900
rect 27672 25848 27678 25900
rect 27706 25848 27712 25900
rect 27764 25848 27770 25900
rect 27890 25848 27896 25900
rect 27948 25848 27954 25900
rect 29178 25848 29184 25900
rect 29236 25848 29242 25900
rect 30101 25891 30159 25897
rect 30101 25857 30113 25891
rect 30147 25888 30159 25891
rect 30484 25888 30512 25984
rect 30147 25860 30512 25888
rect 30147 25857 30159 25860
rect 30101 25851 30159 25857
rect 31202 25848 31208 25900
rect 31260 25848 31266 25900
rect 31297 25891 31355 25897
rect 31297 25857 31309 25891
rect 31343 25888 31355 25891
rect 31478 25888 31484 25900
rect 31343 25860 31484 25888
rect 31343 25857 31355 25860
rect 31297 25851 31355 25857
rect 31478 25848 31484 25860
rect 31536 25848 31542 25900
rect 29914 25820 29920 25832
rect 27172 25792 29920 25820
rect 27172 25764 27200 25792
rect 29914 25780 29920 25792
rect 29972 25780 29978 25832
rect 30285 25823 30343 25829
rect 30285 25789 30297 25823
rect 30331 25820 30343 25823
rect 30558 25820 30564 25832
rect 30331 25792 30564 25820
rect 30331 25789 30343 25792
rect 30285 25783 30343 25789
rect 30558 25780 30564 25792
rect 30616 25780 30622 25832
rect 31110 25780 31116 25832
rect 31168 25780 31174 25832
rect 26973 25755 27031 25761
rect 26973 25721 26985 25755
rect 27019 25721 27031 25755
rect 26973 25715 27031 25721
rect 27154 25712 27160 25764
rect 27212 25712 27218 25764
rect 27540 25724 28764 25752
rect 23109 25687 23167 25693
rect 23109 25653 23121 25687
rect 23155 25684 23167 25687
rect 23198 25684 23204 25696
rect 23155 25656 23204 25684
rect 23155 25653 23167 25656
rect 23109 25647 23167 25653
rect 23198 25644 23204 25656
rect 23256 25644 23262 25696
rect 24026 25644 24032 25696
rect 24084 25684 24090 25696
rect 24581 25687 24639 25693
rect 24581 25684 24593 25687
rect 24084 25656 24593 25684
rect 24084 25644 24090 25656
rect 24581 25653 24593 25656
rect 24627 25653 24639 25687
rect 24581 25647 24639 25653
rect 25314 25644 25320 25696
rect 25372 25644 25378 25696
rect 26694 25644 26700 25696
rect 26752 25644 26758 25696
rect 27540 25693 27568 25724
rect 27525 25687 27583 25693
rect 27525 25653 27537 25687
rect 27571 25653 27583 25687
rect 27525 25647 27583 25653
rect 27798 25644 27804 25696
rect 27856 25684 27862 25696
rect 28077 25687 28135 25693
rect 28077 25684 28089 25687
rect 27856 25656 28089 25684
rect 27856 25644 27862 25656
rect 28077 25653 28089 25656
rect 28123 25653 28135 25687
rect 28736 25684 28764 25724
rect 28810 25712 28816 25764
rect 28868 25752 28874 25764
rect 28868 25724 30696 25752
rect 28868 25712 28874 25724
rect 30668 25696 30696 25724
rect 29270 25684 29276 25696
rect 28736 25656 29276 25684
rect 28077 25647 28135 25653
rect 29270 25644 29276 25656
rect 29328 25644 29334 25696
rect 29362 25644 29368 25696
rect 29420 25644 29426 25696
rect 30650 25644 30656 25696
rect 30708 25684 30714 25696
rect 30929 25687 30987 25693
rect 30929 25684 30941 25687
rect 30708 25656 30941 25684
rect 30708 25644 30714 25656
rect 30929 25653 30941 25656
rect 30975 25653 30987 25687
rect 30929 25647 30987 25653
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 12710 25440 12716 25492
rect 12768 25480 12774 25492
rect 13633 25483 13691 25489
rect 13633 25480 13645 25483
rect 12768 25452 13645 25480
rect 12768 25440 12774 25452
rect 13633 25449 13645 25452
rect 13679 25449 13691 25483
rect 13633 25443 13691 25449
rect 14274 25440 14280 25492
rect 14332 25480 14338 25492
rect 14369 25483 14427 25489
rect 14369 25480 14381 25483
rect 14332 25452 14381 25480
rect 14332 25440 14338 25452
rect 14369 25449 14381 25452
rect 14415 25449 14427 25483
rect 14369 25443 14427 25449
rect 16298 25440 16304 25492
rect 16356 25440 16362 25492
rect 22830 25480 22836 25492
rect 22020 25452 22836 25480
rect 12618 25372 12624 25424
rect 12676 25412 12682 25424
rect 13449 25415 13507 25421
rect 13449 25412 13461 25415
rect 12676 25384 13461 25412
rect 12676 25372 12682 25384
rect 13449 25381 13461 25384
rect 13495 25412 13507 25415
rect 14645 25415 14703 25421
rect 13495 25384 13676 25412
rect 13495 25381 13507 25384
rect 13449 25375 13507 25381
rect 9766 25304 9772 25356
rect 9824 25344 9830 25356
rect 10137 25347 10195 25353
rect 10137 25344 10149 25347
rect 9824 25316 10149 25344
rect 9824 25304 9830 25316
rect 10137 25313 10149 25316
rect 10183 25344 10195 25347
rect 10410 25344 10416 25356
rect 10183 25316 10416 25344
rect 10183 25313 10195 25316
rect 10137 25307 10195 25313
rect 10410 25304 10416 25316
rect 10468 25344 10474 25356
rect 10962 25344 10968 25356
rect 10468 25316 10968 25344
rect 10468 25304 10474 25316
rect 10962 25304 10968 25316
rect 11020 25304 11026 25356
rect 11885 25347 11943 25353
rect 11885 25313 11897 25347
rect 11931 25344 11943 25347
rect 12713 25347 12771 25353
rect 12713 25344 12725 25347
rect 11931 25316 12725 25344
rect 11931 25313 11943 25316
rect 11885 25307 11943 25313
rect 12713 25313 12725 25316
rect 12759 25344 12771 25347
rect 12759 25316 13584 25344
rect 12759 25313 12771 25316
rect 12713 25307 12771 25313
rect 13280 25285 13308 25316
rect 13265 25279 13323 25285
rect 13265 25245 13277 25279
rect 13311 25245 13323 25279
rect 13265 25239 13323 25245
rect 13354 25236 13360 25288
rect 13412 25236 13418 25288
rect 13556 25285 13584 25316
rect 13648 25285 13676 25384
rect 14645 25381 14657 25415
rect 14691 25381 14703 25415
rect 14645 25375 14703 25381
rect 13998 25344 14004 25356
rect 13832 25316 14004 25344
rect 13832 25285 13860 25316
rect 13998 25304 14004 25316
rect 14056 25304 14062 25356
rect 13541 25279 13599 25285
rect 13541 25245 13553 25279
rect 13587 25245 13599 25279
rect 13541 25239 13599 25245
rect 13633 25279 13691 25285
rect 13633 25245 13645 25279
rect 13679 25245 13691 25279
rect 13633 25239 13691 25245
rect 13817 25279 13875 25285
rect 13817 25245 13829 25279
rect 13863 25245 13875 25279
rect 13817 25239 13875 25245
rect 13906 25236 13912 25288
rect 13964 25236 13970 25288
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25276 14611 25279
rect 14660 25276 14688 25375
rect 15289 25347 15347 25353
rect 15289 25313 15301 25347
rect 15335 25344 15347 25347
rect 15746 25344 15752 25356
rect 15335 25316 15752 25344
rect 15335 25313 15347 25316
rect 15289 25307 15347 25313
rect 15746 25304 15752 25316
rect 15804 25304 15810 25356
rect 17954 25304 17960 25356
rect 18012 25344 18018 25356
rect 19058 25344 19064 25356
rect 18012 25316 19064 25344
rect 18012 25304 18018 25316
rect 19058 25304 19064 25316
rect 19116 25344 19122 25356
rect 19245 25347 19303 25353
rect 19245 25344 19257 25347
rect 19116 25316 19257 25344
rect 19116 25304 19122 25316
rect 19245 25313 19257 25316
rect 19291 25313 19303 25347
rect 19245 25307 19303 25313
rect 14599 25248 14688 25276
rect 14599 25245 14611 25248
rect 14553 25239 14611 25245
rect 16022 25236 16028 25288
rect 16080 25236 16086 25288
rect 16393 25279 16451 25285
rect 16393 25276 16405 25279
rect 16224 25248 16405 25276
rect 10413 25211 10471 25217
rect 10413 25177 10425 25211
rect 10459 25177 10471 25211
rect 10413 25171 10471 25177
rect 10428 25140 10456 25171
rect 11146 25168 11152 25220
rect 11204 25168 11210 25220
rect 13081 25211 13139 25217
rect 13081 25177 13093 25211
rect 13127 25208 13139 25211
rect 13924 25208 13952 25236
rect 16224 25220 16252 25248
rect 16393 25245 16405 25248
rect 16439 25245 16451 25279
rect 16393 25239 16451 25245
rect 16666 25236 16672 25288
rect 16724 25276 16730 25288
rect 17972 25276 18000 25304
rect 16724 25248 18000 25276
rect 16724 25236 16730 25248
rect 18690 25236 18696 25288
rect 18748 25236 18754 25288
rect 22020 25285 22048 25452
rect 22830 25440 22836 25452
rect 22888 25480 22894 25492
rect 23290 25480 23296 25492
rect 22888 25452 23296 25480
rect 22888 25440 22894 25452
rect 23290 25440 23296 25452
rect 23348 25440 23354 25492
rect 23566 25440 23572 25492
rect 23624 25440 23630 25492
rect 24762 25440 24768 25492
rect 24820 25480 24826 25492
rect 25133 25483 25191 25489
rect 25133 25480 25145 25483
rect 24820 25452 25145 25480
rect 24820 25440 24826 25452
rect 25133 25449 25145 25452
rect 25179 25449 25191 25483
rect 25133 25443 25191 25449
rect 27525 25483 27583 25489
rect 27525 25449 27537 25483
rect 27571 25480 27583 25483
rect 27614 25480 27620 25492
rect 27571 25452 27620 25480
rect 27571 25449 27583 25452
rect 27525 25443 27583 25449
rect 27614 25440 27620 25452
rect 27672 25440 27678 25492
rect 29270 25440 29276 25492
rect 29328 25440 29334 25492
rect 29362 25440 29368 25492
rect 29420 25440 29426 25492
rect 31849 25483 31907 25489
rect 31849 25449 31861 25483
rect 31895 25480 31907 25483
rect 32125 25483 32183 25489
rect 32125 25480 32137 25483
rect 31895 25452 32137 25480
rect 31895 25449 31907 25452
rect 31849 25443 31907 25449
rect 32125 25449 32137 25452
rect 32171 25449 32183 25483
rect 32125 25443 32183 25449
rect 22738 25412 22744 25424
rect 22480 25384 22744 25412
rect 22097 25347 22155 25353
rect 22097 25313 22109 25347
rect 22143 25344 22155 25347
rect 22278 25344 22284 25356
rect 22143 25316 22284 25344
rect 22143 25313 22155 25316
rect 22097 25307 22155 25313
rect 22278 25304 22284 25316
rect 22336 25304 22342 25356
rect 22480 25344 22508 25384
rect 22738 25372 22744 25384
rect 22796 25412 22802 25424
rect 27433 25415 27491 25421
rect 22796 25384 24532 25412
rect 22796 25372 22802 25384
rect 24397 25347 24455 25353
rect 24397 25344 24409 25347
rect 22388 25316 22508 25344
rect 22572 25316 22968 25344
rect 22005 25279 22063 25285
rect 22005 25245 22017 25279
rect 22051 25245 22063 25279
rect 22005 25239 22063 25245
rect 22189 25279 22247 25285
rect 22189 25245 22201 25279
rect 22235 25276 22247 25279
rect 22388 25276 22416 25316
rect 22235 25248 22416 25276
rect 22465 25279 22523 25285
rect 22235 25245 22247 25248
rect 22189 25239 22247 25245
rect 22465 25245 22477 25279
rect 22511 25278 22523 25279
rect 22572 25278 22600 25316
rect 22511 25250 22600 25278
rect 22833 25279 22891 25285
rect 22511 25245 22523 25250
rect 22465 25239 22523 25245
rect 22833 25245 22845 25279
rect 22879 25245 22891 25279
rect 22833 25239 22891 25245
rect 13127 25180 13952 25208
rect 15013 25211 15071 25217
rect 13127 25177 13139 25180
rect 13081 25171 13139 25177
rect 15013 25177 15025 25211
rect 15059 25208 15071 25211
rect 15473 25211 15531 25217
rect 15473 25208 15485 25211
rect 15059 25180 15485 25208
rect 15059 25177 15071 25180
rect 15013 25171 15071 25177
rect 15473 25177 15485 25180
rect 15519 25177 15531 25211
rect 15473 25171 15531 25177
rect 16206 25168 16212 25220
rect 16264 25168 16270 25220
rect 16574 25168 16580 25220
rect 16632 25208 16638 25220
rect 16914 25211 16972 25217
rect 16914 25208 16926 25211
rect 16632 25180 16926 25208
rect 16632 25168 16638 25180
rect 16914 25177 16926 25180
rect 16960 25177 16972 25211
rect 16914 25171 16972 25177
rect 17954 25168 17960 25220
rect 18012 25208 18018 25220
rect 18141 25211 18199 25217
rect 18141 25208 18153 25211
rect 18012 25180 18153 25208
rect 18012 25168 18018 25180
rect 18141 25177 18153 25180
rect 18187 25177 18199 25211
rect 18141 25171 18199 25177
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 19521 25211 19579 25217
rect 19521 25208 19533 25211
rect 19484 25180 19533 25208
rect 19484 25168 19490 25180
rect 19521 25177 19533 25180
rect 19567 25177 19579 25211
rect 19521 25171 19579 25177
rect 19978 25168 19984 25220
rect 20036 25168 20042 25220
rect 21450 25168 21456 25220
rect 21508 25208 21514 25220
rect 21508 25180 22324 25208
rect 21508 25168 21514 25180
rect 11974 25140 11980 25152
rect 10428 25112 11980 25140
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12158 25100 12164 25152
rect 12216 25100 12222 25152
rect 12434 25100 12440 25152
rect 12492 25140 12498 25152
rect 12897 25143 12955 25149
rect 12897 25140 12909 25143
rect 12492 25112 12909 25140
rect 12492 25100 12498 25112
rect 12897 25109 12909 25112
rect 12943 25109 12955 25143
rect 12897 25103 12955 25109
rect 15105 25143 15163 25149
rect 15105 25109 15117 25143
rect 15151 25140 15163 25143
rect 16482 25140 16488 25152
rect 15151 25112 16488 25140
rect 15151 25109 15163 25112
rect 15105 25103 15163 25109
rect 16482 25100 16488 25112
rect 16540 25100 16546 25152
rect 18046 25100 18052 25152
rect 18104 25100 18110 25152
rect 20806 25100 20812 25152
rect 20864 25140 20870 25152
rect 22296 25149 22324 25180
rect 22554 25168 22560 25220
rect 22612 25168 22618 25220
rect 22646 25168 22652 25220
rect 22704 25168 22710 25220
rect 20993 25143 21051 25149
rect 20993 25140 21005 25143
rect 20864 25112 21005 25140
rect 20864 25100 20870 25112
rect 20993 25109 21005 25112
rect 21039 25109 21051 25143
rect 20993 25103 21051 25109
rect 22281 25143 22339 25149
rect 22281 25109 22293 25143
rect 22327 25109 22339 25143
rect 22848 25140 22876 25239
rect 22940 25208 22968 25316
rect 23032 25316 24409 25344
rect 23032 25285 23060 25316
rect 24397 25313 24409 25316
rect 24443 25313 24455 25347
rect 24397 25307 24455 25313
rect 23017 25279 23075 25285
rect 23017 25245 23029 25279
rect 23063 25245 23075 25279
rect 23017 25239 23075 25245
rect 23290 25236 23296 25288
rect 23348 25236 23354 25288
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25276 23443 25279
rect 23845 25279 23903 25285
rect 23431 25248 23704 25276
rect 23431 25245 23443 25248
rect 23385 25239 23443 25245
rect 23676 25220 23704 25248
rect 23845 25245 23857 25279
rect 23891 25276 23903 25279
rect 24210 25276 24216 25288
rect 23891 25248 24216 25276
rect 23891 25245 23903 25248
rect 23845 25239 23903 25245
rect 24210 25236 24216 25248
rect 24268 25236 24274 25288
rect 24504 25276 24532 25384
rect 27433 25381 27445 25415
rect 27479 25412 27491 25415
rect 27890 25412 27896 25424
rect 27479 25384 27896 25412
rect 27479 25381 27491 25384
rect 27433 25375 27491 25381
rect 27890 25372 27896 25384
rect 27948 25372 27954 25424
rect 24854 25304 24860 25356
rect 24912 25344 24918 25356
rect 26050 25344 26056 25356
rect 24912 25316 26056 25344
rect 24912 25304 24918 25316
rect 26050 25304 26056 25316
rect 26108 25304 26114 25356
rect 27706 25304 27712 25356
rect 27764 25304 27770 25356
rect 27908 25344 27936 25372
rect 27985 25347 28043 25353
rect 27985 25344 27997 25347
rect 27908 25316 27997 25344
rect 27985 25313 27997 25316
rect 28031 25313 28043 25347
rect 27985 25307 28043 25313
rect 28074 25304 28080 25356
rect 28132 25304 28138 25356
rect 28718 25344 28724 25356
rect 28644 25316 28724 25344
rect 24949 25279 25007 25285
rect 24949 25276 24961 25279
rect 24504 25248 24961 25276
rect 24949 25245 24961 25248
rect 24995 25276 25007 25279
rect 25038 25276 25044 25288
rect 24995 25248 25044 25276
rect 24995 25245 25007 25248
rect 24949 25239 25007 25245
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 25314 25285 25320 25288
rect 25312 25276 25320 25285
rect 25275 25248 25320 25276
rect 25312 25239 25320 25248
rect 25314 25236 25320 25239
rect 25372 25236 25378 25288
rect 25590 25236 25596 25288
rect 25648 25285 25654 25288
rect 25648 25279 25687 25285
rect 25675 25245 25687 25279
rect 25648 25239 25687 25245
rect 25648 25236 25654 25239
rect 25774 25236 25780 25288
rect 25832 25236 25838 25288
rect 26320 25279 26378 25285
rect 26320 25245 26332 25279
rect 26366 25276 26378 25279
rect 26694 25276 26700 25288
rect 26366 25248 26700 25276
rect 26366 25245 26378 25248
rect 26320 25239 26378 25245
rect 26694 25236 26700 25248
rect 26752 25236 26758 25288
rect 27798 25236 27804 25288
rect 27856 25236 27862 25288
rect 27893 25279 27951 25285
rect 27893 25245 27905 25279
rect 27939 25276 27951 25279
rect 28092 25276 28120 25304
rect 28644 25285 28672 25316
rect 28718 25304 28724 25316
rect 28776 25344 28782 25356
rect 28776 25316 29132 25344
rect 28776 25304 28782 25316
rect 27939 25248 28120 25276
rect 27939 25245 27951 25248
rect 27893 25239 27951 25245
rect 23201 25211 23259 25217
rect 23201 25208 23213 25211
rect 22940 25180 23213 25208
rect 23201 25177 23213 25180
rect 23247 25177 23259 25211
rect 23201 25171 23259 25177
rect 23014 25140 23020 25152
rect 22848 25112 23020 25140
rect 22281 25103 22339 25109
rect 23014 25100 23020 25112
rect 23072 25100 23078 25152
rect 23216 25140 23244 25171
rect 23658 25168 23664 25220
rect 23716 25168 23722 25220
rect 25056 25208 25084 25236
rect 25406 25208 25412 25220
rect 25056 25180 25412 25208
rect 25406 25168 25412 25180
rect 25464 25168 25470 25220
rect 25498 25168 25504 25220
rect 25556 25168 25562 25220
rect 27816 25208 27844 25236
rect 27724 25180 27844 25208
rect 28092 25208 28120 25248
rect 28629 25279 28687 25285
rect 28629 25245 28641 25279
rect 28675 25245 28687 25279
rect 28629 25239 28687 25245
rect 28810 25236 28816 25288
rect 28868 25236 28874 25288
rect 29104 25285 29132 25316
rect 28905 25279 28963 25285
rect 28905 25245 28917 25279
rect 28951 25245 28963 25279
rect 28905 25239 28963 25245
rect 29089 25279 29147 25285
rect 29089 25245 29101 25279
rect 29135 25245 29147 25279
rect 29380 25276 29408 25440
rect 30926 25372 30932 25424
rect 30984 25412 30990 25424
rect 32493 25415 32551 25421
rect 32493 25412 32505 25415
rect 30984 25384 31432 25412
rect 30984 25372 30990 25384
rect 31113 25347 31171 25353
rect 31113 25313 31125 25347
rect 31159 25344 31171 25347
rect 31159 25316 31340 25344
rect 31159 25313 31171 25316
rect 31113 25307 31171 25313
rect 29380 25248 30052 25276
rect 29089 25239 29147 25245
rect 28920 25208 28948 25239
rect 30024 25208 30052 25248
rect 30374 25236 30380 25288
rect 30432 25276 30438 25288
rect 30929 25279 30987 25285
rect 30929 25276 30941 25279
rect 30432 25248 30941 25276
rect 30432 25236 30438 25248
rect 30929 25245 30941 25248
rect 30975 25245 30987 25279
rect 30929 25239 30987 25245
rect 31202 25236 31208 25288
rect 31260 25236 31266 25288
rect 31312 25285 31340 25316
rect 31297 25279 31355 25285
rect 31297 25245 31309 25279
rect 31343 25245 31355 25279
rect 31404 25276 31432 25384
rect 31864 25384 32505 25412
rect 31665 25279 31723 25285
rect 31665 25276 31677 25279
rect 31404 25248 31677 25276
rect 31297 25239 31355 25245
rect 31665 25245 31677 25248
rect 31711 25245 31723 25279
rect 31665 25239 31723 25245
rect 31864 25220 31892 25384
rect 32493 25381 32505 25384
rect 32539 25381 32551 25415
rect 32493 25375 32551 25381
rect 33778 25236 33784 25288
rect 33836 25276 33842 25288
rect 33873 25279 33931 25285
rect 33873 25276 33885 25279
rect 33836 25248 33885 25276
rect 33836 25236 33842 25248
rect 33873 25245 33885 25248
rect 33919 25245 33931 25279
rect 33873 25239 33931 25245
rect 35526 25236 35532 25288
rect 35584 25276 35590 25288
rect 36081 25279 36139 25285
rect 36081 25276 36093 25279
rect 35584 25248 36093 25276
rect 35584 25236 35590 25248
rect 36081 25245 36093 25248
rect 36127 25245 36139 25279
rect 36081 25239 36139 25245
rect 36265 25279 36323 25285
rect 36265 25245 36277 25279
rect 36311 25276 36323 25279
rect 37274 25276 37280 25288
rect 36311 25248 37280 25276
rect 36311 25245 36323 25248
rect 36265 25239 36323 25245
rect 37274 25236 37280 25248
rect 37332 25236 37338 25288
rect 30662 25211 30720 25217
rect 30662 25208 30674 25211
rect 28092 25180 29408 25208
rect 30024 25180 30674 25208
rect 27724 25152 27752 25180
rect 24029 25143 24087 25149
rect 24029 25140 24041 25143
rect 23216 25112 24041 25140
rect 24029 25109 24041 25112
rect 24075 25109 24087 25143
rect 24029 25103 24087 25109
rect 27706 25100 27712 25152
rect 27764 25100 27770 25152
rect 28721 25143 28779 25149
rect 28721 25109 28733 25143
rect 28767 25140 28779 25143
rect 29086 25140 29092 25152
rect 28767 25112 29092 25140
rect 28767 25109 28779 25112
rect 28721 25103 28779 25109
rect 29086 25100 29092 25112
rect 29144 25100 29150 25152
rect 29380 25140 29408 25180
rect 30662 25177 30674 25180
rect 30708 25177 30720 25211
rect 31478 25208 31484 25220
rect 30662 25171 30720 25177
rect 30760 25180 31484 25208
rect 30760 25152 30788 25180
rect 31478 25168 31484 25180
rect 31536 25168 31542 25220
rect 31573 25211 31631 25217
rect 31573 25177 31585 25211
rect 31619 25208 31631 25211
rect 31846 25208 31852 25220
rect 31619 25180 31852 25208
rect 31619 25177 31631 25180
rect 31573 25171 31631 25177
rect 31846 25168 31852 25180
rect 31904 25168 31910 25220
rect 31941 25211 31999 25217
rect 31941 25177 31953 25211
rect 31987 25177 31999 25211
rect 31941 25171 31999 25177
rect 29549 25143 29607 25149
rect 29549 25140 29561 25143
rect 29380 25112 29561 25140
rect 29549 25109 29561 25112
rect 29595 25109 29607 25143
rect 29549 25103 29607 25109
rect 30742 25100 30748 25152
rect 30800 25100 30806 25152
rect 31754 25100 31760 25152
rect 31812 25140 31818 25152
rect 31956 25140 31984 25171
rect 33318 25168 33324 25220
rect 33376 25208 33382 25220
rect 33606 25211 33664 25217
rect 33606 25208 33618 25211
rect 33376 25180 33618 25208
rect 33376 25168 33382 25180
rect 33606 25177 33618 25180
rect 33652 25177 33664 25211
rect 33606 25171 33664 25177
rect 31812 25112 31984 25140
rect 31812 25100 31818 25112
rect 32122 25100 32128 25152
rect 32180 25149 32186 25152
rect 32180 25143 32199 25149
rect 32187 25109 32199 25143
rect 32180 25103 32199 25109
rect 32180 25100 32186 25103
rect 32306 25100 32312 25152
rect 32364 25100 32370 25152
rect 36170 25100 36176 25152
rect 36228 25100 36234 25152
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 11146 24896 11152 24948
rect 11204 24896 11210 24948
rect 11974 24896 11980 24948
rect 12032 24896 12038 24948
rect 12158 24896 12164 24948
rect 12216 24936 12222 24948
rect 12345 24939 12403 24945
rect 12345 24936 12357 24939
rect 12216 24908 12357 24936
rect 12216 24896 12222 24908
rect 12345 24905 12357 24908
rect 12391 24905 12403 24939
rect 12345 24899 12403 24905
rect 13998 24896 14004 24948
rect 14056 24896 14062 24948
rect 15381 24939 15439 24945
rect 15381 24905 15393 24939
rect 15427 24936 15439 24939
rect 16022 24936 16028 24948
rect 15427 24908 16028 24936
rect 15427 24905 15439 24908
rect 15381 24899 15439 24905
rect 16022 24896 16028 24908
rect 16080 24896 16086 24948
rect 16485 24939 16543 24945
rect 16485 24905 16497 24939
rect 16531 24936 16543 24939
rect 16574 24936 16580 24948
rect 16531 24908 16580 24936
rect 16531 24905 16543 24908
rect 16485 24899 16543 24905
rect 16574 24896 16580 24908
rect 16632 24896 16638 24948
rect 16666 24896 16672 24948
rect 16724 24896 16730 24948
rect 19426 24896 19432 24948
rect 19484 24896 19490 24948
rect 19613 24939 19671 24945
rect 19613 24905 19625 24939
rect 19659 24936 19671 24939
rect 19978 24936 19984 24948
rect 19659 24908 19984 24936
rect 19659 24905 19671 24908
rect 19613 24899 19671 24905
rect 19978 24896 19984 24908
rect 20036 24896 20042 24948
rect 22465 24939 22523 24945
rect 22465 24905 22477 24939
rect 22511 24936 22523 24939
rect 22554 24936 22560 24948
rect 22511 24908 22560 24936
rect 22511 24905 22523 24908
rect 22465 24899 22523 24905
rect 22554 24896 22560 24908
rect 22612 24896 22618 24948
rect 22646 24896 22652 24948
rect 22704 24896 22710 24948
rect 23106 24896 23112 24948
rect 23164 24936 23170 24948
rect 24946 24936 24952 24948
rect 23164 24908 24952 24936
rect 23164 24896 23170 24908
rect 9306 24828 9312 24880
rect 9364 24828 9370 24880
rect 11238 24868 11244 24880
rect 10980 24840 11244 24868
rect 10134 24760 10140 24812
rect 10192 24800 10198 24812
rect 10980 24800 11008 24840
rect 11238 24828 11244 24840
rect 11296 24868 11302 24880
rect 11517 24871 11575 24877
rect 11517 24868 11529 24871
rect 11296 24840 11529 24868
rect 11296 24828 11302 24840
rect 11517 24837 11529 24840
rect 11563 24837 11575 24871
rect 11517 24831 11575 24837
rect 11733 24871 11791 24877
rect 11733 24837 11745 24871
rect 11779 24868 11791 24871
rect 12802 24868 12808 24880
rect 11779 24840 12296 24868
rect 11779 24837 11791 24840
rect 11733 24831 11791 24837
rect 10192 24772 11008 24800
rect 11057 24803 11115 24809
rect 10192 24760 10198 24772
rect 11057 24769 11069 24803
rect 11103 24800 11115 24803
rect 11146 24800 11152 24812
rect 11103 24772 11152 24800
rect 11103 24769 11115 24772
rect 11057 24763 11115 24769
rect 11146 24760 11152 24772
rect 11204 24760 11210 24812
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 11900 24772 12173 24800
rect 8297 24735 8355 24741
rect 8297 24701 8309 24735
rect 8343 24701 8355 24735
rect 8297 24695 8355 24701
rect 8573 24735 8631 24741
rect 8573 24701 8585 24735
rect 8619 24732 8631 24735
rect 9858 24732 9864 24744
rect 8619 24704 9864 24732
rect 8619 24701 8631 24704
rect 8573 24695 8631 24701
rect 7926 24556 7932 24608
rect 7984 24596 7990 24608
rect 8312 24596 8340 24695
rect 9858 24692 9864 24704
rect 9916 24692 9922 24744
rect 10045 24735 10103 24741
rect 10045 24701 10057 24735
rect 10091 24732 10103 24735
rect 10413 24735 10471 24741
rect 10413 24732 10425 24735
rect 10091 24704 10425 24732
rect 10091 24701 10103 24704
rect 10045 24695 10103 24701
rect 10413 24701 10425 24704
rect 10459 24732 10471 24735
rect 11514 24732 11520 24744
rect 10459 24704 11520 24732
rect 10459 24701 10471 24704
rect 10413 24695 10471 24701
rect 11514 24692 11520 24704
rect 11572 24692 11578 24744
rect 9582 24624 9588 24676
rect 9640 24624 9646 24676
rect 11900 24673 11928 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 11885 24667 11943 24673
rect 11885 24633 11897 24667
rect 11931 24633 11943 24667
rect 11885 24627 11943 24633
rect 9600 24596 9628 24624
rect 7984 24568 9628 24596
rect 7984 24556 7990 24568
rect 10778 24556 10784 24608
rect 10836 24596 10842 24608
rect 10965 24599 11023 24605
rect 10965 24596 10977 24599
rect 10836 24568 10977 24596
rect 10836 24556 10842 24568
rect 10965 24565 10977 24568
rect 11011 24565 11023 24599
rect 10965 24559 11023 24565
rect 11701 24599 11759 24605
rect 11701 24565 11713 24599
rect 11747 24596 11759 24599
rect 11974 24596 11980 24608
rect 11747 24568 11980 24596
rect 11747 24565 11759 24568
rect 11701 24559 11759 24565
rect 11974 24556 11980 24568
rect 12032 24556 12038 24608
rect 12268 24596 12296 24840
rect 12452 24840 12808 24868
rect 12452 24809 12480 24840
rect 12802 24828 12808 24840
rect 12860 24828 12866 24880
rect 14016 24868 14044 24896
rect 13740 24840 14044 24868
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24769 12495 24803
rect 12437 24763 12495 24769
rect 13081 24803 13139 24809
rect 13081 24769 13093 24803
rect 13127 24800 13139 24803
rect 13740 24800 13768 24840
rect 13127 24772 13768 24800
rect 13127 24769 13139 24772
rect 13081 24763 13139 24769
rect 13814 24760 13820 24812
rect 13872 24800 13878 24812
rect 14274 24809 14280 24812
rect 14001 24803 14059 24809
rect 14001 24800 14013 24803
rect 13872 24772 14013 24800
rect 13872 24760 13878 24772
rect 14001 24769 14013 24772
rect 14047 24769 14059 24803
rect 14001 24763 14059 24769
rect 14268 24763 14280 24809
rect 14274 24760 14280 24763
rect 14332 24760 14338 24812
rect 16298 24760 16304 24812
rect 16356 24760 16362 24812
rect 16684 24809 16712 24896
rect 22281 24871 22339 24877
rect 22281 24837 22293 24871
rect 22327 24868 22339 24871
rect 22664 24868 22692 24896
rect 23216 24877 23244 24908
rect 24946 24896 24952 24908
rect 25004 24896 25010 24948
rect 25406 24896 25412 24948
rect 25464 24896 25470 24948
rect 25498 24896 25504 24948
rect 25556 24936 25562 24948
rect 25685 24939 25743 24945
rect 25685 24936 25697 24939
rect 25556 24908 25697 24936
rect 25556 24896 25562 24908
rect 25685 24905 25697 24908
rect 25731 24905 25743 24939
rect 25685 24899 25743 24905
rect 29086 24896 29092 24948
rect 29144 24936 29150 24948
rect 29523 24939 29581 24945
rect 29523 24936 29535 24939
rect 29144 24908 29535 24936
rect 29144 24896 29150 24908
rect 29523 24905 29535 24908
rect 29569 24905 29581 24939
rect 29523 24899 29581 24905
rect 30742 24896 30748 24948
rect 30800 24936 30806 24948
rect 30929 24939 30987 24945
rect 30929 24936 30941 24939
rect 30800 24908 30941 24936
rect 30800 24896 30806 24908
rect 30929 24905 30941 24908
rect 30975 24905 30987 24939
rect 30929 24899 30987 24905
rect 31202 24896 31208 24948
rect 31260 24936 31266 24948
rect 32214 24936 32220 24948
rect 31260 24908 32220 24936
rect 31260 24896 31266 24908
rect 32214 24896 32220 24908
rect 32272 24896 32278 24948
rect 32306 24896 32312 24948
rect 32364 24896 32370 24948
rect 33045 24939 33103 24945
rect 33045 24905 33057 24939
rect 33091 24936 33103 24939
rect 33318 24936 33324 24948
rect 33091 24908 33324 24936
rect 33091 24905 33103 24908
rect 33045 24899 33103 24905
rect 33318 24896 33324 24908
rect 33376 24896 33382 24948
rect 22327 24840 22692 24868
rect 23201 24871 23259 24877
rect 22327 24837 22339 24840
rect 22281 24831 22339 24837
rect 23201 24837 23213 24871
rect 23247 24837 23259 24871
rect 23201 24831 23259 24837
rect 23431 24837 23489 24843
rect 23431 24834 23443 24837
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 16758 24760 16764 24812
rect 16816 24800 16822 24812
rect 16925 24803 16983 24809
rect 16925 24800 16937 24803
rect 16816 24772 16937 24800
rect 16816 24760 16822 24772
rect 16925 24769 16937 24772
rect 16971 24769 16983 24803
rect 16925 24763 16983 24769
rect 18046 24760 18052 24812
rect 18104 24800 18110 24812
rect 18693 24803 18751 24809
rect 18693 24800 18705 24803
rect 18104 24772 18705 24800
rect 18104 24760 18110 24772
rect 18693 24769 18705 24772
rect 18739 24769 18751 24803
rect 18693 24763 18751 24769
rect 19242 24760 19248 24812
rect 19300 24760 19306 24812
rect 19521 24803 19579 24809
rect 19521 24769 19533 24803
rect 19567 24800 19579 24803
rect 19567 24772 20208 24800
rect 19567 24769 19579 24772
rect 19521 24763 19579 24769
rect 20180 24744 20208 24772
rect 20806 24760 20812 24812
rect 20864 24800 20870 24812
rect 21453 24803 21511 24809
rect 21453 24800 21465 24803
rect 20864 24772 21465 24800
rect 20864 24760 20870 24772
rect 21453 24769 21465 24772
rect 21499 24800 21511 24803
rect 21542 24800 21548 24812
rect 21499 24772 21548 24800
rect 21499 24769 21511 24772
rect 21453 24763 21511 24769
rect 21542 24760 21548 24772
rect 21600 24760 21606 24812
rect 21726 24760 21732 24812
rect 21784 24800 21790 24812
rect 22005 24803 22063 24809
rect 22005 24800 22017 24803
rect 21784 24772 22017 24800
rect 21784 24760 21790 24772
rect 22005 24769 22017 24772
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 22152 24772 22201 24800
rect 22152 24760 22158 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24701 13323 24735
rect 13265 24695 13323 24701
rect 12618 24596 12624 24608
rect 12268 24568 12624 24596
rect 12618 24556 12624 24568
rect 12676 24556 12682 24608
rect 12894 24556 12900 24608
rect 12952 24556 12958 24608
rect 13280 24596 13308 24695
rect 20162 24692 20168 24744
rect 20220 24692 20226 24744
rect 20530 24692 20536 24744
rect 20588 24692 20594 24744
rect 22204 24732 22232 24763
rect 22370 24760 22376 24812
rect 22428 24800 22434 24812
rect 23416 24803 23443 24834
rect 23477 24803 23489 24837
rect 23566 24828 23572 24880
rect 23624 24868 23630 24880
rect 23937 24871 23995 24877
rect 23937 24868 23949 24871
rect 23624 24840 23949 24868
rect 23624 24828 23630 24840
rect 23937 24837 23949 24840
rect 23983 24837 23995 24871
rect 23937 24831 23995 24837
rect 24578 24828 24584 24880
rect 24636 24828 24642 24880
rect 23416 24800 23489 24803
rect 22428 24797 23489 24800
rect 25424 24800 25452 24896
rect 29733 24871 29791 24877
rect 29733 24868 29745 24871
rect 28276 24840 29745 24868
rect 25593 24803 25651 24809
rect 25593 24800 25605 24803
rect 22428 24772 23444 24797
rect 25424 24772 25605 24800
rect 22428 24760 22434 24772
rect 25593 24769 25605 24772
rect 25639 24769 25651 24803
rect 25593 24763 25651 24769
rect 25774 24760 25780 24812
rect 25832 24760 25838 24812
rect 27614 24760 27620 24812
rect 27672 24760 27678 24812
rect 28074 24760 28080 24812
rect 28132 24800 28138 24812
rect 28276 24809 28304 24840
rect 29733 24837 29745 24840
rect 29779 24837 29791 24871
rect 29733 24831 29791 24837
rect 31846 24828 31852 24880
rect 31904 24868 31910 24880
rect 31941 24871 31999 24877
rect 31941 24868 31953 24871
rect 31904 24840 31953 24868
rect 31904 24828 31910 24840
rect 31941 24837 31953 24840
rect 31987 24837 31999 24871
rect 32324 24868 32352 24896
rect 35980 24871 36038 24877
rect 32324 24840 32904 24868
rect 31941 24831 31999 24837
rect 28261 24803 28319 24809
rect 28261 24800 28273 24803
rect 28132 24772 28273 24800
rect 28132 24760 28138 24772
rect 28261 24769 28273 24772
rect 28307 24769 28319 24803
rect 28261 24763 28319 24769
rect 28445 24803 28503 24809
rect 28445 24769 28457 24803
rect 28491 24800 28503 24803
rect 28718 24800 28724 24812
rect 28491 24772 28724 24800
rect 28491 24769 28503 24772
rect 28445 24763 28503 24769
rect 28718 24760 28724 24772
rect 28776 24760 28782 24812
rect 30650 24760 30656 24812
rect 30708 24800 30714 24812
rect 30837 24803 30895 24809
rect 30837 24800 30849 24803
rect 30708 24772 30849 24800
rect 30708 24760 30714 24772
rect 30837 24769 30849 24772
rect 30883 24769 30895 24803
rect 30837 24763 30895 24769
rect 30926 24760 30932 24812
rect 30984 24800 30990 24812
rect 31021 24803 31079 24809
rect 31021 24800 31033 24803
rect 30984 24772 31033 24800
rect 30984 24760 30990 24772
rect 31021 24769 31033 24772
rect 31067 24769 31079 24803
rect 31021 24763 31079 24769
rect 31481 24803 31539 24809
rect 31481 24769 31493 24803
rect 31527 24769 31539 24803
rect 31481 24763 31539 24769
rect 31665 24803 31723 24809
rect 31665 24769 31677 24803
rect 31711 24800 31723 24803
rect 32214 24800 32220 24812
rect 31711 24772 32220 24800
rect 31711 24769 31723 24772
rect 31665 24763 31723 24769
rect 23017 24735 23075 24741
rect 23017 24732 23029 24735
rect 22204 24704 23029 24732
rect 23017 24701 23029 24704
rect 23063 24701 23075 24735
rect 23017 24695 23075 24701
rect 23661 24735 23719 24741
rect 23661 24701 23673 24735
rect 23707 24701 23719 24735
rect 27632 24732 27660 24760
rect 28166 24732 28172 24744
rect 27632 24704 28172 24732
rect 23661 24695 23719 24701
rect 15746 24624 15752 24676
rect 15804 24624 15810 24676
rect 18690 24664 18696 24676
rect 18064 24636 18696 24664
rect 15764 24596 15792 24624
rect 13280 24568 15792 24596
rect 16666 24556 16672 24608
rect 16724 24596 16730 24608
rect 18064 24605 18092 24636
rect 18690 24624 18696 24636
rect 18748 24624 18754 24676
rect 23566 24624 23572 24676
rect 23624 24624 23630 24676
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 16724 24568 18061 24596
rect 16724 24556 16730 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 18138 24556 18144 24608
rect 18196 24556 18202 24608
rect 19886 24556 19892 24608
rect 19944 24556 19950 24608
rect 20714 24556 20720 24608
rect 20772 24596 20778 24608
rect 20901 24599 20959 24605
rect 20901 24596 20913 24599
rect 20772 24568 20913 24596
rect 20772 24556 20778 24568
rect 20901 24565 20913 24568
rect 20947 24565 20959 24599
rect 20901 24559 20959 24565
rect 21910 24556 21916 24608
rect 21968 24556 21974 24608
rect 23290 24556 23296 24608
rect 23348 24596 23354 24608
rect 23385 24599 23443 24605
rect 23385 24596 23397 24599
rect 23348 24568 23397 24596
rect 23348 24556 23354 24568
rect 23385 24565 23397 24568
rect 23431 24565 23443 24599
rect 23676 24596 23704 24695
rect 28166 24692 28172 24704
rect 28224 24732 28230 24744
rect 28537 24735 28595 24741
rect 28537 24732 28549 24735
rect 28224 24704 28549 24732
rect 28224 24692 28230 24704
rect 28537 24701 28549 24704
rect 28583 24701 28595 24735
rect 28537 24695 28595 24701
rect 31110 24692 31116 24744
rect 31168 24732 31174 24744
rect 31168 24704 31340 24732
rect 31168 24692 31174 24704
rect 29178 24624 29184 24676
rect 29236 24664 29242 24676
rect 31312 24673 31340 24704
rect 29365 24667 29423 24673
rect 29365 24664 29377 24667
rect 29236 24636 29377 24664
rect 29236 24624 29242 24636
rect 29365 24633 29377 24636
rect 29411 24633 29423 24667
rect 29365 24627 29423 24633
rect 31297 24667 31355 24673
rect 31297 24633 31309 24667
rect 31343 24633 31355 24667
rect 31496 24664 31524 24763
rect 32214 24760 32220 24772
rect 32272 24800 32278 24812
rect 32401 24803 32459 24809
rect 32401 24800 32413 24803
rect 32272 24772 32413 24800
rect 32272 24760 32278 24772
rect 32401 24769 32413 24772
rect 32447 24769 32459 24803
rect 32401 24763 32459 24769
rect 32490 24760 32496 24812
rect 32548 24760 32554 24812
rect 32582 24760 32588 24812
rect 32640 24760 32646 24812
rect 32876 24809 32904 24840
rect 34348 24840 34652 24868
rect 34348 24812 34376 24840
rect 32861 24803 32919 24809
rect 32861 24769 32873 24803
rect 32907 24769 32919 24803
rect 32861 24763 32919 24769
rect 33778 24760 33784 24812
rect 33836 24800 33842 24812
rect 34241 24803 34299 24809
rect 34241 24800 34253 24803
rect 33836 24772 34253 24800
rect 33836 24760 33842 24772
rect 34241 24769 34253 24772
rect 34287 24800 34299 24803
rect 34330 24800 34336 24812
rect 34287 24772 34336 24800
rect 34287 24769 34299 24772
rect 34241 24763 34299 24769
rect 34330 24760 34336 24772
rect 34388 24760 34394 24812
rect 34514 24809 34520 24812
rect 34508 24763 34520 24809
rect 34514 24760 34520 24763
rect 34572 24760 34578 24812
rect 34624 24800 34652 24840
rect 35980 24837 35992 24871
rect 36026 24868 36038 24871
rect 36170 24868 36176 24880
rect 36026 24840 36176 24868
rect 36026 24837 36038 24840
rect 35980 24831 36038 24837
rect 36170 24828 36176 24840
rect 36228 24828 36234 24880
rect 35713 24803 35771 24809
rect 35713 24800 35725 24803
rect 34624 24772 35725 24800
rect 35713 24769 35725 24772
rect 35759 24769 35771 24803
rect 35713 24763 35771 24769
rect 31846 24692 31852 24744
rect 31904 24732 31910 24744
rect 32769 24735 32827 24741
rect 32769 24732 32781 24735
rect 31904 24704 32781 24732
rect 31904 24692 31910 24704
rect 32769 24701 32781 24704
rect 32815 24701 32827 24735
rect 37277 24735 37335 24741
rect 37277 24732 37289 24735
rect 32769 24695 32827 24701
rect 37108 24704 37289 24732
rect 32582 24664 32588 24676
rect 31496 24636 32588 24664
rect 31297 24627 31355 24633
rect 32582 24624 32588 24636
rect 32640 24624 32646 24676
rect 37108 24673 37136 24704
rect 37277 24701 37289 24704
rect 37323 24701 37335 24735
rect 37277 24695 37335 24701
rect 37093 24667 37151 24673
rect 37093 24633 37105 24667
rect 37139 24633 37151 24667
rect 37093 24627 37151 24633
rect 24670 24596 24676 24608
rect 23676 24568 24676 24596
rect 23385 24559 23443 24565
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 28074 24556 28080 24608
rect 28132 24556 28138 24608
rect 29546 24556 29552 24608
rect 29604 24596 29610 24608
rect 31754 24596 31760 24608
rect 29604 24568 31760 24596
rect 29604 24556 29610 24568
rect 31754 24556 31760 24568
rect 31812 24556 31818 24608
rect 31849 24599 31907 24605
rect 31849 24565 31861 24599
rect 31895 24596 31907 24599
rect 32490 24596 32496 24608
rect 31895 24568 32496 24596
rect 31895 24565 31907 24568
rect 31849 24559 31907 24565
rect 32490 24556 32496 24568
rect 32548 24556 32554 24608
rect 35621 24599 35679 24605
rect 35621 24565 35633 24599
rect 35667 24596 35679 24599
rect 35986 24596 35992 24608
rect 35667 24568 35992 24596
rect 35667 24565 35679 24568
rect 35621 24559 35679 24565
rect 35986 24556 35992 24568
rect 36044 24556 36050 24608
rect 36078 24556 36084 24608
rect 36136 24596 36142 24608
rect 37108 24596 37136 24627
rect 36136 24568 37136 24596
rect 36136 24556 36142 24568
rect 37918 24556 37924 24608
rect 37976 24556 37982 24608
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 9306 24352 9312 24404
rect 9364 24392 9370 24404
rect 9401 24395 9459 24401
rect 9401 24392 9413 24395
rect 9364 24364 9413 24392
rect 9364 24352 9370 24364
rect 9401 24361 9413 24364
rect 9447 24361 9459 24395
rect 9401 24355 9459 24361
rect 9858 24352 9864 24404
rect 9916 24392 9922 24404
rect 10689 24395 10747 24401
rect 10689 24392 10701 24395
rect 9916 24364 10701 24392
rect 9916 24352 9922 24364
rect 10689 24361 10701 24364
rect 10735 24361 10747 24395
rect 10689 24355 10747 24361
rect 12621 24395 12679 24401
rect 12621 24361 12633 24395
rect 12667 24392 12679 24395
rect 12802 24392 12808 24404
rect 12667 24364 12808 24392
rect 12667 24361 12679 24364
rect 12621 24355 12679 24361
rect 12802 24352 12808 24364
rect 12860 24352 12866 24404
rect 12894 24352 12900 24404
rect 12952 24352 12958 24404
rect 13173 24395 13231 24401
rect 13173 24361 13185 24395
rect 13219 24392 13231 24395
rect 13998 24392 14004 24404
rect 13219 24364 14004 24392
rect 13219 24361 13231 24364
rect 13173 24355 13231 24361
rect 13998 24352 14004 24364
rect 14056 24352 14062 24404
rect 14274 24352 14280 24404
rect 14332 24392 14338 24404
rect 14461 24395 14519 24401
rect 14461 24392 14473 24395
rect 14332 24364 14473 24392
rect 14332 24352 14338 24364
rect 14461 24361 14473 24364
rect 14507 24361 14519 24395
rect 14461 24355 14519 24361
rect 16485 24395 16543 24401
rect 16485 24361 16497 24395
rect 16531 24392 16543 24395
rect 16758 24392 16764 24404
rect 16531 24364 16764 24392
rect 16531 24361 16543 24364
rect 16485 24355 16543 24361
rect 16758 24352 16764 24364
rect 16816 24352 16822 24404
rect 18138 24352 18144 24404
rect 18196 24352 18202 24404
rect 19242 24352 19248 24404
rect 19300 24392 19306 24404
rect 19613 24395 19671 24401
rect 19613 24392 19625 24395
rect 19300 24364 19625 24392
rect 19300 24352 19306 24364
rect 19613 24361 19625 24364
rect 19659 24361 19671 24395
rect 20806 24392 20812 24404
rect 19613 24355 19671 24361
rect 20272 24364 20812 24392
rect 10318 24284 10324 24336
rect 10376 24324 10382 24336
rect 10376 24296 11652 24324
rect 10376 24284 10382 24296
rect 9309 24191 9367 24197
rect 9309 24188 9321 24191
rect 8864 24160 9321 24188
rect 8864 24064 8892 24160
rect 9309 24157 9321 24160
rect 9355 24188 9367 24191
rect 9355 24160 9674 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9646 24120 9674 24160
rect 9950 24148 9956 24200
rect 10008 24148 10014 24200
rect 10502 24148 10508 24200
rect 10560 24188 10566 24200
rect 10873 24191 10931 24197
rect 10873 24188 10885 24191
rect 10560 24160 10885 24188
rect 10560 24148 10566 24160
rect 10873 24157 10885 24160
rect 10919 24157 10931 24191
rect 10873 24151 10931 24157
rect 10965 24191 11023 24197
rect 10965 24157 10977 24191
rect 11011 24157 11023 24191
rect 10965 24151 11023 24157
rect 9646 24092 10732 24120
rect 8846 24012 8852 24064
rect 8904 24012 8910 24064
rect 10594 24012 10600 24064
rect 10652 24012 10658 24064
rect 10704 24052 10732 24092
rect 10778 24080 10784 24132
rect 10836 24120 10842 24132
rect 10980 24120 11008 24151
rect 11238 24148 11244 24200
rect 11296 24148 11302 24200
rect 11330 24148 11336 24200
rect 11388 24148 11394 24200
rect 11514 24148 11520 24200
rect 11572 24148 11578 24200
rect 10836 24092 11008 24120
rect 11057 24123 11115 24129
rect 10836 24080 10842 24092
rect 11057 24089 11069 24123
rect 11103 24120 11115 24123
rect 11425 24123 11483 24129
rect 11425 24120 11437 24123
rect 11103 24092 11437 24120
rect 11103 24089 11115 24092
rect 11057 24083 11115 24089
rect 11425 24089 11437 24092
rect 11471 24089 11483 24123
rect 11624 24120 11652 24296
rect 12618 24256 12624 24268
rect 12176 24228 12624 24256
rect 12176 24197 12204 24228
rect 12618 24216 12624 24228
rect 12676 24216 12682 24268
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24157 12219 24191
rect 12161 24151 12219 24157
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24188 12495 24191
rect 12912 24188 12940 24352
rect 16853 24327 16911 24333
rect 16853 24293 16865 24327
rect 16899 24324 16911 24327
rect 18156 24324 18184 24352
rect 16899 24296 17540 24324
rect 16899 24293 16911 24296
rect 16853 24287 16911 24293
rect 15473 24259 15531 24265
rect 15473 24256 15485 24259
rect 14476 24228 15485 24256
rect 12483 24160 12940 24188
rect 12483 24157 12495 24160
rect 12437 24151 12495 24157
rect 12452 24120 12480 24151
rect 13078 24148 13084 24200
rect 13136 24148 13142 24200
rect 14476 24197 14504 24228
rect 15473 24225 15485 24228
rect 15519 24225 15531 24259
rect 15473 24219 15531 24225
rect 15746 24216 15752 24268
rect 15804 24216 15810 24268
rect 17512 24265 17540 24296
rect 17604 24296 18184 24324
rect 16945 24259 17003 24265
rect 16945 24256 16957 24259
rect 16500 24228 16957 24256
rect 13265 24191 13323 24197
rect 13265 24188 13277 24191
rect 13188 24160 13277 24188
rect 12713 24123 12771 24129
rect 12713 24120 12725 24123
rect 11624 24092 12480 24120
rect 12544 24092 12725 24120
rect 11425 24083 11483 24089
rect 11146 24052 11152 24064
rect 10704 24024 11152 24052
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 11238 24012 11244 24064
rect 11296 24052 11302 24064
rect 12253 24055 12311 24061
rect 12253 24052 12265 24055
rect 11296 24024 12265 24052
rect 11296 24012 11302 24024
rect 12253 24021 12265 24024
rect 12299 24052 12311 24055
rect 12544 24052 12572 24092
rect 12713 24089 12725 24092
rect 12759 24089 12771 24123
rect 12713 24083 12771 24089
rect 12894 24080 12900 24132
rect 12952 24080 12958 24132
rect 13188 24064 13216 24160
rect 13265 24157 13277 24160
rect 13311 24157 13323 24191
rect 13265 24151 13323 24157
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14645 24191 14703 24197
rect 14645 24157 14657 24191
rect 14691 24157 14703 24191
rect 14645 24151 14703 24157
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24188 15439 24191
rect 15764 24188 15792 24216
rect 15427 24160 15792 24188
rect 15427 24157 15439 24160
rect 15381 24151 15439 24157
rect 14660 24120 14688 24151
rect 15930 24148 15936 24200
rect 15988 24188 15994 24200
rect 16500 24197 16528 24228
rect 16945 24225 16957 24228
rect 16991 24225 17003 24259
rect 16945 24219 17003 24225
rect 17497 24259 17555 24265
rect 17497 24225 17509 24259
rect 17543 24225 17555 24259
rect 17497 24219 17555 24225
rect 16025 24191 16083 24197
rect 16025 24188 16037 24191
rect 15988 24160 16037 24188
rect 15988 24148 15994 24160
rect 16025 24157 16037 24160
rect 16071 24157 16083 24191
rect 16025 24151 16083 24157
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24157 16359 24191
rect 16301 24151 16359 24157
rect 16485 24191 16543 24197
rect 16485 24157 16497 24191
rect 16531 24157 16543 24191
rect 16485 24151 16543 24157
rect 16316 24120 16344 24151
rect 16574 24148 16580 24200
rect 16632 24148 16638 24200
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 17604 24188 17632 24296
rect 19058 24216 19064 24268
rect 19116 24216 19122 24268
rect 20272 24265 20300 24364
rect 20806 24352 20812 24364
rect 20864 24352 20870 24404
rect 22373 24395 22431 24401
rect 22373 24361 22385 24395
rect 22419 24361 22431 24395
rect 22373 24355 22431 24361
rect 21910 24284 21916 24336
rect 21968 24284 21974 24336
rect 22186 24284 22192 24336
rect 22244 24324 22250 24336
rect 22388 24324 22416 24355
rect 24578 24352 24584 24404
rect 24636 24392 24642 24404
rect 24673 24395 24731 24401
rect 24673 24392 24685 24395
rect 24636 24364 24685 24392
rect 24636 24352 24642 24364
rect 24673 24361 24685 24364
rect 24719 24361 24731 24395
rect 24673 24355 24731 24361
rect 30558 24352 30564 24404
rect 30616 24352 30622 24404
rect 30745 24395 30803 24401
rect 30745 24361 30757 24395
rect 30791 24392 30803 24395
rect 30926 24392 30932 24404
rect 30791 24364 30932 24392
rect 30791 24361 30803 24364
rect 30745 24355 30803 24361
rect 30926 24352 30932 24364
rect 30984 24352 30990 24404
rect 32122 24352 32128 24404
rect 32180 24392 32186 24404
rect 32401 24395 32459 24401
rect 32401 24392 32413 24395
rect 32180 24364 32413 24392
rect 32180 24352 32186 24364
rect 32401 24361 32413 24364
rect 32447 24361 32459 24395
rect 33134 24392 33140 24404
rect 32401 24355 32459 24361
rect 32692 24364 33140 24392
rect 22244 24296 22416 24324
rect 22244 24284 22250 24296
rect 29914 24284 29920 24336
rect 29972 24324 29978 24336
rect 32692 24324 32720 24364
rect 33134 24352 33140 24364
rect 33192 24392 33198 24404
rect 33192 24364 34468 24392
rect 33192 24352 33198 24364
rect 29972 24296 32720 24324
rect 34440 24324 34468 24364
rect 34514 24352 34520 24404
rect 34572 24392 34578 24404
rect 34977 24395 35035 24401
rect 34977 24392 34989 24395
rect 34572 24364 34989 24392
rect 34572 24352 34578 24364
rect 34977 24361 34989 24364
rect 35023 24361 35035 24395
rect 34977 24355 35035 24361
rect 37274 24352 37280 24404
rect 37332 24352 37338 24404
rect 37918 24352 37924 24404
rect 37976 24352 37982 24404
rect 34440 24296 37228 24324
rect 29972 24284 29978 24296
rect 20257 24259 20315 24265
rect 20257 24225 20269 24259
rect 20303 24225 20315 24259
rect 20257 24219 20315 24225
rect 20717 24259 20775 24265
rect 20717 24225 20729 24259
rect 20763 24256 20775 24259
rect 21450 24256 21456 24268
rect 20763 24228 21456 24256
rect 20763 24225 20775 24228
rect 20717 24219 20775 24225
rect 21450 24216 21456 24228
rect 21508 24216 21514 24268
rect 16899 24160 17632 24188
rect 19076 24188 19104 24216
rect 20441 24191 20499 24197
rect 20441 24188 20453 24191
rect 19076 24160 20453 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 20441 24157 20453 24160
rect 20487 24157 20499 24191
rect 21928 24188 21956 24284
rect 27433 24259 27491 24265
rect 21850 24160 21956 24188
rect 22066 24228 24624 24256
rect 20441 24151 20499 24157
rect 14660 24092 16344 24120
rect 16592 24120 16620 24148
rect 17494 24120 17500 24132
rect 16592 24092 17500 24120
rect 15396 24064 15424 24092
rect 17494 24080 17500 24092
rect 17552 24080 17558 24132
rect 18506 24080 18512 24132
rect 18564 24120 18570 24132
rect 18794 24123 18852 24129
rect 18794 24120 18806 24123
rect 18564 24092 18806 24120
rect 18564 24080 18570 24092
rect 18794 24089 18806 24092
rect 18840 24089 18852 24123
rect 18794 24083 18852 24089
rect 19886 24080 19892 24132
rect 19944 24120 19950 24132
rect 19981 24123 20039 24129
rect 19981 24120 19993 24123
rect 19944 24092 19993 24120
rect 19944 24080 19950 24092
rect 19981 24089 19993 24092
rect 20027 24089 20039 24123
rect 19981 24083 20039 24089
rect 12299 24024 12572 24052
rect 12299 24021 12311 24024
rect 12253 24015 12311 24021
rect 13170 24012 13176 24064
rect 13228 24012 13234 24064
rect 14734 24012 14740 24064
rect 14792 24012 14798 24064
rect 15378 24012 15384 24064
rect 15436 24012 15442 24064
rect 16666 24012 16672 24064
rect 16724 24012 16730 24064
rect 17218 24012 17224 24064
rect 17276 24052 17282 24064
rect 17681 24055 17739 24061
rect 17681 24052 17693 24055
rect 17276 24024 17693 24052
rect 17276 24012 17282 24024
rect 17681 24021 17693 24024
rect 17727 24021 17739 24055
rect 17681 24015 17739 24021
rect 20070 24012 20076 24064
rect 20128 24012 20134 24064
rect 21726 24012 21732 24064
rect 21784 24052 21790 24064
rect 22066 24052 22094 24228
rect 22186 24148 22192 24200
rect 22244 24148 22250 24200
rect 22646 24148 22652 24200
rect 22704 24148 22710 24200
rect 24596 24197 24624 24228
rect 27433 24225 27445 24259
rect 27479 24256 27491 24259
rect 27614 24256 27620 24268
rect 27479 24228 27620 24256
rect 27479 24225 27491 24228
rect 27433 24219 27491 24225
rect 27614 24216 27620 24228
rect 27672 24256 27678 24268
rect 28074 24256 28080 24268
rect 27672 24228 28080 24256
rect 27672 24216 27678 24228
rect 28074 24216 28080 24228
rect 28132 24216 28138 24268
rect 29270 24216 29276 24268
rect 29328 24216 29334 24268
rect 31846 24216 31852 24268
rect 31904 24256 31910 24268
rect 31941 24259 31999 24265
rect 31941 24256 31953 24259
rect 31904 24228 31953 24256
rect 31904 24216 31910 24228
rect 31941 24225 31953 24228
rect 31987 24225 31999 24259
rect 31941 24219 31999 24225
rect 32125 24259 32183 24265
rect 32125 24225 32137 24259
rect 32171 24256 32183 24259
rect 32490 24256 32496 24268
rect 32171 24228 32496 24256
rect 32171 24225 32183 24228
rect 32125 24219 32183 24225
rect 22741 24191 22799 24197
rect 22741 24157 22753 24191
rect 22787 24157 22799 24191
rect 22741 24151 22799 24157
rect 24581 24191 24639 24197
rect 24581 24157 24593 24191
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 25409 24191 25467 24197
rect 25409 24157 25421 24191
rect 25455 24188 25467 24191
rect 25682 24188 25688 24200
rect 25455 24160 25688 24188
rect 25455 24157 25467 24160
rect 25409 24151 25467 24157
rect 22204 24061 22232 24148
rect 22278 24080 22284 24132
rect 22336 24080 22342 24132
rect 21784 24024 22094 24052
rect 22189 24055 22247 24061
rect 21784 24012 21790 24024
rect 22189 24021 22201 24055
rect 22235 24052 22247 24055
rect 22756 24052 22784 24151
rect 25682 24148 25688 24160
rect 25740 24148 25746 24200
rect 27338 24148 27344 24200
rect 27396 24148 27402 24200
rect 27982 24148 27988 24200
rect 28040 24188 28046 24200
rect 28040 24160 28120 24188
rect 28040 24148 28046 24160
rect 28092 24129 28120 24160
rect 28166 24148 28172 24200
rect 28224 24188 28230 24200
rect 28261 24191 28319 24197
rect 28261 24188 28273 24191
rect 28224 24160 28273 24188
rect 28224 24148 28230 24160
rect 28261 24157 28273 24160
rect 28307 24157 28319 24191
rect 28261 24151 28319 24157
rect 28350 24148 28356 24200
rect 28408 24148 28414 24200
rect 29288 24188 29316 24216
rect 32324 24200 32352 24228
rect 32490 24216 32496 24228
rect 32548 24216 32554 24268
rect 32692 24265 32720 24296
rect 37200 24265 37228 24296
rect 32677 24259 32735 24265
rect 32677 24225 32689 24259
rect 32723 24225 32735 24259
rect 32677 24219 32735 24225
rect 37185 24259 37243 24265
rect 37185 24225 37197 24259
rect 37231 24225 37243 24259
rect 37185 24219 37243 24225
rect 30190 24188 30196 24200
rect 29288 24160 30196 24188
rect 30190 24148 30196 24160
rect 30248 24188 30254 24200
rect 30285 24191 30343 24197
rect 30285 24188 30297 24191
rect 30248 24160 30297 24188
rect 30248 24148 30254 24160
rect 30285 24157 30297 24160
rect 30331 24157 30343 24191
rect 30285 24151 30343 24157
rect 32033 24191 32091 24197
rect 32033 24157 32045 24191
rect 32079 24157 32091 24191
rect 32033 24151 32091 24157
rect 28077 24123 28135 24129
rect 28077 24089 28089 24123
rect 28123 24089 28135 24123
rect 32048 24120 32076 24151
rect 32214 24148 32220 24200
rect 32272 24148 32278 24200
rect 32306 24148 32312 24200
rect 32364 24148 32370 24200
rect 32858 24148 32864 24200
rect 32916 24148 32922 24200
rect 32950 24148 32956 24200
rect 33008 24148 33014 24200
rect 34330 24148 34336 24200
rect 34388 24188 34394 24200
rect 34425 24191 34483 24197
rect 34425 24188 34437 24191
rect 34388 24160 34437 24188
rect 34388 24148 34394 24160
rect 34425 24157 34437 24160
rect 34471 24157 34483 24191
rect 34425 24151 34483 24157
rect 35158 24148 35164 24200
rect 35216 24148 35222 24200
rect 35437 24191 35495 24197
rect 35437 24157 35449 24191
rect 35483 24188 35495 24191
rect 35526 24188 35532 24200
rect 35483 24160 35532 24188
rect 35483 24157 35495 24160
rect 35437 24151 35495 24157
rect 35526 24148 35532 24160
rect 35584 24148 35590 24200
rect 35621 24191 35679 24197
rect 35621 24157 35633 24191
rect 35667 24188 35679 24191
rect 35713 24191 35771 24197
rect 35713 24188 35725 24191
rect 35667 24160 35725 24188
rect 35667 24157 35679 24160
rect 35621 24151 35679 24157
rect 35713 24157 35725 24160
rect 35759 24157 35771 24191
rect 35713 24151 35771 24157
rect 35986 24148 35992 24200
rect 36044 24188 36050 24200
rect 36354 24188 36360 24200
rect 36044 24160 36360 24188
rect 36044 24148 36050 24160
rect 36354 24148 36360 24160
rect 36412 24188 36418 24200
rect 37001 24191 37059 24197
rect 37001 24188 37013 24191
rect 36412 24160 37013 24188
rect 36412 24148 36418 24160
rect 37001 24157 37013 24160
rect 37047 24157 37059 24191
rect 37001 24151 37059 24157
rect 37090 24148 37096 24200
rect 37148 24188 37154 24200
rect 37369 24191 37427 24197
rect 37369 24188 37381 24191
rect 37148 24160 37381 24188
rect 37148 24148 37154 24160
rect 37369 24157 37381 24160
rect 37415 24157 37427 24191
rect 37369 24151 37427 24157
rect 37461 24191 37519 24197
rect 37461 24157 37473 24191
rect 37507 24188 37519 24191
rect 37936 24188 37964 24352
rect 37507 24160 37964 24188
rect 37507 24157 37519 24160
rect 37461 24151 37519 24157
rect 32582 24120 32588 24132
rect 32048 24092 32588 24120
rect 28077 24083 28135 24089
rect 32582 24080 32588 24092
rect 32640 24120 32646 24132
rect 32640 24092 33088 24120
rect 32640 24080 32646 24092
rect 33060 24064 33088 24092
rect 34054 24080 34060 24132
rect 34112 24120 34118 24132
rect 34158 24123 34216 24129
rect 34158 24120 34170 24123
rect 34112 24092 34170 24120
rect 34112 24080 34118 24092
rect 34158 24089 34170 24092
rect 34204 24089 34216 24123
rect 34158 24083 34216 24089
rect 22235 24024 22784 24052
rect 22235 24021 22247 24024
rect 22189 24015 22247 24021
rect 22922 24012 22928 24064
rect 22980 24012 22986 24064
rect 25314 24012 25320 24064
rect 25372 24012 25378 24064
rect 26970 24012 26976 24064
rect 27028 24012 27034 24064
rect 27890 24012 27896 24064
rect 27948 24012 27954 24064
rect 28534 24012 28540 24064
rect 28592 24012 28598 24064
rect 32674 24012 32680 24064
rect 32732 24012 32738 24064
rect 33042 24012 33048 24064
rect 33100 24012 33106 24064
rect 36446 24012 36452 24064
rect 36504 24012 36510 24064
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 9677 23851 9735 23857
rect 9677 23817 9689 23851
rect 9723 23848 9735 23851
rect 9950 23848 9956 23860
rect 9723 23820 9956 23848
rect 9723 23817 9735 23820
rect 9677 23811 9735 23817
rect 9950 23808 9956 23820
rect 10008 23808 10014 23860
rect 10042 23808 10048 23860
rect 10100 23848 10106 23860
rect 10137 23851 10195 23857
rect 10137 23848 10149 23851
rect 10100 23820 10149 23848
rect 10100 23808 10106 23820
rect 10137 23817 10149 23820
rect 10183 23817 10195 23851
rect 10137 23811 10195 23817
rect 10502 23808 10508 23860
rect 10560 23808 10566 23860
rect 10594 23808 10600 23860
rect 10652 23848 10658 23860
rect 10689 23851 10747 23857
rect 10689 23848 10701 23851
rect 10652 23820 10701 23848
rect 10652 23808 10658 23820
rect 10689 23817 10701 23820
rect 10735 23817 10747 23851
rect 11330 23848 11336 23860
rect 10689 23811 10747 23817
rect 11256 23820 11336 23848
rect 8938 23740 8944 23792
rect 8996 23740 9002 23792
rect 11256 23789 11284 23820
rect 11330 23808 11336 23820
rect 11388 23808 11394 23860
rect 11885 23851 11943 23857
rect 11885 23817 11897 23851
rect 11931 23848 11943 23851
rect 11974 23848 11980 23860
rect 11931 23820 11980 23848
rect 11931 23817 11943 23820
rect 11885 23811 11943 23817
rect 11974 23808 11980 23820
rect 12032 23848 12038 23860
rect 12032 23820 12434 23848
rect 12032 23808 12038 23820
rect 11241 23783 11299 23789
rect 11241 23780 11253 23783
rect 10060 23752 11253 23780
rect 10060 23721 10088 23752
rect 11241 23749 11253 23752
rect 11287 23749 11299 23783
rect 11241 23743 11299 23749
rect 11514 23740 11520 23792
rect 11572 23740 11578 23792
rect 11717 23783 11775 23789
rect 11717 23780 11729 23783
rect 11624 23752 11729 23780
rect 10045 23715 10103 23721
rect 10045 23681 10057 23715
rect 10091 23681 10103 23715
rect 10045 23675 10103 23681
rect 10318 23672 10324 23724
rect 10376 23672 10382 23724
rect 10502 23672 10508 23724
rect 10560 23712 10566 23724
rect 10597 23715 10655 23721
rect 10597 23712 10609 23715
rect 10560 23684 10609 23712
rect 10560 23672 10566 23684
rect 10597 23681 10609 23684
rect 10643 23681 10655 23715
rect 10597 23675 10655 23681
rect 10873 23715 10931 23721
rect 10873 23681 10885 23715
rect 10919 23712 10931 23715
rect 11054 23712 11060 23724
rect 10919 23684 11060 23712
rect 10919 23681 10931 23684
rect 10873 23675 10931 23681
rect 11054 23672 11060 23684
rect 11112 23672 11118 23724
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 7926 23604 7932 23656
rect 7984 23604 7990 23656
rect 8205 23647 8263 23653
rect 8205 23613 8217 23647
rect 8251 23644 8263 23647
rect 8251 23616 11100 23644
rect 8251 23613 8263 23616
rect 8205 23607 8263 23613
rect 9950 23536 9956 23588
rect 10008 23536 10014 23588
rect 11072 23585 11100 23616
rect 11057 23579 11115 23585
rect 11057 23545 11069 23579
rect 11103 23545 11115 23579
rect 11057 23539 11115 23545
rect 9968 23508 9996 23536
rect 11164 23508 11192 23675
rect 11330 23672 11336 23724
rect 11388 23712 11394 23724
rect 11624 23712 11652 23752
rect 11717 23749 11729 23752
rect 11763 23749 11775 23783
rect 12406 23780 12434 23820
rect 12894 23808 12900 23860
rect 12952 23808 12958 23860
rect 16298 23808 16304 23860
rect 16356 23848 16362 23860
rect 16945 23851 17003 23857
rect 16945 23848 16957 23851
rect 16356 23820 16957 23848
rect 16356 23808 16362 23820
rect 16945 23817 16957 23820
rect 16991 23817 17003 23851
rect 16945 23811 17003 23817
rect 17954 23808 17960 23860
rect 18012 23808 18018 23860
rect 18506 23808 18512 23860
rect 18564 23808 18570 23860
rect 20530 23808 20536 23860
rect 20588 23848 20594 23860
rect 20993 23851 21051 23857
rect 20993 23848 21005 23851
rect 20588 23820 21005 23848
rect 20588 23808 20594 23820
rect 20993 23817 21005 23820
rect 21039 23817 21051 23851
rect 20993 23811 21051 23817
rect 24302 23808 24308 23860
rect 24360 23848 24366 23860
rect 24581 23851 24639 23857
rect 24581 23848 24593 23851
rect 24360 23820 24593 23848
rect 24360 23808 24366 23820
rect 24581 23817 24593 23820
rect 24627 23817 24639 23851
rect 24581 23811 24639 23817
rect 25314 23808 25320 23860
rect 25372 23848 25378 23860
rect 25409 23851 25467 23857
rect 25409 23848 25421 23851
rect 25372 23820 25421 23848
rect 25372 23808 25378 23820
rect 25409 23817 25421 23820
rect 25455 23817 25467 23851
rect 25409 23811 25467 23817
rect 25682 23808 25688 23860
rect 25740 23808 25746 23860
rect 26970 23808 26976 23860
rect 27028 23808 27034 23860
rect 27338 23808 27344 23860
rect 27396 23808 27402 23860
rect 27709 23851 27767 23857
rect 27709 23817 27721 23851
rect 27755 23848 27767 23851
rect 28166 23848 28172 23860
rect 27755 23820 28172 23848
rect 27755 23817 27767 23820
rect 27709 23811 27767 23817
rect 28166 23808 28172 23820
rect 28224 23808 28230 23860
rect 28534 23808 28540 23860
rect 28592 23808 28598 23860
rect 32674 23808 32680 23860
rect 32732 23848 32738 23860
rect 32732 23820 33916 23848
rect 32732 23808 32738 23820
rect 13354 23780 13360 23792
rect 12406 23752 13360 23780
rect 11717 23743 11775 23749
rect 13354 23740 13360 23752
rect 13412 23740 13418 23792
rect 17972 23780 18000 23808
rect 16500 23752 18000 23780
rect 19720 23752 22094 23780
rect 11388 23684 11652 23712
rect 12713 23715 12771 23721
rect 11388 23672 11394 23684
rect 12713 23681 12725 23715
rect 12759 23712 12771 23715
rect 12986 23712 12992 23724
rect 12759 23684 12992 23712
rect 12759 23681 12771 23684
rect 12713 23675 12771 23681
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 13078 23672 13084 23724
rect 13136 23672 13142 23724
rect 16500 23721 16528 23752
rect 14645 23715 14703 23721
rect 14645 23681 14657 23715
rect 14691 23712 14703 23715
rect 14737 23715 14795 23721
rect 14737 23712 14749 23715
rect 14691 23684 14749 23712
rect 14691 23681 14703 23684
rect 14645 23675 14703 23681
rect 14737 23681 14749 23684
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 16485 23715 16543 23721
rect 16485 23681 16497 23715
rect 16531 23681 16543 23715
rect 16485 23675 16543 23681
rect 17129 23715 17187 23721
rect 17129 23681 17141 23715
rect 17175 23712 17187 23715
rect 17175 23684 17448 23712
rect 17175 23681 17187 23684
rect 17129 23675 17187 23681
rect 12526 23604 12532 23656
rect 12584 23644 12590 23656
rect 13096 23644 13124 23672
rect 12584 23616 13124 23644
rect 12584 23604 12590 23616
rect 13262 23604 13268 23656
rect 13320 23644 13326 23656
rect 14001 23647 14059 23653
rect 14001 23644 14013 23647
rect 13320 23616 14013 23644
rect 13320 23604 13326 23616
rect 14001 23613 14013 23616
rect 14047 23613 14059 23647
rect 14001 23607 14059 23613
rect 16209 23647 16267 23653
rect 16209 23613 16221 23647
rect 16255 23644 16267 23647
rect 17218 23644 17224 23656
rect 16255 23616 17224 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 17218 23604 17224 23616
rect 17276 23644 17282 23656
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 17276 23616 17325 23644
rect 17276 23604 17282 23616
rect 17313 23613 17325 23616
rect 17359 23613 17371 23647
rect 17420 23644 17448 23684
rect 17494 23672 17500 23724
rect 17552 23712 17558 23724
rect 17589 23715 17647 23721
rect 17589 23712 17601 23715
rect 17552 23684 17601 23712
rect 17552 23672 17558 23684
rect 17589 23681 17601 23684
rect 17635 23681 17647 23715
rect 17589 23675 17647 23681
rect 17773 23715 17831 23721
rect 17773 23681 17785 23715
rect 17819 23681 17831 23715
rect 17773 23675 17831 23681
rect 17420 23616 17632 23644
rect 17313 23607 17371 23613
rect 16393 23579 16451 23585
rect 16393 23545 16405 23579
rect 16439 23576 16451 23579
rect 16942 23576 16948 23588
rect 16439 23548 16948 23576
rect 16439 23545 16451 23548
rect 16393 23539 16451 23545
rect 16942 23536 16948 23548
rect 17000 23536 17006 23588
rect 11606 23508 11612 23520
rect 9968 23480 11612 23508
rect 11606 23468 11612 23480
rect 11664 23508 11670 23520
rect 11701 23511 11759 23517
rect 11701 23508 11713 23511
rect 11664 23480 11713 23508
rect 11664 23468 11670 23480
rect 11701 23477 11713 23480
rect 11747 23477 11759 23511
rect 11701 23471 11759 23477
rect 14366 23468 14372 23520
rect 14424 23508 14430 23520
rect 14829 23511 14887 23517
rect 14829 23508 14841 23511
rect 14424 23480 14841 23508
rect 14424 23468 14430 23480
rect 14829 23477 14841 23480
rect 14875 23477 14887 23511
rect 14829 23471 14887 23477
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 17604 23517 17632 23616
rect 17788 23576 17816 23675
rect 18046 23672 18052 23724
rect 18104 23672 18110 23724
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 18325 23715 18383 23721
rect 18325 23712 18337 23715
rect 18279 23684 18337 23712
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 18325 23681 18337 23684
rect 18371 23681 18383 23715
rect 18325 23675 18383 23681
rect 19058 23672 19064 23724
rect 19116 23712 19122 23724
rect 19613 23715 19671 23721
rect 19613 23712 19625 23715
rect 19116 23684 19625 23712
rect 19116 23672 19122 23684
rect 19613 23681 19625 23684
rect 19659 23681 19671 23715
rect 19613 23675 19671 23681
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18598 23644 18604 23656
rect 17911 23616 18604 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18598 23604 18604 23616
rect 18656 23644 18662 23656
rect 19720 23644 19748 23752
rect 19880 23715 19938 23721
rect 19880 23681 19892 23715
rect 19926 23712 19938 23715
rect 20254 23712 20260 23724
rect 19926 23684 20260 23712
rect 19926 23681 19938 23684
rect 19880 23675 19938 23681
rect 20254 23672 20260 23684
rect 20312 23672 20318 23724
rect 18656 23616 19748 23644
rect 18656 23604 18662 23616
rect 18322 23576 18328 23588
rect 17788 23548 18328 23576
rect 18322 23536 18328 23548
rect 18380 23576 18386 23588
rect 19426 23576 19432 23588
rect 18380 23548 19432 23576
rect 18380 23536 18386 23548
rect 19426 23536 19432 23548
rect 19484 23536 19490 23588
rect 22066 23576 22094 23752
rect 22738 23672 22744 23724
rect 22796 23712 22802 23724
rect 23382 23712 23388 23724
rect 22796 23684 23388 23712
rect 22796 23672 22802 23684
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 25317 23715 25375 23721
rect 25317 23712 25329 23715
rect 23492 23684 25329 23712
rect 22373 23647 22431 23653
rect 22373 23613 22385 23647
rect 22419 23644 22431 23647
rect 22462 23644 22468 23656
rect 22419 23616 22468 23644
rect 22419 23613 22431 23616
rect 22373 23607 22431 23613
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 22646 23604 22652 23656
rect 22704 23604 22710 23656
rect 22830 23604 22836 23656
rect 22888 23644 22894 23656
rect 23492 23644 23520 23684
rect 25317 23681 25329 23684
rect 25363 23681 25375 23715
rect 25317 23675 25375 23681
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23681 25651 23715
rect 25593 23675 25651 23681
rect 22888 23616 23520 23644
rect 22888 23604 22894 23616
rect 25038 23604 25044 23656
rect 25096 23644 25102 23656
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 25096 23616 25145 23644
rect 25096 23604 25102 23616
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 25222 23604 25228 23656
rect 25280 23644 25286 23656
rect 25608 23644 25636 23675
rect 25774 23672 25780 23724
rect 25832 23712 25838 23724
rect 26237 23715 26295 23721
rect 26237 23712 26249 23715
rect 25832 23684 26249 23712
rect 25832 23672 25838 23684
rect 26237 23681 26249 23684
rect 26283 23681 26295 23715
rect 26237 23675 26295 23681
rect 26510 23672 26516 23724
rect 26568 23672 26574 23724
rect 26697 23715 26755 23721
rect 26697 23681 26709 23715
rect 26743 23712 26755 23715
rect 26988 23712 27016 23808
rect 26743 23684 27016 23712
rect 26743 23681 26755 23684
rect 26697 23675 26755 23681
rect 26878 23644 26884 23656
rect 25280 23616 26884 23644
rect 25280 23604 25286 23616
rect 26878 23604 26884 23616
rect 26936 23604 26942 23656
rect 26973 23647 27031 23653
rect 26973 23613 26985 23647
rect 27019 23644 27031 23647
rect 27356 23644 27384 23808
rect 28552 23780 28580 23808
rect 28822 23783 28880 23789
rect 28822 23780 28834 23783
rect 28552 23752 28834 23780
rect 28822 23749 28834 23752
rect 28868 23749 28880 23783
rect 28822 23743 28880 23749
rect 32950 23740 32956 23792
rect 33008 23780 33014 23792
rect 33888 23789 33916 23820
rect 35158 23808 35164 23860
rect 35216 23848 35222 23860
rect 35805 23851 35863 23857
rect 35805 23848 35817 23851
rect 35216 23820 35817 23848
rect 35216 23808 35222 23820
rect 35805 23817 35817 23820
rect 35851 23817 35863 23851
rect 35805 23811 35863 23817
rect 33137 23783 33195 23789
rect 33137 23780 33149 23783
rect 33008 23752 33149 23780
rect 33008 23740 33014 23752
rect 33137 23749 33149 23752
rect 33183 23749 33195 23783
rect 33137 23743 33195 23749
rect 33873 23783 33931 23789
rect 33873 23749 33885 23783
rect 33919 23749 33931 23783
rect 36262 23780 36268 23792
rect 33873 23743 33931 23749
rect 36004 23752 36268 23780
rect 33152 23712 33180 23743
rect 34057 23715 34115 23721
rect 34057 23712 34069 23715
rect 33152 23684 34069 23712
rect 34057 23681 34069 23684
rect 34103 23681 34115 23715
rect 34057 23675 34115 23681
rect 34146 23672 34152 23724
rect 34204 23672 34210 23724
rect 36004 23721 36032 23752
rect 36262 23740 36268 23752
rect 36320 23780 36326 23792
rect 36320 23752 37136 23780
rect 36320 23740 36326 23752
rect 37108 23724 37136 23752
rect 35989 23715 36047 23721
rect 35989 23681 36001 23715
rect 36035 23681 36047 23715
rect 35989 23675 36047 23681
rect 36173 23715 36231 23721
rect 36173 23681 36185 23715
rect 36219 23712 36231 23715
rect 36354 23712 36360 23724
rect 36219 23684 36360 23712
rect 36219 23681 36231 23684
rect 36173 23675 36231 23681
rect 36354 23672 36360 23684
rect 36412 23672 36418 23724
rect 36538 23672 36544 23724
rect 36596 23672 36602 23724
rect 37090 23672 37096 23724
rect 37148 23672 37154 23724
rect 27019 23616 27384 23644
rect 27617 23647 27675 23653
rect 27019 23613 27031 23616
rect 26973 23607 27031 23613
rect 27617 23613 27629 23647
rect 27663 23644 27675 23647
rect 27706 23644 27712 23656
rect 27663 23616 27712 23644
rect 27663 23613 27675 23616
rect 27617 23607 27675 23613
rect 27706 23604 27712 23616
rect 27764 23604 27770 23656
rect 29086 23604 29092 23656
rect 29144 23604 29150 23656
rect 29917 23647 29975 23653
rect 29917 23613 29929 23647
rect 29963 23644 29975 23647
rect 30558 23644 30564 23656
rect 29963 23616 30564 23644
rect 29963 23613 29975 23616
rect 29917 23607 29975 23613
rect 30558 23604 30564 23616
rect 30616 23644 30622 23656
rect 30926 23644 30932 23656
rect 30616 23616 30932 23644
rect 30616 23604 30622 23616
rect 30926 23604 30932 23616
rect 30984 23644 30990 23656
rect 31021 23647 31079 23653
rect 31021 23644 31033 23647
rect 30984 23616 31033 23644
rect 30984 23604 30990 23616
rect 31021 23613 31033 23616
rect 31067 23613 31079 23647
rect 31021 23607 31079 23613
rect 33042 23604 33048 23656
rect 33100 23644 33106 23656
rect 33689 23647 33747 23653
rect 33689 23644 33701 23647
rect 33100 23616 33701 23644
rect 33100 23604 33106 23616
rect 33689 23613 33701 23616
rect 33735 23613 33747 23647
rect 33689 23607 33747 23613
rect 33870 23604 33876 23656
rect 33928 23644 33934 23656
rect 33928 23616 34192 23644
rect 33928 23604 33934 23616
rect 27154 23576 27160 23588
rect 22066 23548 27160 23576
rect 27154 23536 27160 23548
rect 27212 23576 27218 23588
rect 27522 23576 27528 23588
rect 27212 23548 27528 23576
rect 27212 23536 27218 23548
rect 27522 23536 27528 23548
rect 27580 23536 27586 23588
rect 30190 23536 30196 23588
rect 30248 23536 30254 23588
rect 30377 23579 30435 23585
rect 30377 23545 30389 23579
rect 30423 23576 30435 23579
rect 32582 23576 32588 23588
rect 30423 23548 32588 23576
rect 30423 23545 30435 23548
rect 30377 23539 30435 23545
rect 32582 23536 32588 23548
rect 32640 23536 32646 23588
rect 34054 23536 34060 23588
rect 34112 23536 34118 23588
rect 34164 23576 34192 23616
rect 36078 23604 36084 23656
rect 36136 23604 36142 23656
rect 36265 23647 36323 23653
rect 36265 23613 36277 23647
rect 36311 23613 36323 23647
rect 36372 23644 36400 23672
rect 36722 23644 36728 23656
rect 36372 23616 36728 23644
rect 36265 23607 36323 23613
rect 36280 23576 36308 23607
rect 36722 23604 36728 23616
rect 36780 23604 36786 23656
rect 36814 23604 36820 23656
rect 36872 23604 36878 23656
rect 36354 23576 36360 23588
rect 34164 23548 36360 23576
rect 36354 23536 36360 23548
rect 36412 23536 36418 23588
rect 36630 23536 36636 23588
rect 36688 23536 36694 23588
rect 16301 23511 16359 23517
rect 16301 23508 16313 23511
rect 15988 23480 16313 23508
rect 15988 23468 15994 23480
rect 16301 23477 16313 23480
rect 16347 23477 16359 23511
rect 16301 23471 16359 23477
rect 17589 23511 17647 23517
rect 17589 23477 17601 23511
rect 17635 23508 17647 23511
rect 18414 23508 18420 23520
rect 17635 23480 18420 23508
rect 17635 23477 17647 23480
rect 17589 23471 17647 23477
rect 18414 23468 18420 23480
rect 18472 23468 18478 23520
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 23290 23508 23296 23520
rect 20036 23480 23296 23508
rect 20036 23468 20042 23480
rect 23290 23468 23296 23480
rect 23348 23508 23354 23520
rect 24578 23508 24584 23520
rect 23348 23480 24584 23508
rect 23348 23468 23354 23480
rect 24578 23468 24584 23480
rect 24636 23468 24642 23520
rect 25590 23468 25596 23520
rect 25648 23468 25654 23520
rect 26694 23468 26700 23520
rect 26752 23468 26758 23520
rect 30466 23468 30472 23520
rect 30524 23468 30530 23520
rect 33873 23511 33931 23517
rect 33873 23477 33885 23511
rect 33919 23508 33931 23511
rect 34072 23508 34100 23536
rect 33919 23480 34100 23508
rect 36725 23511 36783 23517
rect 33919 23477 33931 23480
rect 33873 23471 33931 23477
rect 36725 23477 36737 23511
rect 36771 23508 36783 23511
rect 37274 23508 37280 23520
rect 36771 23480 37280 23508
rect 36771 23477 36783 23480
rect 36725 23471 36783 23477
rect 37274 23468 37280 23480
rect 37332 23468 37338 23520
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 8938 23264 8944 23316
rect 8996 23304 9002 23316
rect 9033 23307 9091 23313
rect 9033 23304 9045 23307
rect 8996 23276 9045 23304
rect 8996 23264 9002 23276
rect 9033 23273 9045 23276
rect 9079 23273 9091 23307
rect 9033 23267 9091 23273
rect 11054 23264 11060 23316
rect 11112 23304 11118 23316
rect 11149 23307 11207 23313
rect 11149 23304 11161 23307
rect 11112 23276 11161 23304
rect 11112 23264 11118 23276
rect 11149 23273 11161 23276
rect 11195 23273 11207 23307
rect 11149 23267 11207 23273
rect 11333 23307 11391 23313
rect 11333 23273 11345 23307
rect 11379 23304 11391 23307
rect 12989 23307 13047 23313
rect 11379 23276 11744 23304
rect 11379 23273 11391 23276
rect 11333 23267 11391 23273
rect 11606 23196 11612 23248
rect 11664 23196 11670 23248
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8864 23072 8953 23100
rect 8864 23044 8892 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 10134 23060 10140 23112
rect 10192 23060 10198 23112
rect 11624 23109 11652 23196
rect 11716 23109 11744 23276
rect 12989 23273 13001 23307
rect 13035 23304 13047 23307
rect 13170 23304 13176 23316
rect 13035 23276 13176 23304
rect 13035 23273 13047 23276
rect 12989 23267 13047 23273
rect 13170 23264 13176 23276
rect 13228 23304 13234 23316
rect 14918 23304 14924 23316
rect 13228 23276 14924 23304
rect 13228 23264 13234 23276
rect 14918 23264 14924 23276
rect 14976 23304 14982 23316
rect 16574 23304 16580 23316
rect 14976 23276 16580 23304
rect 14976 23264 14982 23276
rect 16574 23264 16580 23276
rect 16632 23264 16638 23316
rect 16684 23276 17632 23304
rect 16684 23248 16712 23276
rect 16666 23196 16672 23248
rect 16724 23196 16730 23248
rect 17126 23196 17132 23248
rect 17184 23196 17190 23248
rect 11882 23128 11888 23180
rect 11940 23168 11946 23180
rect 12526 23168 12532 23180
rect 11940 23140 12532 23168
rect 11940 23128 11946 23140
rect 12526 23128 12532 23140
rect 12584 23128 12590 23180
rect 12621 23171 12679 23177
rect 12621 23137 12633 23171
rect 12667 23168 12679 23171
rect 12667 23140 12940 23168
rect 12667 23137 12679 23140
rect 12621 23131 12679 23137
rect 11609 23103 11667 23109
rect 11609 23069 11621 23103
rect 11655 23069 11667 23103
rect 11609 23063 11667 23069
rect 11701 23103 11759 23109
rect 11701 23069 11713 23103
rect 11747 23100 11759 23103
rect 12437 23103 12495 23109
rect 12437 23100 12449 23103
rect 11747 23072 12449 23100
rect 11747 23069 11759 23072
rect 11701 23063 11759 23069
rect 12437 23069 12449 23072
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 12802 23060 12808 23112
rect 12860 23060 12866 23112
rect 8846 22992 8852 23044
rect 8904 22992 8910 23044
rect 10594 22992 10600 23044
rect 10652 23032 10658 23044
rect 11330 23041 11336 23044
rect 11317 23035 11336 23041
rect 10652 23004 10824 23032
rect 10652 22992 10658 23004
rect 10686 22924 10692 22976
rect 10744 22924 10750 22976
rect 10796 22964 10824 23004
rect 11317 23001 11329 23035
rect 11317 22995 11336 23001
rect 11330 22992 11336 22995
rect 11388 22992 11394 23044
rect 11517 23035 11575 23041
rect 11517 23001 11529 23035
rect 11563 23032 11575 23035
rect 11882 23032 11888 23044
rect 11563 23004 11888 23032
rect 11563 23001 11575 23004
rect 11517 22995 11575 23001
rect 11882 22992 11888 23004
rect 11940 22992 11946 23044
rect 12912 23032 12940 23140
rect 13814 23128 13820 23180
rect 13872 23168 13878 23180
rect 14090 23168 14096 23180
rect 13872 23140 14096 23168
rect 13872 23128 13878 23140
rect 14090 23128 14096 23140
rect 14148 23168 14154 23180
rect 14550 23168 14556 23180
rect 14148 23140 14556 23168
rect 14148 23128 14154 23140
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 15948 23140 16896 23168
rect 15948 23112 15976 23140
rect 13170 23060 13176 23112
rect 13228 23060 13234 23112
rect 14366 23060 14372 23112
rect 14424 23060 14430 23112
rect 14461 23103 14519 23109
rect 14461 23069 14473 23103
rect 14507 23100 14519 23103
rect 15930 23100 15936 23112
rect 14507 23072 15936 23100
rect 14507 23069 14519 23072
rect 14461 23063 14519 23069
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 16114 23060 16120 23112
rect 16172 23060 16178 23112
rect 16868 23109 16896 23140
rect 17494 23128 17500 23180
rect 17552 23128 17558 23180
rect 17604 23168 17632 23276
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 18141 23307 18199 23313
rect 18141 23304 18153 23307
rect 18104 23276 18153 23304
rect 18104 23264 18110 23276
rect 18141 23273 18153 23276
rect 18187 23273 18199 23307
rect 18141 23267 18199 23273
rect 20254 23264 20260 23316
rect 20312 23304 20318 23316
rect 20349 23307 20407 23313
rect 20349 23304 20361 23307
rect 20312 23276 20361 23304
rect 20312 23264 20318 23276
rect 20349 23273 20361 23276
rect 20395 23273 20407 23307
rect 25222 23304 25228 23316
rect 20349 23267 20407 23273
rect 20456 23276 25228 23304
rect 18233 23171 18291 23177
rect 18233 23168 18245 23171
rect 17604 23140 18245 23168
rect 18233 23137 18245 23140
rect 18279 23137 18291 23171
rect 20456 23168 20484 23276
rect 25222 23264 25228 23276
rect 25280 23264 25286 23316
rect 25774 23264 25780 23316
rect 25832 23304 25838 23316
rect 25961 23307 26019 23313
rect 25961 23304 25973 23307
rect 25832 23276 25973 23304
rect 25832 23264 25838 23276
rect 25961 23273 25973 23276
rect 26007 23273 26019 23307
rect 25961 23267 26019 23273
rect 27433 23307 27491 23313
rect 27433 23273 27445 23307
rect 27479 23304 27491 23307
rect 27706 23304 27712 23316
rect 27479 23276 27712 23304
rect 27479 23273 27491 23276
rect 27433 23267 27491 23273
rect 27706 23264 27712 23276
rect 27764 23264 27770 23316
rect 27890 23264 27896 23316
rect 27948 23304 27954 23316
rect 27985 23307 28043 23313
rect 27985 23304 27997 23307
rect 27948 23276 27997 23304
rect 27948 23264 27954 23276
rect 27985 23273 27997 23276
rect 28031 23273 28043 23307
rect 27985 23267 28043 23273
rect 28169 23307 28227 23313
rect 28169 23273 28181 23307
rect 28215 23304 28227 23307
rect 28350 23304 28356 23316
rect 28215 23276 28356 23304
rect 28215 23273 28227 23276
rect 28169 23267 28227 23273
rect 28350 23264 28356 23276
rect 28408 23264 28414 23316
rect 28445 23307 28503 23313
rect 28445 23273 28457 23307
rect 28491 23304 28503 23307
rect 29546 23304 29552 23316
rect 28491 23276 29552 23304
rect 28491 23273 28503 23276
rect 28445 23267 28503 23273
rect 27614 23196 27620 23248
rect 27672 23196 27678 23248
rect 28460 23168 28488 23267
rect 29546 23264 29552 23276
rect 29604 23264 29610 23316
rect 30926 23264 30932 23316
rect 30984 23264 30990 23316
rect 31389 23307 31447 23313
rect 31389 23273 31401 23307
rect 31435 23304 31447 23307
rect 31478 23304 31484 23316
rect 31435 23276 31484 23304
rect 31435 23273 31447 23276
rect 31389 23267 31447 23273
rect 31478 23264 31484 23276
rect 31536 23264 31542 23316
rect 32585 23307 32643 23313
rect 32585 23273 32597 23307
rect 32631 23273 32643 23307
rect 32585 23267 32643 23273
rect 32769 23307 32827 23313
rect 32769 23273 32781 23307
rect 32815 23304 32827 23307
rect 32858 23304 32864 23316
rect 32815 23276 32864 23304
rect 32815 23273 32827 23276
rect 32769 23267 32827 23273
rect 32600 23236 32628 23267
rect 32858 23264 32864 23276
rect 32916 23264 32922 23316
rect 32950 23264 32956 23316
rect 33008 23264 33014 23316
rect 35342 23264 35348 23316
rect 35400 23304 35406 23316
rect 35437 23307 35495 23313
rect 35437 23304 35449 23307
rect 35400 23276 35449 23304
rect 35400 23264 35406 23276
rect 35437 23273 35449 23276
rect 35483 23273 35495 23307
rect 35437 23267 35495 23273
rect 35526 23264 35532 23316
rect 35584 23264 35590 23316
rect 36081 23307 36139 23313
rect 36081 23273 36093 23307
rect 36127 23304 36139 23307
rect 36630 23304 36636 23316
rect 36127 23276 36636 23304
rect 36127 23273 36139 23276
rect 36081 23267 36139 23273
rect 36630 23264 36636 23276
rect 36688 23264 36694 23316
rect 35253 23239 35311 23245
rect 32232 23208 34100 23236
rect 32232 23180 32260 23208
rect 18233 23131 18291 23137
rect 20180 23140 20484 23168
rect 28000 23140 28488 23168
rect 16853 23103 16911 23109
rect 16853 23069 16865 23103
rect 16899 23069 16911 23103
rect 16853 23063 16911 23069
rect 17129 23103 17187 23109
rect 17129 23069 17141 23103
rect 17175 23100 17187 23103
rect 17218 23100 17224 23112
rect 17175 23072 17224 23100
rect 17175 23069 17187 23072
rect 17129 23063 17187 23069
rect 17218 23060 17224 23072
rect 17276 23100 17282 23112
rect 17586 23100 17592 23112
rect 17276 23072 17592 23100
rect 17276 23060 17282 23072
rect 17586 23060 17592 23072
rect 17644 23100 17650 23112
rect 17681 23103 17739 23109
rect 17681 23100 17693 23103
rect 17644 23072 17693 23100
rect 17644 23060 17650 23072
rect 17681 23069 17693 23072
rect 17727 23069 17739 23103
rect 17681 23063 17739 23069
rect 18414 23060 18420 23112
rect 18472 23060 18478 23112
rect 20180 23109 20208 23140
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23100 18659 23103
rect 18693 23103 18751 23109
rect 18693 23100 18705 23103
rect 18647 23072 18705 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 18693 23069 18705 23072
rect 18739 23069 18751 23103
rect 20165 23103 20223 23109
rect 20165 23100 20177 23103
rect 18693 23063 18751 23069
rect 19306 23072 20177 23100
rect 14826 23041 14832 23044
rect 12406 23004 12940 23032
rect 12406 22964 12434 23004
rect 12912 22976 12940 23004
rect 14185 23035 14243 23041
rect 14185 23001 14197 23035
rect 14231 23032 14243 23035
rect 14231 23004 14412 23032
rect 14231 23001 14243 23004
rect 14185 22995 14243 23001
rect 10796 22936 12434 22964
rect 12526 22924 12532 22976
rect 12584 22924 12590 22976
rect 12710 22924 12716 22976
rect 12768 22924 12774 22976
rect 12894 22924 12900 22976
rect 12952 22924 12958 22976
rect 14274 22924 14280 22976
rect 14332 22973 14338 22976
rect 14332 22927 14341 22973
rect 14384 22964 14412 23004
rect 14820 22995 14832 23041
rect 14826 22992 14832 22995
rect 14884 22992 14890 23044
rect 19306 23032 19334 23072
rect 20165 23069 20177 23072
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 20349 23103 20407 23109
rect 20349 23069 20361 23103
rect 20395 23100 20407 23103
rect 22830 23100 22836 23112
rect 20395 23072 22836 23100
rect 20395 23069 20407 23072
rect 20349 23063 20407 23069
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 23106 23060 23112 23112
rect 23164 23100 23170 23112
rect 23201 23103 23259 23109
rect 23201 23100 23213 23103
rect 23164 23072 23213 23100
rect 23164 23060 23170 23072
rect 23201 23069 23213 23072
rect 23247 23069 23259 23103
rect 23201 23063 23259 23069
rect 24118 23060 24124 23112
rect 24176 23060 24182 23112
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23100 24639 23103
rect 24670 23100 24676 23112
rect 24627 23072 24676 23100
rect 24627 23069 24639 23072
rect 24581 23063 24639 23069
rect 24670 23060 24676 23072
rect 24728 23100 24734 23112
rect 26050 23100 26056 23112
rect 24728 23072 26056 23100
rect 24728 23060 24734 23072
rect 26050 23060 26056 23072
rect 26108 23060 26114 23112
rect 26320 23103 26378 23109
rect 26320 23069 26332 23103
rect 26366 23100 26378 23103
rect 26694 23100 26700 23112
rect 26366 23072 26700 23100
rect 26366 23069 26378 23072
rect 26320 23063 26378 23069
rect 26694 23060 26700 23072
rect 26752 23060 26758 23112
rect 15120 23004 19334 23032
rect 15010 22964 15016 22976
rect 14384 22936 15016 22964
rect 14332 22924 14338 22927
rect 15010 22924 15016 22936
rect 15068 22964 15074 22976
rect 15120 22964 15148 23004
rect 23014 22992 23020 23044
rect 23072 23032 23078 23044
rect 23569 23035 23627 23041
rect 23569 23032 23581 23035
rect 23072 23004 23581 23032
rect 23072 22992 23078 23004
rect 23569 23001 23581 23004
rect 23615 23001 23627 23035
rect 23569 22995 23627 23001
rect 24848 23035 24906 23041
rect 24848 23001 24860 23035
rect 24894 23032 24906 23035
rect 25590 23032 25596 23044
rect 24894 23004 25596 23032
rect 24894 23001 24906 23004
rect 24848 22995 24906 23001
rect 25590 22992 25596 23004
rect 25648 22992 25654 23044
rect 28000 23041 28028 23140
rect 29086 23128 29092 23180
rect 29144 23168 29150 23180
rect 29549 23171 29607 23177
rect 29549 23168 29561 23171
rect 29144 23140 29561 23168
rect 29144 23128 29150 23140
rect 29549 23137 29561 23140
rect 29595 23137 29607 23171
rect 29549 23131 29607 23137
rect 32214 23128 32220 23180
rect 32272 23128 32278 23180
rect 32398 23128 32404 23180
rect 32456 23168 32462 23180
rect 34072 23177 34100 23208
rect 35253 23205 35265 23239
rect 35299 23236 35311 23239
rect 35544 23236 35572 23264
rect 35299 23208 35572 23236
rect 36173 23239 36231 23245
rect 35299 23205 35311 23208
rect 35253 23199 35311 23205
rect 36173 23205 36185 23239
rect 36219 23236 36231 23239
rect 36538 23236 36544 23248
rect 36219 23208 36544 23236
rect 36219 23205 36231 23208
rect 36173 23199 36231 23205
rect 36538 23196 36544 23208
rect 36596 23196 36602 23248
rect 33689 23171 33747 23177
rect 33689 23168 33701 23171
rect 32456 23140 33701 23168
rect 32456 23128 32462 23140
rect 33689 23137 33701 23140
rect 33735 23137 33747 23171
rect 34057 23171 34115 23177
rect 33689 23131 33747 23137
rect 33796 23140 34008 23168
rect 31202 23060 31208 23112
rect 31260 23060 31266 23112
rect 31481 23103 31539 23109
rect 31481 23069 31493 23103
rect 31527 23100 31539 23103
rect 31665 23103 31723 23109
rect 31665 23100 31677 23103
rect 31527 23072 31677 23100
rect 31527 23069 31539 23072
rect 31481 23063 31539 23069
rect 31665 23069 31677 23072
rect 31711 23069 31723 23103
rect 31665 23063 31723 23069
rect 32306 23060 32312 23112
rect 32364 23100 32370 23112
rect 33226 23100 33232 23112
rect 32364 23072 33232 23100
rect 32364 23060 32370 23072
rect 27985 23035 28043 23041
rect 27985 23001 27997 23035
rect 28031 23032 28043 23035
rect 28074 23032 28080 23044
rect 28031 23004 28080 23032
rect 28031 23001 28043 23004
rect 27985 22995 28043 23001
rect 28074 22992 28080 23004
rect 28132 22992 28138 23044
rect 28258 22992 28264 23044
rect 28316 22992 28322 23044
rect 29362 22992 29368 23044
rect 29420 23032 29426 23044
rect 32416 23041 32444 23072
rect 33226 23060 33232 23072
rect 33284 23100 33290 23112
rect 33505 23103 33563 23109
rect 33505 23100 33517 23103
rect 33284 23072 33517 23100
rect 33284 23060 33290 23072
rect 33505 23069 33517 23072
rect 33551 23069 33563 23103
rect 33505 23063 33563 23069
rect 29794 23035 29852 23041
rect 29794 23032 29806 23035
rect 29420 23004 29806 23032
rect 29420 22992 29426 23004
rect 29794 23001 29806 23004
rect 29840 23001 29852 23035
rect 29794 22995 29852 23001
rect 32401 23035 32459 23041
rect 32401 23001 32413 23035
rect 32447 23001 32459 23035
rect 32401 22995 32459 23001
rect 32858 22992 32864 23044
rect 32916 23032 32922 23044
rect 33796 23032 33824 23140
rect 33873 23103 33931 23109
rect 33873 23069 33885 23103
rect 33919 23069 33931 23103
rect 33980 23100 34008 23140
rect 34057 23137 34069 23171
rect 34103 23137 34115 23171
rect 34057 23131 34115 23137
rect 35897 23171 35955 23177
rect 35897 23137 35909 23171
rect 35943 23168 35955 23171
rect 36446 23168 36452 23180
rect 35943 23140 36452 23168
rect 35943 23137 35955 23140
rect 35897 23131 35955 23137
rect 36446 23128 36452 23140
rect 36504 23128 36510 23180
rect 36722 23168 36728 23180
rect 36556 23140 36728 23168
rect 34146 23100 34152 23112
rect 33980 23072 34152 23100
rect 33873 23063 33931 23069
rect 32916 23004 33824 23032
rect 32916 22992 32922 23004
rect 15068 22936 15148 22964
rect 15068 22924 15074 22936
rect 15194 22924 15200 22976
rect 15252 22964 15258 22976
rect 15933 22967 15991 22973
rect 15933 22964 15945 22967
rect 15252 22936 15945 22964
rect 15252 22924 15258 22936
rect 15933 22933 15945 22936
rect 15979 22964 15991 22967
rect 16114 22964 16120 22976
rect 15979 22936 16120 22964
rect 15979 22933 15991 22936
rect 15933 22927 15991 22933
rect 16114 22924 16120 22936
rect 16172 22924 16178 22976
rect 16761 22967 16819 22973
rect 16761 22933 16773 22967
rect 16807 22964 16819 22967
rect 16945 22967 17003 22973
rect 16945 22964 16957 22967
rect 16807 22936 16957 22964
rect 16807 22933 16819 22936
rect 16761 22927 16819 22933
rect 16945 22933 16957 22936
rect 16991 22933 17003 22967
rect 16945 22927 17003 22933
rect 17770 22924 17776 22976
rect 17828 22924 17834 22976
rect 18877 22967 18935 22973
rect 18877 22933 18889 22967
rect 18923 22964 18935 22967
rect 19334 22964 19340 22976
rect 18923 22936 19340 22964
rect 18923 22933 18935 22936
rect 18877 22927 18935 22933
rect 19334 22924 19340 22936
rect 19392 22924 19398 22976
rect 23290 22924 23296 22976
rect 23348 22924 23354 22976
rect 28350 22924 28356 22976
rect 28408 22964 28414 22976
rect 28461 22967 28519 22973
rect 28461 22964 28473 22967
rect 28408 22936 28473 22964
rect 28408 22924 28414 22936
rect 28461 22933 28473 22936
rect 28507 22933 28519 22967
rect 28461 22927 28519 22933
rect 28629 22967 28687 22973
rect 28629 22933 28641 22967
rect 28675 22964 28687 22967
rect 29178 22964 29184 22976
rect 28675 22936 29184 22964
rect 28675 22933 28687 22936
rect 28629 22927 28687 22933
rect 29178 22924 29184 22936
rect 29236 22924 29242 22976
rect 31018 22924 31024 22976
rect 31076 22924 31082 22976
rect 32582 22924 32588 22976
rect 32640 22973 32646 22976
rect 32640 22967 32669 22973
rect 32657 22964 32669 22967
rect 33888 22964 33916 23063
rect 34146 23060 34152 23072
rect 34204 23060 34210 23112
rect 34333 23103 34391 23109
rect 34333 23069 34345 23103
rect 34379 23100 34391 23103
rect 34422 23100 34428 23112
rect 34379 23072 34428 23100
rect 34379 23069 34391 23072
rect 34333 23063 34391 23069
rect 34422 23060 34428 23072
rect 34480 23060 34486 23112
rect 35713 23103 35771 23109
rect 35713 23100 35725 23103
rect 35544 23072 35725 23100
rect 34238 22992 34244 23044
rect 34296 22992 34302 23044
rect 35544 22976 35572 23072
rect 35713 23069 35725 23072
rect 35759 23069 35771 23103
rect 35713 23063 35771 23069
rect 36078 23060 36084 23112
rect 36136 23060 36142 23112
rect 36170 23060 36176 23112
rect 36228 23100 36234 23112
rect 36556 23109 36584 23140
rect 36722 23128 36728 23140
rect 36780 23128 36786 23180
rect 36541 23103 36599 23109
rect 36228 23072 36492 23100
rect 36228 23060 36234 23072
rect 35621 23035 35679 23041
rect 35621 23001 35633 23035
rect 35667 23032 35679 23035
rect 35805 23035 35863 23041
rect 35805 23032 35817 23035
rect 35667 23004 35817 23032
rect 35667 23001 35679 23004
rect 35621 22995 35679 23001
rect 35805 23001 35817 23004
rect 35851 23032 35863 23035
rect 36188 23032 36216 23060
rect 35851 23004 36216 23032
rect 35851 23001 35863 23004
rect 35805 22995 35863 23001
rect 36262 22992 36268 23044
rect 36320 23032 36326 23044
rect 36464 23041 36492 23072
rect 36541 23069 36553 23103
rect 36587 23069 36599 23103
rect 36541 23063 36599 23069
rect 36630 23060 36636 23112
rect 36688 23100 36694 23112
rect 37274 23109 37280 23112
rect 37001 23103 37059 23109
rect 37001 23100 37013 23103
rect 36688 23072 37013 23100
rect 36688 23060 36694 23072
rect 37001 23069 37013 23072
rect 37047 23069 37059 23103
rect 37268 23100 37280 23109
rect 37235 23072 37280 23100
rect 37001 23063 37059 23069
rect 37268 23063 37280 23072
rect 37274 23060 37280 23063
rect 37332 23060 37338 23112
rect 36357 23035 36415 23041
rect 36357 23032 36369 23035
rect 36320 23004 36369 23032
rect 36320 22992 36326 23004
rect 36357 23001 36369 23004
rect 36403 23001 36415 23035
rect 36357 22995 36415 23001
rect 36449 23035 36507 23041
rect 36449 23001 36461 23035
rect 36495 23001 36507 23035
rect 36449 22995 36507 23001
rect 36725 23035 36783 23041
rect 36725 23001 36737 23035
rect 36771 23001 36783 23035
rect 36725 22995 36783 23001
rect 35434 22973 35440 22976
rect 32657 22936 33916 22964
rect 35421 22967 35440 22973
rect 32657 22933 32669 22936
rect 32640 22927 32669 22933
rect 35421 22933 35433 22967
rect 35421 22927 35440 22933
rect 32640 22924 32646 22927
rect 35434 22924 35440 22927
rect 35492 22924 35498 22976
rect 35526 22924 35532 22976
rect 35584 22964 35590 22976
rect 36280 22964 36308 22992
rect 35584 22936 36308 22964
rect 36740 22964 36768 22995
rect 38378 22964 38384 22976
rect 36740 22936 38384 22964
rect 35584 22924 35590 22936
rect 38378 22924 38384 22936
rect 38436 22924 38442 22976
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 10042 22720 10048 22772
rect 10100 22720 10106 22772
rect 10686 22720 10692 22772
rect 10744 22720 10750 22772
rect 11057 22763 11115 22769
rect 11057 22729 11069 22763
rect 11103 22760 11115 22763
rect 11330 22760 11336 22772
rect 11103 22732 11336 22760
rect 11103 22729 11115 22732
rect 11057 22723 11115 22729
rect 11330 22720 11336 22732
rect 11388 22720 11394 22772
rect 11606 22720 11612 22772
rect 11664 22720 11670 22772
rect 13081 22763 13139 22769
rect 13081 22729 13093 22763
rect 13127 22760 13139 22763
rect 13170 22760 13176 22772
rect 13127 22732 13176 22760
rect 13127 22729 13139 22732
rect 13081 22723 13139 22729
rect 13170 22720 13176 22732
rect 13228 22720 13234 22772
rect 13262 22720 13268 22772
rect 13320 22720 13326 22772
rect 14274 22720 14280 22772
rect 14332 22720 14338 22772
rect 14826 22720 14832 22772
rect 14884 22720 14890 22772
rect 15010 22720 15016 22772
rect 15068 22720 15074 22772
rect 17126 22720 17132 22772
rect 17184 22720 17190 22772
rect 21913 22763 21971 22769
rect 21913 22729 21925 22763
rect 21959 22760 21971 22763
rect 22738 22760 22744 22772
rect 21959 22732 22744 22760
rect 21959 22729 21971 22732
rect 21913 22723 21971 22729
rect 22738 22720 22744 22732
rect 22796 22720 22802 22772
rect 23290 22720 23296 22772
rect 23348 22720 23354 22772
rect 23382 22720 23388 22772
rect 23440 22760 23446 22772
rect 23440 22732 23796 22760
rect 23440 22720 23446 22732
rect 8938 22652 8944 22704
rect 8996 22652 9002 22704
rect 10060 22692 10088 22720
rect 10318 22701 10324 22704
rect 10137 22695 10195 22701
rect 10137 22692 10149 22695
rect 9876 22664 10149 22692
rect 9876 22636 9904 22664
rect 10137 22661 10149 22664
rect 10183 22661 10195 22695
rect 10137 22655 10195 22661
rect 10275 22695 10324 22701
rect 10275 22661 10287 22695
rect 10321 22661 10324 22695
rect 10275 22655 10324 22661
rect 10318 22652 10324 22655
rect 10376 22652 10382 22704
rect 10704 22692 10732 22720
rect 10428 22664 10732 22692
rect 10781 22695 10839 22701
rect 7926 22584 7932 22636
rect 7984 22584 7990 22636
rect 9858 22584 9864 22636
rect 9916 22584 9922 22636
rect 9950 22584 9956 22636
rect 10008 22584 10014 22636
rect 10428 22633 10456 22664
rect 10781 22661 10793 22695
rect 10827 22692 10839 22695
rect 10827 22664 11192 22692
rect 10827 22661 10839 22664
rect 10781 22655 10839 22661
rect 11164 22636 11192 22664
rect 10045 22627 10103 22633
rect 10045 22593 10057 22627
rect 10091 22593 10103 22627
rect 10045 22587 10103 22593
rect 10413 22627 10471 22633
rect 10413 22593 10425 22627
rect 10459 22593 10471 22627
rect 10413 22587 10471 22593
rect 8205 22559 8263 22565
rect 8205 22525 8217 22559
rect 8251 22556 8263 22559
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 8251 22528 9781 22556
rect 8251 22525 8263 22528
rect 8205 22519 8263 22525
rect 9769 22525 9781 22528
rect 9815 22525 9827 22559
rect 10060 22556 10088 22587
rect 10594 22584 10600 22636
rect 10652 22624 10658 22636
rect 10689 22627 10747 22633
rect 10689 22624 10701 22627
rect 10652 22596 10701 22624
rect 10652 22584 10658 22596
rect 10689 22593 10701 22596
rect 10735 22593 10747 22627
rect 10689 22587 10747 22593
rect 10870 22584 10876 22636
rect 10928 22584 10934 22636
rect 11146 22584 11152 22636
rect 11204 22584 11210 22636
rect 11348 22633 11376 22720
rect 11333 22627 11391 22633
rect 11333 22593 11345 22627
rect 11379 22593 11391 22627
rect 11624 22624 11652 22720
rect 12161 22695 12219 22701
rect 12161 22692 12173 22695
rect 11992 22664 12173 22692
rect 11992 22633 12020 22664
rect 12161 22661 12173 22664
rect 12207 22692 12219 22695
rect 14292 22692 14320 22720
rect 14378 22695 14436 22701
rect 14378 22692 14390 22695
rect 12207 22664 13676 22692
rect 14292 22664 14390 22692
rect 12207 22661 12219 22664
rect 12161 22655 12219 22661
rect 11701 22627 11759 22633
rect 11701 22624 11713 22627
rect 11624 22596 11713 22624
rect 11333 22587 11391 22593
rect 11701 22593 11713 22596
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 11977 22627 12035 22633
rect 11977 22593 11989 22627
rect 12023 22593 12035 22627
rect 11977 22587 12035 22593
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22624 12127 22627
rect 12345 22627 12403 22633
rect 12115 22596 12204 22624
rect 12115 22593 12127 22596
rect 12069 22587 12127 22593
rect 12176 22568 12204 22596
rect 12345 22593 12357 22627
rect 12391 22624 12403 22627
rect 12434 22624 12440 22636
rect 12391 22596 12440 22624
rect 12391 22593 12403 22596
rect 12345 22587 12403 22593
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12529 22627 12587 22633
rect 12529 22593 12541 22627
rect 12575 22624 12587 22627
rect 12621 22627 12679 22633
rect 12621 22624 12633 22627
rect 12575 22596 12633 22624
rect 12575 22593 12587 22596
rect 12529 22587 12587 22593
rect 12621 22593 12633 22596
rect 12667 22593 12679 22627
rect 12621 22587 12679 22593
rect 12894 22584 12900 22636
rect 12952 22584 12958 22636
rect 11241 22559 11299 22565
rect 11241 22556 11253 22559
rect 10060 22528 11253 22556
rect 9769 22519 9827 22525
rect 11241 22525 11253 22528
rect 11287 22525 11299 22559
rect 11241 22519 11299 22525
rect 11606 22516 11612 22568
rect 11664 22516 11670 22568
rect 11885 22559 11943 22565
rect 11885 22556 11897 22559
rect 11716 22528 11897 22556
rect 9677 22491 9735 22497
rect 9677 22457 9689 22491
rect 9723 22488 9735 22491
rect 10134 22488 10140 22500
rect 9723 22460 10140 22488
rect 9723 22457 9735 22460
rect 9677 22451 9735 22457
rect 10134 22448 10140 22460
rect 10192 22488 10198 22500
rect 10505 22491 10563 22497
rect 10505 22488 10517 22491
rect 10192 22460 10517 22488
rect 10192 22448 10198 22460
rect 10505 22457 10517 22460
rect 10551 22488 10563 22491
rect 11716 22488 11744 22528
rect 11885 22525 11897 22528
rect 11931 22556 11943 22559
rect 12158 22556 12164 22568
rect 11931 22528 12164 22556
rect 11931 22525 11943 22528
rect 11885 22519 11943 22525
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 12713 22559 12771 22565
rect 12713 22556 12725 22559
rect 12406 22528 12725 22556
rect 10551 22460 11744 22488
rect 11793 22491 11851 22497
rect 10551 22457 10563 22460
rect 10505 22451 10563 22457
rect 11793 22457 11805 22491
rect 11839 22488 11851 22491
rect 12406 22488 12434 22528
rect 12713 22525 12725 22528
rect 12759 22525 12771 22559
rect 12713 22519 12771 22525
rect 11839 22460 12434 22488
rect 11839 22457 11851 22460
rect 11793 22451 11851 22457
rect 12894 22380 12900 22432
rect 12952 22380 12958 22432
rect 13648 22420 13676 22664
rect 14378 22661 14390 22664
rect 14424 22661 14436 22695
rect 14378 22655 14436 22661
rect 14550 22584 14556 22636
rect 14608 22624 14614 22636
rect 14645 22627 14703 22633
rect 14645 22624 14657 22627
rect 14608 22596 14657 22624
rect 14608 22584 14614 22596
rect 14645 22593 14657 22596
rect 14691 22593 14703 22627
rect 14645 22587 14703 22593
rect 14844 22556 14872 22720
rect 15028 22633 15056 22720
rect 15841 22695 15899 22701
rect 15841 22692 15853 22695
rect 15212 22664 15853 22692
rect 15212 22633 15240 22664
rect 15841 22661 15853 22664
rect 15887 22661 15899 22695
rect 16666 22692 16672 22704
rect 15841 22655 15899 22661
rect 16408 22664 16672 22692
rect 15013 22627 15071 22633
rect 15013 22593 15025 22627
rect 15059 22593 15071 22627
rect 15013 22587 15071 22593
rect 15197 22627 15255 22633
rect 15197 22593 15209 22627
rect 15243 22593 15255 22627
rect 15197 22587 15255 22593
rect 15470 22584 15476 22636
rect 15528 22624 15534 22636
rect 15749 22627 15807 22633
rect 15528 22596 15700 22624
rect 15528 22584 15534 22596
rect 15105 22559 15163 22565
rect 15105 22556 15117 22559
rect 14844 22528 15117 22556
rect 15105 22525 15117 22528
rect 15151 22525 15163 22559
rect 15672 22556 15700 22596
rect 15749 22593 15761 22627
rect 15795 22624 15807 22627
rect 16408 22624 16436 22664
rect 16666 22652 16672 22664
rect 16724 22652 16730 22704
rect 15795 22596 16436 22624
rect 16485 22627 16543 22633
rect 15795 22593 15807 22596
rect 15749 22587 15807 22593
rect 16485 22593 16497 22627
rect 16531 22624 16543 22627
rect 17144 22624 17172 22720
rect 18509 22695 18567 22701
rect 16531 22596 17172 22624
rect 17236 22664 17724 22692
rect 16531 22593 16543 22596
rect 16485 22587 16543 22593
rect 17236 22556 17264 22664
rect 17586 22584 17592 22636
rect 17644 22584 17650 22636
rect 17696 22633 17724 22664
rect 18509 22661 18521 22695
rect 18555 22692 18567 22695
rect 19058 22692 19064 22704
rect 18555 22664 19064 22692
rect 18555 22661 18567 22664
rect 18509 22655 18567 22661
rect 19058 22652 19064 22664
rect 19116 22652 19122 22704
rect 19168 22664 22094 22692
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22593 17739 22627
rect 17681 22587 17739 22593
rect 17865 22627 17923 22633
rect 17865 22593 17877 22627
rect 17911 22593 17923 22627
rect 17865 22587 17923 22593
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22624 18107 22627
rect 19168 22624 19196 22664
rect 18095 22596 19196 22624
rect 18095 22593 18107 22596
rect 18049 22587 18107 22593
rect 15672 22528 17264 22556
rect 17313 22559 17371 22565
rect 15105 22519 15163 22525
rect 17313 22525 17325 22559
rect 17359 22556 17371 22559
rect 17405 22559 17463 22565
rect 17405 22556 17417 22559
rect 17359 22528 17417 22556
rect 17359 22525 17371 22528
rect 17313 22519 17371 22525
rect 17405 22525 17417 22528
rect 17451 22525 17463 22559
rect 17880 22556 17908 22587
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 19484 22596 20024 22624
rect 19484 22584 19490 22596
rect 17405 22519 17463 22525
rect 17604 22528 17908 22556
rect 15381 22491 15439 22497
rect 15381 22457 15393 22491
rect 15427 22457 15439 22491
rect 15381 22451 15439 22457
rect 15657 22491 15715 22497
rect 15657 22457 15669 22491
rect 15703 22488 15715 22491
rect 17604 22488 17632 22528
rect 19702 22516 19708 22568
rect 19760 22516 19766 22568
rect 19996 22556 20024 22596
rect 20070 22584 20076 22636
rect 20128 22624 20134 22636
rect 20533 22627 20591 22633
rect 20533 22624 20545 22627
rect 20128 22596 20545 22624
rect 20128 22584 20134 22596
rect 20533 22593 20545 22596
rect 20579 22593 20591 22627
rect 20533 22587 20591 22593
rect 20714 22584 20720 22636
rect 20772 22584 20778 22636
rect 21082 22584 21088 22636
rect 21140 22624 21146 22636
rect 21269 22627 21327 22633
rect 21269 22624 21281 22627
rect 21140 22596 21281 22624
rect 21140 22584 21146 22596
rect 21269 22593 21281 22596
rect 21315 22624 21327 22627
rect 21726 22624 21732 22636
rect 21315 22596 21732 22624
rect 21315 22593 21327 22596
rect 21269 22587 21327 22593
rect 21726 22584 21732 22596
rect 21784 22584 21790 22636
rect 22066 22624 22094 22664
rect 23014 22652 23020 22704
rect 23072 22701 23078 22704
rect 23072 22695 23095 22701
rect 23083 22661 23095 22695
rect 23308 22692 23336 22720
rect 23308 22664 23612 22692
rect 23072 22655 23095 22661
rect 23072 22652 23078 22655
rect 23198 22624 23204 22636
rect 22066 22596 23204 22624
rect 23198 22584 23204 22596
rect 23256 22624 23262 22636
rect 23584 22633 23612 22664
rect 23768 22633 23796 22732
rect 23842 22720 23848 22772
rect 23900 22720 23906 22772
rect 24029 22763 24087 22769
rect 24029 22729 24041 22763
rect 24075 22760 24087 22763
rect 24118 22760 24124 22772
rect 24075 22732 24124 22760
rect 24075 22729 24087 22732
rect 24029 22723 24087 22729
rect 24118 22720 24124 22732
rect 24176 22720 24182 22772
rect 24302 22720 24308 22772
rect 24360 22760 24366 22772
rect 25130 22760 25136 22772
rect 24360 22732 25136 22760
rect 24360 22720 24366 22732
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 28261 22763 28319 22769
rect 25976 22732 26832 22760
rect 23860 22692 23888 22720
rect 24762 22692 24768 22704
rect 23860 22664 24768 22692
rect 24762 22652 24768 22664
rect 24820 22692 24826 22704
rect 25976 22692 26004 22732
rect 24820 22664 26004 22692
rect 24820 22652 24826 22664
rect 26050 22652 26056 22704
rect 26108 22652 26114 22704
rect 26804 22701 26832 22732
rect 28261 22729 28273 22763
rect 28307 22760 28319 22763
rect 28350 22760 28356 22772
rect 28307 22732 28356 22760
rect 28307 22729 28319 22732
rect 28261 22723 28319 22729
rect 28350 22720 28356 22732
rect 28408 22720 28414 22772
rect 29362 22720 29368 22772
rect 29420 22720 29426 22772
rect 30650 22760 30656 22772
rect 29656 22732 30656 22760
rect 26789 22695 26847 22701
rect 26789 22661 26801 22695
rect 26835 22692 26847 22695
rect 27893 22695 27951 22701
rect 27893 22692 27905 22695
rect 26835 22664 27905 22692
rect 26835 22661 26847 22664
rect 26789 22655 26847 22661
rect 27893 22661 27905 22664
rect 27939 22692 27951 22695
rect 27939 22664 29224 22692
rect 27939 22661 27951 22664
rect 27893 22655 27951 22661
rect 23385 22627 23443 22633
rect 23385 22624 23397 22627
rect 23256 22596 23397 22624
rect 23256 22584 23262 22596
rect 23385 22593 23397 22596
rect 23431 22593 23443 22627
rect 23385 22587 23443 22593
rect 23569 22627 23627 22633
rect 23569 22593 23581 22627
rect 23615 22593 23627 22627
rect 23569 22587 23627 22593
rect 23753 22627 23811 22633
rect 23753 22593 23765 22627
rect 23799 22593 23811 22627
rect 23753 22587 23811 22593
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22624 23903 22627
rect 24210 22624 24216 22636
rect 23891 22596 24216 22624
rect 23891 22593 23903 22596
rect 23845 22587 23903 22593
rect 24210 22584 24216 22596
rect 24268 22584 24274 22636
rect 24670 22584 24676 22636
rect 24728 22584 24734 22636
rect 25429 22627 25487 22633
rect 25429 22593 25441 22627
rect 25475 22624 25487 22627
rect 25685 22627 25743 22633
rect 25475 22596 25636 22624
rect 25475 22593 25487 22596
rect 25429 22587 25487 22593
rect 20898 22556 20904 22568
rect 19996 22528 20904 22556
rect 20898 22516 20904 22528
rect 20956 22516 20962 22568
rect 23293 22559 23351 22565
rect 23293 22525 23305 22559
rect 23339 22556 23351 22559
rect 24688 22556 24716 22584
rect 23339 22528 24716 22556
rect 25608 22556 25636 22596
rect 25685 22593 25697 22627
rect 25731 22624 25743 22627
rect 26068 22624 26096 22652
rect 27065 22627 27123 22633
rect 27065 22624 27077 22627
rect 25731 22596 27077 22624
rect 25731 22593 25743 22596
rect 25685 22587 25743 22593
rect 27065 22593 27077 22596
rect 27111 22624 27123 22627
rect 29086 22624 29092 22636
rect 27111 22596 29092 22624
rect 27111 22593 27123 22596
rect 27065 22587 27123 22593
rect 29086 22584 29092 22596
rect 29144 22584 29150 22636
rect 26053 22559 26111 22565
rect 25608 22528 26004 22556
rect 23339 22525 23351 22528
rect 23293 22519 23351 22525
rect 15703 22460 17632 22488
rect 17773 22491 17831 22497
rect 15703 22457 15715 22460
rect 15657 22451 15715 22457
rect 17773 22457 17785 22491
rect 17819 22457 17831 22491
rect 17773 22451 17831 22457
rect 15396 22420 15424 22451
rect 13648 22392 15424 22420
rect 16666 22380 16672 22432
rect 16724 22380 16730 22432
rect 16942 22380 16948 22432
rect 17000 22420 17006 22432
rect 17788 22420 17816 22451
rect 23658 22448 23664 22500
rect 23716 22448 23722 22500
rect 25976 22488 26004 22528
rect 26053 22525 26065 22559
rect 26099 22556 26111 22559
rect 26326 22556 26332 22568
rect 26099 22528 26332 22556
rect 26099 22525 26111 22528
rect 26053 22519 26111 22525
rect 26326 22516 26332 22528
rect 26384 22516 26390 22568
rect 28810 22516 28816 22568
rect 28868 22516 28874 22568
rect 29196 22556 29224 22664
rect 29270 22584 29276 22636
rect 29328 22624 29334 22636
rect 29656 22633 29684 22732
rect 30650 22720 30656 22732
rect 30708 22720 30714 22772
rect 31757 22763 31815 22769
rect 31757 22729 31769 22763
rect 31803 22760 31815 22763
rect 32214 22760 32220 22772
rect 31803 22732 32220 22760
rect 31803 22729 31815 22732
rect 31757 22723 31815 22729
rect 32214 22720 32220 22732
rect 32272 22720 32278 22772
rect 34238 22760 34244 22772
rect 32324 22732 34244 22760
rect 29748 22664 31754 22692
rect 29549 22627 29607 22633
rect 29549 22624 29561 22627
rect 29328 22596 29561 22624
rect 29328 22584 29334 22596
rect 29549 22593 29561 22596
rect 29595 22593 29607 22627
rect 29549 22587 29607 22593
rect 29641 22627 29699 22633
rect 29641 22593 29653 22627
rect 29687 22593 29699 22627
rect 29641 22587 29699 22593
rect 29748 22556 29776 22664
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22593 29883 22627
rect 29825 22587 29883 22593
rect 29917 22627 29975 22633
rect 29917 22593 29929 22627
rect 29963 22624 29975 22627
rect 30466 22624 30472 22636
rect 29963 22596 30472 22624
rect 29963 22593 29975 22596
rect 29917 22587 29975 22593
rect 29196 22528 29776 22556
rect 26418 22488 26424 22500
rect 25976 22460 26424 22488
rect 26418 22448 26424 22460
rect 26476 22448 26482 22500
rect 17000 22392 17816 22420
rect 20625 22423 20683 22429
rect 17000 22380 17006 22392
rect 20625 22389 20637 22423
rect 20671 22420 20683 22423
rect 20714 22420 20720 22432
rect 20671 22392 20720 22420
rect 20671 22389 20683 22392
rect 20625 22383 20683 22389
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 21358 22380 21364 22432
rect 21416 22380 21422 22432
rect 25498 22380 25504 22432
rect 25556 22420 25562 22432
rect 29840 22420 29868 22587
rect 30466 22584 30472 22596
rect 30524 22584 30530 22636
rect 30644 22627 30702 22633
rect 30644 22593 30656 22627
rect 30690 22624 30702 22627
rect 31018 22624 31024 22636
rect 30690 22596 31024 22624
rect 30690 22593 30702 22596
rect 30644 22587 30702 22593
rect 31018 22584 31024 22596
rect 31076 22584 31082 22636
rect 30374 22516 30380 22568
rect 30432 22516 30438 22568
rect 31726 22556 31754 22664
rect 32324 22633 32352 22732
rect 34238 22720 34244 22732
rect 34296 22720 34302 22772
rect 36078 22720 36084 22772
rect 36136 22760 36142 22772
rect 37277 22763 37335 22769
rect 37277 22760 37289 22763
rect 36136 22732 37289 22760
rect 36136 22720 36142 22732
rect 37277 22729 37289 22732
rect 37323 22729 37335 22763
rect 37277 22723 37335 22729
rect 38378 22720 38384 22772
rect 38436 22720 38442 22772
rect 33597 22695 33655 22701
rect 33597 22661 33609 22695
rect 33643 22692 33655 22695
rect 33870 22692 33876 22704
rect 33643 22664 33876 22692
rect 33643 22661 33655 22664
rect 33597 22655 33655 22661
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22593 32367 22627
rect 32769 22627 32827 22633
rect 32769 22624 32781 22627
rect 32309 22587 32367 22593
rect 32416 22596 32781 22624
rect 32416 22556 32444 22596
rect 32769 22593 32781 22596
rect 32815 22624 32827 22627
rect 33318 22624 33324 22636
rect 32815 22596 33324 22624
rect 32815 22593 32827 22596
rect 32769 22587 32827 22593
rect 33318 22584 33324 22596
rect 33376 22584 33382 22636
rect 33796 22633 33824 22664
rect 33870 22652 33876 22664
rect 33928 22692 33934 22704
rect 34330 22692 34336 22704
rect 33928 22664 34336 22692
rect 33928 22652 33934 22664
rect 34330 22652 34336 22664
rect 34388 22652 34394 22704
rect 36417 22695 36475 22701
rect 36417 22692 36429 22695
rect 35820 22664 36429 22692
rect 33781 22627 33839 22633
rect 33781 22593 33793 22627
rect 33827 22624 33839 22627
rect 34048 22627 34106 22633
rect 33827 22596 33861 22624
rect 33827 22593 33839 22596
rect 33781 22587 33839 22593
rect 34048 22593 34060 22627
rect 34094 22624 34106 22627
rect 34514 22624 34520 22636
rect 34094 22596 34520 22624
rect 34094 22593 34106 22596
rect 34048 22587 34106 22593
rect 34514 22584 34520 22596
rect 34572 22584 34578 22636
rect 31726 22528 32444 22556
rect 32585 22559 32643 22565
rect 32585 22525 32597 22559
rect 32631 22556 32643 22559
rect 32950 22556 32956 22568
rect 32631 22528 32956 22556
rect 32631 22525 32643 22528
rect 32585 22519 32643 22525
rect 32950 22516 32956 22528
rect 33008 22516 33014 22568
rect 35618 22516 35624 22568
rect 35676 22556 35682 22568
rect 35820 22565 35848 22664
rect 36417 22661 36429 22664
rect 36463 22661 36475 22695
rect 36417 22655 36475 22661
rect 36633 22695 36691 22701
rect 36633 22661 36645 22695
rect 36679 22692 36691 22695
rect 38010 22692 38016 22704
rect 36679 22664 38016 22692
rect 36679 22661 36691 22664
rect 36633 22655 36691 22661
rect 38010 22652 38016 22664
rect 38068 22652 38074 22704
rect 37921 22627 37979 22633
rect 37921 22593 37933 22627
rect 37967 22624 37979 22627
rect 38396 22624 38424 22720
rect 37967 22596 38424 22624
rect 37967 22593 37979 22596
rect 37921 22587 37979 22593
rect 35805 22559 35863 22565
rect 35805 22556 35817 22559
rect 35676 22528 35817 22556
rect 35676 22516 35682 22528
rect 35805 22525 35817 22528
rect 35851 22525 35863 22559
rect 35805 22519 35863 22525
rect 35161 22491 35219 22497
rect 31726 22460 32628 22488
rect 31726 22420 31754 22460
rect 32600 22432 32628 22460
rect 35161 22457 35173 22491
rect 35207 22488 35219 22491
rect 35342 22488 35348 22500
rect 35207 22460 35348 22488
rect 35207 22457 35219 22460
rect 35161 22451 35219 22457
rect 35342 22448 35348 22460
rect 35400 22488 35406 22500
rect 35636 22488 35664 22516
rect 37936 22488 37964 22587
rect 35400 22460 35664 22488
rect 36464 22460 37964 22488
rect 35400 22448 35406 22460
rect 25556 22392 31754 22420
rect 25556 22380 25562 22392
rect 32122 22380 32128 22432
rect 32180 22380 32186 22432
rect 32398 22380 32404 22432
rect 32456 22420 32462 22432
rect 32493 22423 32551 22429
rect 32493 22420 32505 22423
rect 32456 22392 32505 22420
rect 32456 22380 32462 22392
rect 32493 22389 32505 22392
rect 32539 22389 32551 22423
rect 32493 22383 32551 22389
rect 32582 22380 32588 22432
rect 32640 22380 32646 22432
rect 35250 22380 35256 22432
rect 35308 22380 35314 22432
rect 35986 22380 35992 22432
rect 36044 22420 36050 22432
rect 36464 22429 36492 22460
rect 36265 22423 36323 22429
rect 36265 22420 36277 22423
rect 36044 22392 36277 22420
rect 36044 22380 36050 22392
rect 36265 22389 36277 22392
rect 36311 22389 36323 22423
rect 36265 22383 36323 22389
rect 36449 22423 36507 22429
rect 36449 22389 36461 22423
rect 36495 22389 36507 22423
rect 36449 22383 36507 22389
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 8938 22176 8944 22228
rect 8996 22216 9002 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 8996 22188 9045 22216
rect 8996 22176 9002 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9033 22179 9091 22185
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10229 22219 10287 22225
rect 10229 22216 10241 22219
rect 10008 22188 10241 22216
rect 10008 22176 10014 22188
rect 10229 22185 10241 22188
rect 10275 22185 10287 22219
rect 10229 22179 10287 22185
rect 12158 22176 12164 22228
rect 12216 22216 12222 22228
rect 12621 22219 12679 22225
rect 12621 22216 12633 22219
rect 12216 22188 12633 22216
rect 12216 22176 12222 22188
rect 12621 22185 12633 22188
rect 12667 22185 12679 22219
rect 12894 22216 12900 22228
rect 12621 22179 12679 22185
rect 12728 22188 12900 22216
rect 10689 22083 10747 22089
rect 10689 22049 10701 22083
rect 10735 22080 10747 22083
rect 12176 22080 12204 22176
rect 12434 22108 12440 22160
rect 12492 22148 12498 22160
rect 12728 22148 12756 22188
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 15470 22176 15476 22228
rect 15528 22176 15534 22228
rect 16942 22176 16948 22228
rect 17000 22176 17006 22228
rect 19058 22176 19064 22228
rect 19116 22216 19122 22228
rect 19242 22216 19248 22228
rect 19116 22188 19248 22216
rect 19116 22176 19122 22188
rect 19242 22176 19248 22188
rect 19300 22176 19306 22228
rect 19702 22176 19708 22228
rect 19760 22216 19766 22228
rect 25498 22216 25504 22228
rect 19760 22188 25504 22216
rect 19760 22176 19766 22188
rect 25498 22176 25504 22188
rect 25556 22176 25562 22228
rect 26418 22176 26424 22228
rect 26476 22176 26482 22228
rect 29362 22216 29368 22228
rect 28460 22188 29368 22216
rect 12492 22120 12756 22148
rect 12492 22108 12498 22120
rect 13078 22108 13084 22160
rect 13136 22148 13142 22160
rect 13173 22151 13231 22157
rect 13173 22148 13185 22151
rect 13136 22120 13185 22148
rect 13136 22108 13142 22120
rect 13173 22117 13185 22120
rect 13219 22117 13231 22151
rect 13173 22111 13231 22117
rect 18782 22108 18788 22160
rect 18840 22148 18846 22160
rect 19720 22148 19748 22176
rect 18840 22120 19748 22148
rect 18840 22108 18846 22120
rect 22830 22108 22836 22160
rect 22888 22148 22894 22160
rect 23017 22151 23075 22157
rect 23017 22148 23029 22151
rect 22888 22120 23029 22148
rect 22888 22108 22894 22120
rect 23017 22117 23029 22120
rect 23063 22148 23075 22151
rect 24213 22151 24271 22157
rect 23063 22120 23980 22148
rect 23063 22117 23075 22120
rect 23017 22111 23075 22117
rect 10735 22052 12204 22080
rect 12805 22083 12863 22089
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 12805 22049 12817 22083
rect 12851 22080 12863 22083
rect 12851 22052 13216 22080
rect 12851 22049 12863 22052
rect 12805 22043 12863 22049
rect 8846 21972 8852 22024
rect 8904 22012 8910 22024
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8904 21984 8953 22012
rect 8904 21972 8910 21984
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 10428 21944 10456 21975
rect 10502 21972 10508 22024
rect 10560 21972 10566 22024
rect 10594 21972 10600 22024
rect 10652 21972 10658 22024
rect 10870 21972 10876 22024
rect 10928 21972 10934 22024
rect 12526 21972 12532 22024
rect 12584 22012 12590 22024
rect 12621 22015 12679 22021
rect 12621 22012 12633 22015
rect 12584 21984 12633 22012
rect 12584 21972 12590 21984
rect 12621 21981 12633 21984
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 21981 12955 22015
rect 12897 21975 12955 21981
rect 10888 21944 10916 21972
rect 10428 21916 10916 21944
rect 11698 21904 11704 21956
rect 11756 21944 11762 21956
rect 12912 21944 12940 21975
rect 11756 21916 12940 21944
rect 13188 21944 13216 22052
rect 13354 22040 13360 22092
rect 13412 22080 13418 22092
rect 13725 22083 13783 22089
rect 13725 22080 13737 22083
rect 13412 22052 13737 22080
rect 13412 22040 13418 22052
rect 13725 22049 13737 22052
rect 13771 22049 13783 22083
rect 13725 22043 13783 22049
rect 15194 22040 15200 22092
rect 15252 22040 15258 22092
rect 16853 22083 16911 22089
rect 16853 22049 16865 22083
rect 16899 22080 16911 22083
rect 19242 22080 19248 22092
rect 16899 22052 19248 22080
rect 16899 22049 16911 22052
rect 16853 22043 16911 22049
rect 19242 22040 19248 22052
rect 19300 22040 19306 22092
rect 23842 22080 23848 22092
rect 20180 22052 23848 22080
rect 13262 21972 13268 22024
rect 13320 22012 13326 22024
rect 13541 22015 13599 22021
rect 13541 22012 13553 22015
rect 13320 21984 13553 22012
rect 13320 21972 13326 21984
rect 13541 21981 13553 21984
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 13633 22015 13691 22021
rect 13633 21981 13645 22015
rect 13679 22012 13691 22015
rect 15212 22012 15240 22040
rect 13679 21984 15240 22012
rect 13679 21981 13691 21984
rect 13633 21975 13691 21981
rect 16574 21972 16580 22024
rect 16632 22021 16638 22024
rect 16632 21975 16644 22021
rect 16632 21972 16638 21975
rect 17586 21972 17592 22024
rect 17644 21972 17650 22024
rect 17865 22015 17923 22021
rect 17865 21981 17877 22015
rect 17911 21981 17923 22015
rect 17865 21975 17923 21981
rect 17957 22015 18015 22021
rect 17957 21981 17969 22015
rect 18003 22012 18015 22015
rect 18046 22012 18052 22024
rect 18003 21984 18052 22012
rect 18003 21981 18015 21984
rect 17957 21975 18015 21981
rect 13188 21916 14044 21944
rect 11756 21904 11762 21916
rect 14016 21888 14044 21916
rect 10502 21836 10508 21888
rect 10560 21876 10566 21888
rect 11146 21876 11152 21888
rect 10560 21848 11152 21876
rect 10560 21836 10566 21848
rect 11146 21836 11152 21848
rect 11204 21836 11210 21888
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 12434 21876 12440 21888
rect 12032 21848 12440 21876
rect 12032 21836 12038 21848
rect 12434 21836 12440 21848
rect 12492 21836 12498 21888
rect 13081 21879 13139 21885
rect 13081 21845 13093 21879
rect 13127 21876 13139 21879
rect 13538 21876 13544 21888
rect 13127 21848 13544 21876
rect 13127 21845 13139 21848
rect 13081 21839 13139 21845
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 13998 21836 14004 21888
rect 14056 21836 14062 21888
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 17880 21876 17908 21975
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18141 22015 18199 22021
rect 18141 21981 18153 22015
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 17954 21876 17960 21888
rect 17880 21848 17960 21876
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 18156 21876 18184 21975
rect 18248 21944 18276 21975
rect 18414 21972 18420 22024
rect 18472 21972 18478 22024
rect 20180 22012 20208 22052
rect 23842 22040 23848 22052
rect 23900 22040 23906 22092
rect 23952 22031 23980 22120
rect 24213 22117 24225 22151
rect 24259 22148 24271 22151
rect 24673 22151 24731 22157
rect 24259 22120 24624 22148
rect 24259 22117 24271 22120
rect 24213 22111 24271 22117
rect 24596 22080 24624 22120
rect 24673 22117 24685 22151
rect 24719 22148 24731 22151
rect 24719 22120 24900 22148
rect 24719 22117 24731 22120
rect 24673 22111 24731 22117
rect 24765 22083 24823 22089
rect 24765 22080 24777 22083
rect 24596 22052 24777 22080
rect 24765 22049 24777 22052
rect 24811 22049 24823 22083
rect 24765 22043 24823 22049
rect 23937 22025 23995 22031
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 19260 21984 20208 22012
rect 20272 21984 20361 22012
rect 18248 21916 19104 21944
rect 19076 21888 19104 21916
rect 19150 21904 19156 21956
rect 19208 21944 19214 21956
rect 19260 21953 19288 21984
rect 20272 21956 20300 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 20714 21972 20720 22024
rect 20772 21972 20778 22024
rect 23017 22015 23075 22021
rect 23017 22012 23029 22015
rect 22848 21984 23029 22012
rect 22848 21956 22876 21984
rect 23017 21981 23029 21984
rect 23063 21981 23075 22015
rect 23017 21975 23075 21981
rect 23106 21972 23112 22024
rect 23164 21972 23170 22024
rect 23937 21991 23949 22025
rect 23983 21991 23995 22025
rect 23937 21985 23995 21991
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 22012 24087 22015
rect 24302 22012 24308 22024
rect 24075 21984 24308 22012
rect 24075 21981 24087 21984
rect 24029 21975 24087 21981
rect 24302 21972 24308 21984
rect 24360 21972 24366 22024
rect 24394 21972 24400 22024
rect 24452 21972 24458 22024
rect 24872 22012 24900 22120
rect 26878 22108 26884 22160
rect 26936 22108 26942 22160
rect 28460 22148 28488 22188
rect 29362 22176 29368 22188
rect 29420 22176 29426 22228
rect 31202 22176 31208 22228
rect 31260 22176 31266 22228
rect 32490 22216 32496 22228
rect 31772 22188 32496 22216
rect 28368 22120 28488 22148
rect 25409 22083 25467 22089
rect 25409 22049 25421 22083
rect 25455 22080 25467 22083
rect 26896 22080 26924 22108
rect 25455 22052 26464 22080
rect 25455 22049 25467 22052
rect 25409 22043 25467 22049
rect 26436 22021 26464 22052
rect 26703 22052 26924 22080
rect 27065 22083 27123 22089
rect 26237 22015 26295 22021
rect 26237 22012 26249 22015
rect 24872 21984 26249 22012
rect 26237 21981 26249 21984
rect 26283 21981 26295 22015
rect 26237 21975 26295 21981
rect 26421 22015 26479 22021
rect 26421 21981 26433 22015
rect 26467 21981 26479 22015
rect 26421 21975 26479 21981
rect 26617 22015 26675 22021
rect 26617 21981 26629 22015
rect 26663 22012 26675 22015
rect 26703 22012 26731 22052
rect 27065 22049 27077 22083
rect 27111 22080 27123 22083
rect 28368 22080 28396 22120
rect 27111 22052 28396 22080
rect 29365 22083 29423 22089
rect 27111 22049 27123 22052
rect 27065 22043 27123 22049
rect 29365 22049 29377 22083
rect 29411 22080 29423 22083
rect 30374 22080 30380 22092
rect 29411 22052 30380 22080
rect 29411 22049 29423 22052
rect 29365 22043 29423 22049
rect 30374 22040 30380 22052
rect 30432 22040 30438 22092
rect 31220 22080 31248 22176
rect 31665 22083 31723 22089
rect 31665 22080 31677 22083
rect 31220 22052 31677 22080
rect 31665 22049 31677 22052
rect 31711 22049 31723 22083
rect 31665 22043 31723 22049
rect 26663 21984 26731 22012
rect 26881 22015 26939 22021
rect 26663 21981 26675 21984
rect 26617 21975 26675 21981
rect 26881 21981 26893 22015
rect 26927 21981 26939 22015
rect 26881 21975 26939 21981
rect 27157 22015 27215 22021
rect 27157 21981 27169 22015
rect 27203 22012 27215 22015
rect 27203 21984 27292 22012
rect 27203 21981 27215 21984
rect 27157 21975 27215 21981
rect 19245 21947 19303 21953
rect 19245 21944 19257 21947
rect 19208 21916 19257 21944
rect 19208 21904 19214 21916
rect 19245 21913 19257 21916
rect 19291 21913 19303 21947
rect 19245 21907 19303 21913
rect 20073 21947 20131 21953
rect 20073 21913 20085 21947
rect 20119 21944 20131 21947
rect 20254 21944 20260 21956
rect 20119 21916 20260 21944
rect 20119 21913 20131 21916
rect 20073 21907 20131 21913
rect 20254 21904 20260 21916
rect 20312 21904 20318 21956
rect 21266 21904 21272 21956
rect 21324 21904 21330 21956
rect 22830 21904 22836 21956
rect 22888 21904 22894 21956
rect 23293 21947 23351 21953
rect 23293 21913 23305 21947
rect 23339 21944 23351 21947
rect 23382 21944 23388 21956
rect 23339 21916 23388 21944
rect 23339 21913 23351 21916
rect 23293 21907 23351 21913
rect 23382 21904 23388 21916
rect 23440 21904 23446 21956
rect 24210 21904 24216 21956
rect 24268 21904 24274 21956
rect 24670 21904 24676 21956
rect 24728 21904 24734 21956
rect 18690 21876 18696 21888
rect 18156 21848 18696 21876
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 19058 21836 19064 21888
rect 19116 21836 19122 21888
rect 22094 21836 22100 21888
rect 22152 21885 22158 21888
rect 22152 21879 22201 21885
rect 22152 21845 22155 21879
rect 22189 21845 22201 21879
rect 22152 21839 22201 21845
rect 22152 21836 22158 21839
rect 24486 21836 24492 21888
rect 24544 21836 24550 21888
rect 25682 21836 25688 21888
rect 25740 21836 25746 21888
rect 26694 21836 26700 21888
rect 26752 21836 26758 21888
rect 26896 21876 26924 21975
rect 27264 21953 27292 21984
rect 27798 21972 27804 22024
rect 27856 21972 27862 22024
rect 28166 21972 28172 22024
rect 28224 21972 28230 22024
rect 31772 22021 31800 22188
rect 32490 22176 32496 22188
rect 32548 22176 32554 22228
rect 33226 22176 33232 22228
rect 33284 22176 33290 22228
rect 35989 22219 36047 22225
rect 33888 22188 35940 22216
rect 33888 22160 33916 22188
rect 33870 22108 33876 22160
rect 33928 22108 33934 22160
rect 34514 22108 34520 22160
rect 34572 22148 34578 22160
rect 34701 22151 34759 22157
rect 34701 22148 34713 22151
rect 34572 22120 34713 22148
rect 34572 22108 34578 22120
rect 34701 22117 34713 22120
rect 34747 22117 34759 22151
rect 34701 22111 34759 22117
rect 34790 22108 34796 22160
rect 34848 22148 34854 22160
rect 35253 22151 35311 22157
rect 35253 22148 35265 22151
rect 34848 22120 35265 22148
rect 34848 22108 34854 22120
rect 35253 22117 35265 22120
rect 35299 22148 35311 22151
rect 35526 22148 35532 22160
rect 35299 22120 35532 22148
rect 35299 22117 35311 22120
rect 35253 22111 35311 22117
rect 35526 22108 35532 22120
rect 35584 22108 35590 22160
rect 35912 22148 35940 22188
rect 35989 22185 36001 22219
rect 36035 22216 36047 22219
rect 36170 22216 36176 22228
rect 36035 22188 36176 22216
rect 36035 22185 36047 22188
rect 35989 22179 36047 22185
rect 36170 22176 36176 22188
rect 36228 22176 36234 22228
rect 38010 22216 38016 22228
rect 36372 22188 36676 22216
rect 37971 22188 38016 22216
rect 36372 22148 36400 22188
rect 35912 22120 36400 22148
rect 36449 22151 36507 22157
rect 36449 22117 36461 22151
rect 36495 22148 36507 22151
rect 36538 22148 36544 22160
rect 36495 22120 36544 22148
rect 36495 22117 36507 22120
rect 36449 22111 36507 22117
rect 36538 22108 36544 22120
rect 36596 22108 36602 22160
rect 36648 22092 36676 22188
rect 38010 22176 38016 22188
rect 38068 22176 38074 22228
rect 34422 22080 34428 22092
rect 34348 22052 34428 22080
rect 31573 22015 31631 22021
rect 31573 21981 31585 22015
rect 31619 21981 31631 22015
rect 31573 21975 31631 21981
rect 31757 22015 31815 22021
rect 31757 21981 31769 22015
rect 31803 21981 31815 22015
rect 31757 21975 31815 21981
rect 31849 22015 31907 22021
rect 31849 21981 31861 22015
rect 31895 22012 31907 22015
rect 31895 21984 33088 22012
rect 31895 21981 31907 21984
rect 31849 21975 31907 21981
rect 27249 21947 27307 21953
rect 27249 21913 27261 21947
rect 27295 21944 27307 21947
rect 28184 21944 28212 21972
rect 27295 21916 28212 21944
rect 29120 21947 29178 21953
rect 27295 21913 27307 21916
rect 27249 21907 27307 21913
rect 29120 21913 29132 21947
rect 29166 21944 29178 21947
rect 29454 21944 29460 21956
rect 29166 21916 29460 21944
rect 29166 21913 29178 21916
rect 29120 21907 29178 21913
rect 29454 21904 29460 21916
rect 29512 21904 29518 21956
rect 27154 21876 27160 21888
rect 26896 21848 27160 21876
rect 27154 21836 27160 21848
rect 27212 21836 27218 21888
rect 27982 21836 27988 21888
rect 28040 21836 28046 21888
rect 28442 21836 28448 21888
rect 28500 21876 28506 21888
rect 31588 21876 31616 21975
rect 33060 21956 33088 21984
rect 33318 21972 33324 22024
rect 33376 21972 33382 22024
rect 34348 22021 34376 22052
rect 34422 22040 34428 22052
rect 34480 22040 34486 22092
rect 35158 22040 35164 22092
rect 35216 22040 35222 22092
rect 35618 22040 35624 22092
rect 35676 22040 35682 22092
rect 35894 22040 35900 22092
rect 35952 22080 35958 22092
rect 36265 22083 36323 22089
rect 36265 22080 36277 22083
rect 35952 22052 36277 22080
rect 35952 22040 35958 22052
rect 36265 22049 36277 22052
rect 36311 22049 36323 22083
rect 36265 22043 36323 22049
rect 36630 22040 36636 22092
rect 36688 22080 36694 22092
rect 38028 22080 38056 22176
rect 38657 22083 38715 22089
rect 38657 22080 38669 22083
rect 36688 22052 36713 22080
rect 38028 22052 38669 22080
rect 36688 22040 36694 22052
rect 38657 22049 38669 22052
rect 38703 22049 38715 22083
rect 38657 22043 38715 22049
rect 34333 22015 34391 22021
rect 34333 21981 34345 22015
rect 34379 21981 34391 22015
rect 34333 21975 34391 21981
rect 34517 22015 34575 22021
rect 34517 21981 34529 22015
rect 34563 22012 34575 22015
rect 34790 22012 34796 22024
rect 34563 21984 34796 22012
rect 34563 21981 34575 21984
rect 34517 21975 34575 21981
rect 32122 21953 32128 21956
rect 32116 21907 32128 21953
rect 32122 21904 32128 21907
rect 32180 21904 32186 21956
rect 33042 21904 33048 21956
rect 33100 21944 33106 21956
rect 34057 21947 34115 21953
rect 34057 21944 34069 21947
rect 33100 21916 34069 21944
rect 33100 21904 33106 21916
rect 34057 21913 34069 21916
rect 34103 21913 34115 21947
rect 34057 21907 34115 21913
rect 31846 21876 31852 21888
rect 28500 21848 31852 21876
rect 28500 21836 28506 21848
rect 31846 21836 31852 21848
rect 31904 21876 31910 21888
rect 34348 21876 34376 21975
rect 34790 21972 34796 21984
rect 34848 21972 34854 22024
rect 34885 22015 34943 22021
rect 34885 21981 34897 22015
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 35069 22015 35127 22021
rect 35069 21981 35081 22015
rect 35115 22012 35127 22015
rect 35434 22012 35440 22024
rect 35115 21984 35440 22012
rect 35115 21981 35127 21984
rect 35069 21975 35127 21981
rect 35392 21978 35440 21984
rect 34425 21947 34483 21953
rect 34425 21913 34437 21947
rect 34471 21944 34483 21947
rect 34900 21944 34928 21975
rect 35434 21972 35440 21978
rect 35492 21972 35498 22024
rect 36541 22015 36599 22021
rect 36541 21981 36553 22015
rect 36587 22012 36599 22015
rect 36722 22012 36728 22024
rect 36587 21984 36728 22012
rect 36587 21981 36599 21984
rect 36541 21975 36599 21981
rect 36722 21972 36728 21984
rect 36780 22012 36786 22024
rect 38105 22015 38163 22021
rect 38105 22012 38117 22015
rect 36780 21984 38117 22012
rect 36780 21972 36786 21984
rect 38105 21981 38117 21984
rect 38151 21981 38163 22015
rect 38105 21975 38163 21981
rect 35434 21969 35492 21972
rect 35986 21953 35992 21956
rect 34471 21916 34928 21944
rect 35973 21947 35992 21953
rect 34471 21913 34483 21916
rect 34425 21907 34483 21913
rect 35973 21913 35985 21947
rect 35973 21907 35992 21913
rect 35986 21904 35992 21907
rect 36044 21904 36050 21956
rect 36906 21953 36912 21956
rect 36173 21947 36231 21953
rect 36173 21913 36185 21947
rect 36219 21944 36231 21947
rect 36219 21916 36768 21944
rect 36219 21913 36231 21916
rect 36173 21907 36231 21913
rect 31904 21848 34376 21876
rect 31904 21836 31910 21848
rect 35802 21836 35808 21888
rect 35860 21836 35866 21888
rect 36262 21836 36268 21888
rect 36320 21836 36326 21888
rect 36740 21876 36768 21916
rect 36900 21907 36912 21953
rect 36906 21904 36912 21907
rect 36964 21904 36970 21956
rect 36814 21876 36820 21888
rect 36740 21848 36820 21876
rect 36814 21836 36820 21848
rect 36872 21836 36878 21888
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 9217 21675 9275 21681
rect 9217 21641 9229 21675
rect 9263 21641 9275 21675
rect 9217 21635 9275 21641
rect 9677 21675 9735 21681
rect 9677 21641 9689 21675
rect 9723 21672 9735 21675
rect 10318 21672 10324 21684
rect 9723 21644 10324 21672
rect 9723 21641 9735 21644
rect 9677 21635 9735 21641
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21536 8723 21539
rect 9232 21536 9260 21635
rect 10318 21632 10324 21644
rect 10376 21672 10382 21684
rect 10778 21672 10784 21684
rect 10376 21644 10784 21672
rect 10376 21632 10382 21644
rect 10778 21632 10784 21644
rect 10836 21672 10842 21684
rect 11974 21672 11980 21684
rect 10836 21644 11284 21672
rect 10836 21632 10842 21644
rect 8711 21508 9260 21536
rect 9585 21539 9643 21545
rect 8711 21505 8723 21508
rect 8665 21499 8723 21505
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9858 21536 9864 21548
rect 9631 21508 9864 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9858 21496 9864 21508
rect 9916 21536 9922 21548
rect 9916 21508 10272 21536
rect 9916 21496 9922 21508
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21437 9827 21471
rect 10244 21468 10272 21508
rect 10870 21496 10876 21548
rect 10928 21536 10934 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10928 21508 10977 21536
rect 10928 21496 10934 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 10965 21499 11023 21505
rect 11146 21496 11152 21548
rect 11204 21496 11210 21548
rect 11256 21536 11284 21644
rect 11808 21644 11980 21672
rect 11808 21613 11836 21644
rect 11974 21632 11980 21644
rect 12032 21632 12038 21684
rect 13906 21632 13912 21684
rect 13964 21672 13970 21684
rect 14918 21672 14924 21684
rect 13964 21644 14924 21672
rect 13964 21632 13970 21644
rect 14918 21632 14924 21644
rect 14976 21632 14982 21684
rect 18325 21675 18383 21681
rect 18325 21641 18337 21675
rect 18371 21672 18383 21675
rect 18414 21672 18420 21684
rect 18371 21644 18420 21672
rect 18371 21641 18383 21644
rect 18325 21635 18383 21641
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 19334 21632 19340 21684
rect 19392 21632 19398 21684
rect 23106 21632 23112 21684
rect 23164 21672 23170 21684
rect 24121 21675 24179 21681
rect 24121 21672 24133 21675
rect 23164 21644 24133 21672
rect 23164 21632 23170 21644
rect 24121 21641 24133 21644
rect 24167 21641 24179 21675
rect 24121 21635 24179 21641
rect 26326 21632 26332 21684
rect 26384 21632 26390 21684
rect 27982 21632 27988 21684
rect 28040 21632 28046 21684
rect 28629 21675 28687 21681
rect 28629 21641 28641 21675
rect 28675 21672 28687 21675
rect 28810 21672 28816 21684
rect 28675 21644 28816 21672
rect 28675 21641 28687 21644
rect 28629 21635 28687 21641
rect 28810 21632 28816 21644
rect 28868 21632 28874 21684
rect 29454 21632 29460 21684
rect 29512 21632 29518 21684
rect 34793 21675 34851 21681
rect 34793 21641 34805 21675
rect 34839 21641 34851 21675
rect 34793 21635 34851 21641
rect 35069 21675 35127 21681
rect 35069 21641 35081 21675
rect 35115 21672 35127 21675
rect 35342 21672 35348 21684
rect 35115 21644 35348 21672
rect 35115 21641 35127 21644
rect 35069 21635 35127 21641
rect 11333 21607 11391 21613
rect 11333 21573 11345 21607
rect 11379 21604 11391 21607
rect 11793 21607 11851 21613
rect 11793 21604 11805 21607
rect 11379 21576 11805 21604
rect 11379 21573 11391 21576
rect 11333 21567 11391 21573
rect 11793 21573 11805 21576
rect 11839 21573 11851 21607
rect 11793 21567 11851 21573
rect 11882 21564 11888 21616
rect 11940 21564 11946 21616
rect 19150 21604 19156 21616
rect 13372 21576 19156 21604
rect 13372 21548 13400 21576
rect 19150 21564 19156 21576
rect 19208 21564 19214 21616
rect 11256 21508 11652 21536
rect 11330 21468 11336 21480
rect 10244 21440 11336 21468
rect 9769 21431 9827 21437
rect 9784 21400 9812 21431
rect 11330 21428 11336 21440
rect 11388 21428 11394 21480
rect 11624 21468 11652 21508
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 12003 21539 12061 21545
rect 12003 21536 12015 21539
rect 11992 21505 12015 21536
rect 12049 21505 12061 21539
rect 11992 21499 12061 21505
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 12250 21536 12256 21548
rect 12207 21508 12256 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 11992 21468 12020 21499
rect 12250 21496 12256 21508
rect 12308 21536 12314 21548
rect 12710 21536 12716 21548
rect 12308 21508 12716 21536
rect 12308 21496 12314 21508
rect 12710 21496 12716 21508
rect 12768 21496 12774 21548
rect 13354 21496 13360 21548
rect 13412 21496 13418 21548
rect 13817 21539 13875 21545
rect 13817 21505 13829 21539
rect 13863 21536 13875 21539
rect 13906 21536 13912 21548
rect 13863 21508 13912 21536
rect 13863 21505 13875 21508
rect 13817 21499 13875 21505
rect 13906 21496 13912 21508
rect 13964 21496 13970 21548
rect 14001 21539 14059 21545
rect 14001 21505 14013 21539
rect 14047 21536 14059 21539
rect 14734 21536 14740 21548
rect 14047 21508 14740 21536
rect 14047 21505 14059 21508
rect 14001 21499 14059 21505
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 17497 21539 17555 21545
rect 17497 21505 17509 21539
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 11624 21440 12020 21468
rect 12621 21471 12679 21477
rect 12621 21437 12633 21471
rect 12667 21468 12679 21471
rect 14090 21468 14096 21480
rect 12667 21440 14096 21468
rect 12667 21437 12679 21440
rect 12621 21431 12679 21437
rect 14090 21428 14096 21440
rect 14148 21428 14154 21480
rect 17512 21468 17540 21499
rect 17678 21496 17684 21548
rect 17736 21496 17742 21548
rect 19352 21536 19380 21632
rect 20898 21564 20904 21616
rect 20956 21604 20962 21616
rect 26234 21604 26240 21616
rect 20956 21576 26240 21604
rect 20956 21564 20962 21576
rect 26234 21564 26240 21576
rect 26292 21564 26298 21616
rect 19438 21539 19496 21545
rect 19438 21536 19450 21539
rect 19352 21508 19450 21536
rect 19438 21505 19450 21508
rect 19484 21505 19496 21539
rect 19438 21499 19496 21505
rect 19705 21539 19763 21545
rect 19705 21505 19717 21539
rect 19751 21505 19763 21539
rect 19705 21499 19763 21505
rect 23477 21539 23535 21545
rect 23477 21505 23489 21539
rect 23523 21536 23535 21539
rect 23934 21536 23940 21548
rect 23523 21508 23940 21536
rect 23523 21505 23535 21508
rect 23477 21499 23535 21505
rect 18046 21468 18052 21480
rect 17512 21440 18052 21468
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 10870 21400 10876 21412
rect 9784 21372 10876 21400
rect 10870 21360 10876 21372
rect 10928 21360 10934 21412
rect 11882 21360 11888 21412
rect 11940 21400 11946 21412
rect 16022 21400 16028 21412
rect 11940 21372 16028 21400
rect 11940 21360 11946 21372
rect 16022 21360 16028 21372
rect 16080 21360 16086 21412
rect 8478 21292 8484 21344
rect 8536 21292 8542 21344
rect 11146 21292 11152 21344
rect 11204 21332 11210 21344
rect 11517 21335 11575 21341
rect 11517 21332 11529 21335
rect 11204 21304 11529 21332
rect 11204 21292 11210 21304
rect 11517 21301 11529 21304
rect 11563 21301 11575 21335
rect 11517 21295 11575 21301
rect 13909 21335 13967 21341
rect 13909 21301 13921 21335
rect 13955 21332 13967 21335
rect 14274 21332 14280 21344
rect 13955 21304 14280 21332
rect 13955 21301 13967 21304
rect 13909 21295 13967 21301
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 17310 21292 17316 21344
rect 17368 21292 17374 21344
rect 18230 21292 18236 21344
rect 18288 21292 18294 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19720 21332 19748 21499
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24670 21496 24676 21548
rect 24728 21536 24734 21548
rect 24728 21508 25360 21536
rect 24728 21496 24734 21508
rect 20714 21428 20720 21480
rect 20772 21428 20778 21480
rect 22830 21428 22836 21480
rect 22888 21468 22894 21480
rect 23658 21468 23664 21480
rect 22888 21440 23664 21468
rect 22888 21428 22894 21440
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 24486 21428 24492 21480
rect 24544 21468 24550 21480
rect 24765 21471 24823 21477
rect 24765 21468 24777 21471
rect 24544 21440 24777 21468
rect 24544 21428 24550 21440
rect 24765 21437 24777 21440
rect 24811 21468 24823 21471
rect 25222 21468 25228 21480
rect 24811 21440 25228 21468
rect 24811 21437 24823 21440
rect 24765 21431 24823 21437
rect 25222 21428 25228 21440
rect 25280 21428 25286 21480
rect 25332 21468 25360 21508
rect 25406 21496 25412 21548
rect 25464 21536 25470 21548
rect 25501 21539 25559 21545
rect 25501 21536 25513 21539
rect 25464 21508 25513 21536
rect 25464 21496 25470 21508
rect 25501 21505 25513 21508
rect 25547 21505 25559 21539
rect 25501 21499 25559 21505
rect 25590 21496 25596 21548
rect 25648 21496 25654 21548
rect 25682 21496 25688 21548
rect 25740 21536 25746 21548
rect 25777 21539 25835 21545
rect 25777 21536 25789 21539
rect 25740 21508 25789 21536
rect 25740 21496 25746 21508
rect 25777 21505 25789 21508
rect 25823 21505 25835 21539
rect 26344 21536 26372 21632
rect 27516 21607 27574 21613
rect 27516 21573 27528 21607
rect 27562 21604 27574 21607
rect 27706 21604 27712 21616
rect 27562 21576 27712 21604
rect 27562 21573 27574 21576
rect 27516 21567 27574 21573
rect 27706 21564 27712 21576
rect 27764 21564 27770 21616
rect 27249 21539 27307 21545
rect 27249 21536 27261 21539
rect 25777 21499 25835 21505
rect 26252 21508 27261 21536
rect 26252 21480 26280 21508
rect 27249 21505 27261 21508
rect 27295 21505 27307 21539
rect 28000 21536 28028 21632
rect 33870 21604 33876 21616
rect 33428 21576 33876 21604
rect 28000 21508 29040 21536
rect 27249 21499 27307 21505
rect 25869 21471 25927 21477
rect 25869 21468 25881 21471
rect 25332 21440 25881 21468
rect 25869 21437 25881 21440
rect 25915 21437 25927 21471
rect 25869 21431 25927 21437
rect 26234 21428 26240 21480
rect 26292 21428 26298 21480
rect 26418 21428 26424 21480
rect 26476 21428 26482 21480
rect 29012 21468 29040 21508
rect 29178 21496 29184 21548
rect 29236 21536 29242 21548
rect 33428 21545 33456 21576
rect 33870 21564 33876 21576
rect 33928 21564 33934 21616
rect 34808 21604 34836 21635
rect 35342 21632 35348 21644
rect 35400 21632 35406 21684
rect 36262 21632 36268 21684
rect 36320 21672 36326 21684
rect 36320 21644 36952 21672
rect 36320 21632 36326 21644
rect 35434 21604 35440 21616
rect 34808 21576 35440 21604
rect 35434 21564 35440 21576
rect 35492 21564 35498 21616
rect 36722 21564 36728 21616
rect 36780 21564 36786 21616
rect 36924 21613 36952 21644
rect 36909 21607 36967 21613
rect 36909 21573 36921 21607
rect 36955 21573 36967 21607
rect 36909 21567 36967 21573
rect 29641 21539 29699 21545
rect 29641 21536 29653 21539
rect 29236 21508 29653 21536
rect 29236 21496 29242 21508
rect 29641 21505 29653 21508
rect 29687 21505 29699 21539
rect 30938 21539 30996 21545
rect 30938 21536 30950 21539
rect 29641 21499 29699 21505
rect 29748 21508 30950 21536
rect 29270 21468 29276 21480
rect 29012 21440 29276 21468
rect 29270 21428 29276 21440
rect 29328 21428 29334 21480
rect 29362 21428 29368 21480
rect 29420 21468 29426 21480
rect 29748 21468 29776 21508
rect 30938 21505 30950 21508
rect 30984 21505 30996 21539
rect 30938 21499 30996 21505
rect 33413 21539 33471 21545
rect 33413 21505 33425 21539
rect 33459 21505 33471 21539
rect 33413 21499 33471 21505
rect 33680 21539 33738 21545
rect 33680 21505 33692 21539
rect 33726 21536 33738 21539
rect 34238 21536 34244 21548
rect 33726 21508 34244 21536
rect 33726 21505 33738 21508
rect 33680 21499 33738 21505
rect 34238 21496 34244 21508
rect 34296 21496 34302 21548
rect 36630 21496 36636 21548
rect 36688 21496 36694 21548
rect 29420 21440 29776 21468
rect 31205 21471 31263 21477
rect 29420 21428 29426 21440
rect 31205 21437 31217 21471
rect 31251 21468 31263 21471
rect 32030 21468 32036 21480
rect 31251 21440 32036 21468
rect 31251 21437 31263 21440
rect 31205 21431 31263 21437
rect 32030 21428 32036 21440
rect 32088 21468 32094 21480
rect 33042 21468 33048 21480
rect 32088 21440 33048 21468
rect 32088 21428 32094 21440
rect 33042 21428 33048 21440
rect 33100 21428 33106 21480
rect 35529 21471 35587 21477
rect 35529 21468 35541 21471
rect 35360 21440 35541 21468
rect 23382 21360 23388 21412
rect 23440 21400 23446 21412
rect 24210 21400 24216 21412
rect 23440 21372 24216 21400
rect 23440 21360 23446 21372
rect 24210 21360 24216 21372
rect 24268 21400 24274 21412
rect 25317 21403 25375 21409
rect 25317 21400 25329 21403
rect 24268 21372 25329 21400
rect 24268 21360 24274 21372
rect 25317 21369 25329 21372
rect 25363 21369 25375 21403
rect 25317 21363 25375 21369
rect 25590 21360 25596 21412
rect 25648 21400 25654 21412
rect 26602 21400 26608 21412
rect 25648 21372 26608 21400
rect 25648 21360 25654 21372
rect 26602 21360 26608 21372
rect 26660 21360 26666 21412
rect 35360 21344 35388 21440
rect 35529 21437 35541 21440
rect 35575 21437 35587 21471
rect 35529 21431 35587 21437
rect 35713 21471 35771 21477
rect 35713 21437 35725 21471
rect 35759 21437 35771 21471
rect 35713 21431 35771 21437
rect 35728 21344 35756 21431
rect 36906 21360 36912 21412
rect 36964 21360 36970 21412
rect 19392 21304 19748 21332
rect 19392 21292 19398 21304
rect 20070 21292 20076 21344
rect 20128 21292 20134 21344
rect 20990 21292 20996 21344
rect 21048 21292 21054 21344
rect 23293 21335 23351 21341
rect 23293 21301 23305 21335
rect 23339 21332 23351 21335
rect 23474 21332 23480 21344
rect 23339 21304 23480 21332
rect 23339 21301 23351 21304
rect 23293 21295 23351 21301
rect 23474 21292 23480 21304
rect 23532 21292 23538 21344
rect 25774 21292 25780 21344
rect 25832 21292 25838 21344
rect 28718 21292 28724 21344
rect 28776 21292 28782 21344
rect 29825 21335 29883 21341
rect 29825 21301 29837 21335
rect 29871 21332 29883 21335
rect 30190 21332 30196 21344
rect 29871 21304 30196 21332
rect 29871 21301 29883 21304
rect 29825 21295 29883 21301
rect 30190 21292 30196 21304
rect 30248 21292 30254 21344
rect 35342 21292 35348 21344
rect 35400 21292 35406 21344
rect 35710 21292 35716 21344
rect 35768 21292 35774 21344
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 17681 21131 17739 21137
rect 17681 21097 17693 21131
rect 17727 21128 17739 21131
rect 17954 21128 17960 21140
rect 17727 21100 17960 21128
rect 17727 21097 17739 21100
rect 17681 21091 17739 21097
rect 17954 21088 17960 21100
rect 18012 21088 18018 21140
rect 20990 21088 20996 21140
rect 21048 21128 21054 21140
rect 21048 21100 23888 21128
rect 21048 21088 21054 21100
rect 10888 21032 12020 21060
rect 8941 20995 8999 21001
rect 8941 20961 8953 20995
rect 8987 20992 8999 20995
rect 10318 20992 10324 21004
rect 8987 20964 10324 20992
rect 8987 20961 8999 20964
rect 8941 20955 8999 20961
rect 10318 20952 10324 20964
rect 10376 20992 10382 21004
rect 10594 20992 10600 21004
rect 10376 20964 10600 20992
rect 10376 20952 10382 20964
rect 10594 20952 10600 20964
rect 10652 20992 10658 21004
rect 10888 20992 10916 21032
rect 10652 20964 10916 20992
rect 10652 20952 10658 20964
rect 10962 20952 10968 21004
rect 11020 20952 11026 21004
rect 8757 20927 8815 20933
rect 8757 20893 8769 20927
rect 8803 20893 8815 20927
rect 8757 20887 8815 20893
rect 8772 20856 8800 20887
rect 9582 20884 9588 20936
rect 9640 20884 9646 20936
rect 11054 20884 11060 20936
rect 11112 20884 11118 20936
rect 11330 20884 11336 20936
rect 11388 20884 11394 20936
rect 11517 20927 11575 20933
rect 11517 20893 11529 20927
rect 11563 20924 11575 20927
rect 11882 20924 11888 20936
rect 11563 20896 11888 20924
rect 11563 20893 11575 20896
rect 11517 20887 11575 20893
rect 11882 20884 11888 20896
rect 11940 20884 11946 20936
rect 11992 20924 12020 21032
rect 14090 20952 14096 21004
rect 14148 20952 14154 21004
rect 14274 20952 14280 21004
rect 14332 20992 14338 21004
rect 14461 20995 14519 21001
rect 14461 20992 14473 20995
rect 14332 20964 14473 20992
rect 14332 20952 14338 20964
rect 14461 20961 14473 20964
rect 14507 20961 14519 20995
rect 14461 20955 14519 20961
rect 19076 20964 19564 20992
rect 12355 20937 12413 20943
rect 12066 20924 12072 20936
rect 11992 20896 12072 20924
rect 12066 20884 12072 20896
rect 12124 20884 12130 20936
rect 12250 20884 12256 20936
rect 12308 20884 12314 20936
rect 12355 20903 12367 20937
rect 12401 20934 12413 20937
rect 12401 20924 12480 20934
rect 13262 20924 13268 20936
rect 12401 20906 13268 20924
rect 12401 20903 12413 20906
rect 12355 20897 12413 20903
rect 12452 20896 13268 20906
rect 8846 20856 8852 20868
rect 8772 20828 8852 20856
rect 8846 20816 8852 20828
rect 8904 20856 8910 20868
rect 9398 20856 9404 20868
rect 8904 20828 9404 20856
rect 8904 20816 8910 20828
rect 9398 20816 9404 20828
rect 9456 20816 9462 20868
rect 10689 20859 10747 20865
rect 10689 20825 10701 20859
rect 10735 20825 10747 20859
rect 10689 20819 10747 20825
rect 8662 20748 8668 20800
rect 8720 20748 8726 20800
rect 10704 20788 10732 20819
rect 10778 20816 10784 20868
rect 10836 20856 10842 20868
rect 11195 20859 11253 20865
rect 11195 20856 11207 20859
rect 10836 20828 11207 20856
rect 10836 20816 10842 20828
rect 11195 20825 11207 20828
rect 11241 20825 11253 20859
rect 11195 20819 11253 20825
rect 11422 20816 11428 20868
rect 11480 20816 11486 20868
rect 11701 20791 11759 20797
rect 11701 20788 11713 20791
rect 10704 20760 11713 20788
rect 11701 20757 11713 20760
rect 11747 20757 11759 20791
rect 11701 20751 11759 20757
rect 11790 20748 11796 20800
rect 11848 20788 11854 20800
rect 12452 20788 12480 20896
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 13354 20884 13360 20936
rect 13412 20884 13418 20936
rect 17310 20884 17316 20936
rect 17368 20933 17374 20936
rect 19076 20933 19104 20964
rect 17368 20924 17380 20933
rect 17589 20927 17647 20933
rect 17368 20896 17413 20924
rect 17368 20887 17380 20896
rect 17589 20893 17601 20927
rect 17635 20924 17647 20927
rect 19061 20927 19119 20933
rect 19061 20924 19073 20927
rect 17635 20896 19073 20924
rect 17635 20893 17647 20896
rect 17589 20887 17647 20893
rect 19061 20893 19073 20896
rect 19107 20893 19119 20927
rect 19061 20887 19119 20893
rect 17368 20884 17374 20887
rect 12526 20816 12532 20868
rect 12584 20816 12590 20868
rect 14826 20816 14832 20868
rect 14884 20816 14890 20868
rect 17604 20856 17632 20887
rect 19150 20884 19156 20936
rect 19208 20924 19214 20936
rect 19536 20933 19564 20964
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 19208 20896 19257 20924
rect 19208 20884 19214 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20924 19579 20927
rect 20254 20924 20260 20936
rect 19567 20896 20260 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 20254 20884 20260 20896
rect 20312 20924 20318 20936
rect 20993 20927 21051 20933
rect 20993 20924 21005 20927
rect 20312 20896 21005 20924
rect 20312 20884 20318 20896
rect 20993 20893 21005 20896
rect 21039 20924 21051 20927
rect 21542 20924 21548 20936
rect 21039 20896 21548 20924
rect 21039 20893 21051 20896
rect 20993 20887 21051 20893
rect 21542 20884 21548 20896
rect 21600 20884 21606 20936
rect 22833 20927 22891 20933
rect 22833 20893 22845 20927
rect 22879 20924 22891 20927
rect 22922 20924 22928 20936
rect 22879 20896 22928 20924
rect 22879 20893 22891 20896
rect 22833 20887 22891 20893
rect 22922 20884 22928 20896
rect 22980 20884 22986 20936
rect 17420 20828 17632 20856
rect 17420 20800 17448 20828
rect 18230 20816 18236 20868
rect 18288 20856 18294 20868
rect 18794 20859 18852 20865
rect 18794 20856 18806 20859
rect 18288 20828 18806 20856
rect 18288 20816 18294 20828
rect 18794 20825 18806 20828
rect 18840 20825 18852 20859
rect 18794 20819 18852 20825
rect 19788 20859 19846 20865
rect 19788 20825 19800 20859
rect 19834 20856 19846 20859
rect 20070 20856 20076 20868
rect 19834 20828 20076 20856
rect 19834 20825 19846 20828
rect 19788 20819 19846 20825
rect 20070 20816 20076 20828
rect 20128 20816 20134 20868
rect 21260 20859 21318 20865
rect 21260 20825 21272 20859
rect 21306 20856 21318 20859
rect 22462 20856 22468 20868
rect 21306 20828 22468 20856
rect 21306 20825 21318 20828
rect 21260 20819 21318 20825
rect 22462 20816 22468 20828
rect 22520 20816 22526 20868
rect 23106 20865 23112 20868
rect 23100 20819 23112 20865
rect 23106 20816 23112 20819
rect 23164 20816 23170 20868
rect 23860 20856 23888 21100
rect 24210 21088 24216 21140
rect 24268 21128 24274 21140
rect 25406 21128 25412 21140
rect 24268 21100 25412 21128
rect 24268 21088 24274 21100
rect 25406 21088 25412 21100
rect 25464 21088 25470 21140
rect 27798 21088 27804 21140
rect 27856 21088 27862 21140
rect 28169 21131 28227 21137
rect 28169 21097 28181 21131
rect 28215 21128 28227 21131
rect 28718 21128 28724 21140
rect 28215 21100 28724 21128
rect 28215 21097 28227 21100
rect 28169 21091 28227 21097
rect 28718 21088 28724 21100
rect 28776 21088 28782 21140
rect 29270 21088 29276 21140
rect 29328 21088 29334 21140
rect 29362 21088 29368 21140
rect 29420 21088 29426 21140
rect 29546 21088 29552 21140
rect 29604 21088 29610 21140
rect 30190 21088 30196 21140
rect 30248 21128 30254 21140
rect 30248 21100 30512 21128
rect 30248 21088 30254 21100
rect 23934 20952 23940 21004
rect 23992 20952 23998 21004
rect 27816 20992 27844 21088
rect 28353 21063 28411 21069
rect 28353 21029 28365 21063
rect 28399 21060 28411 21063
rect 29178 21060 29184 21072
rect 28399 21032 29184 21060
rect 28399 21029 28411 21032
rect 28353 21023 28411 21029
rect 29178 21020 29184 21032
rect 29236 21020 29242 21072
rect 27816 20964 28580 20992
rect 23952 20924 23980 20952
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 23952 20896 24593 20924
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24670 20884 24676 20936
rect 24728 20884 24734 20936
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 26062 20927 26120 20933
rect 26062 20924 26074 20927
rect 25832 20896 26074 20924
rect 25832 20884 25838 20896
rect 26062 20893 26074 20896
rect 26108 20893 26120 20927
rect 26062 20887 26120 20893
rect 26234 20884 26240 20936
rect 26292 20924 26298 20936
rect 26694 20933 26700 20936
rect 26329 20927 26387 20933
rect 26329 20924 26341 20927
rect 26292 20896 26341 20924
rect 26292 20884 26298 20896
rect 26329 20893 26341 20896
rect 26375 20924 26387 20927
rect 26421 20927 26479 20933
rect 26421 20924 26433 20927
rect 26375 20896 26433 20924
rect 26375 20893 26387 20896
rect 26329 20887 26387 20893
rect 26421 20893 26433 20896
rect 26467 20893 26479 20927
rect 26688 20924 26700 20933
rect 26655 20896 26700 20924
rect 26421 20887 26479 20893
rect 26688 20887 26700 20896
rect 26694 20884 26700 20887
rect 26752 20884 26758 20936
rect 28261 20927 28319 20933
rect 28261 20893 28273 20927
rect 28307 20893 28319 20927
rect 28261 20887 28319 20893
rect 28276 20856 28304 20887
rect 28442 20856 28448 20868
rect 23860 20828 28448 20856
rect 28442 20816 28448 20828
rect 28500 20816 28506 20868
rect 28552 20856 28580 20964
rect 28644 20964 28856 20992
rect 28644 20933 28672 20964
rect 28828 20936 28856 20964
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 28721 20927 28779 20933
rect 28721 20893 28733 20927
rect 28767 20893 28779 20927
rect 28721 20887 28779 20893
rect 28736 20856 28764 20887
rect 28810 20884 28816 20936
rect 28868 20884 28874 20936
rect 29181 20927 29239 20933
rect 29181 20893 29193 20927
rect 29227 20893 29239 20927
rect 29288 20924 29316 21088
rect 29564 20992 29592 21088
rect 29564 20964 30328 20992
rect 29641 20927 29699 20933
rect 29641 20924 29653 20927
rect 29288 20896 29653 20924
rect 29181 20887 29239 20893
rect 29641 20893 29653 20896
rect 29687 20893 29699 20927
rect 29641 20887 29699 20893
rect 30147 20893 30205 20899
rect 28552 20828 28764 20856
rect 29196 20856 29224 20887
rect 30147 20859 30159 20893
rect 30193 20890 30205 20893
rect 30193 20859 30220 20890
rect 30147 20856 30220 20859
rect 29196 20828 30052 20856
rect 15930 20797 15936 20800
rect 11848 20760 12480 20788
rect 15887 20791 15936 20797
rect 11848 20748 11854 20760
rect 15887 20757 15899 20791
rect 15933 20757 15936 20791
rect 15887 20751 15936 20757
rect 15930 20748 15936 20751
rect 15988 20748 15994 20800
rect 16209 20791 16267 20797
rect 16209 20757 16221 20791
rect 16255 20788 16267 20791
rect 17310 20788 17316 20800
rect 16255 20760 17316 20788
rect 16255 20757 16267 20760
rect 16209 20751 16267 20757
rect 17310 20748 17316 20760
rect 17368 20748 17374 20800
rect 17402 20748 17408 20800
rect 17460 20748 17466 20800
rect 19334 20748 19340 20800
rect 19392 20748 19398 20800
rect 20898 20748 20904 20800
rect 20956 20748 20962 20800
rect 22370 20748 22376 20800
rect 22428 20748 22434 20800
rect 24394 20748 24400 20800
rect 24452 20748 24458 20800
rect 24949 20791 25007 20797
rect 24949 20757 24961 20791
rect 24995 20788 25007 20791
rect 25222 20788 25228 20800
rect 24995 20760 25228 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 25222 20748 25228 20760
rect 25280 20748 25286 20800
rect 27890 20748 27896 20800
rect 27948 20748 27954 20800
rect 28537 20791 28595 20797
rect 28537 20757 28549 20791
rect 28583 20788 28595 20791
rect 28813 20791 28871 20797
rect 28813 20788 28825 20791
rect 28583 20760 28825 20788
rect 28583 20757 28595 20760
rect 28537 20751 28595 20757
rect 28813 20757 28825 20760
rect 28859 20757 28871 20791
rect 28813 20751 28871 20757
rect 29270 20748 29276 20800
rect 29328 20788 29334 20800
rect 30024 20797 30052 20828
rect 30116 20828 30220 20856
rect 30300 20856 30328 20964
rect 30484 20924 30512 21100
rect 34238 21088 34244 21140
rect 34296 21088 34302 21140
rect 35894 21128 35900 21140
rect 34348 21100 35900 21128
rect 32769 21063 32827 21069
rect 32769 21029 32781 21063
rect 32815 21029 32827 21063
rect 32769 21023 32827 21029
rect 32784 20992 32812 21023
rect 33134 21020 33140 21072
rect 33192 21060 33198 21072
rect 33870 21060 33876 21072
rect 33192 21032 33876 21060
rect 33192 21020 33198 21032
rect 33870 21020 33876 21032
rect 33928 21060 33934 21072
rect 34348 21060 34376 21100
rect 35894 21088 35900 21100
rect 35952 21088 35958 21140
rect 33928 21032 34376 21060
rect 33928 21020 33934 21032
rect 33413 20995 33471 21001
rect 33413 20992 33425 20995
rect 32784 20964 33425 20992
rect 33413 20961 33425 20964
rect 33459 20992 33471 20995
rect 35342 20992 35348 21004
rect 33459 20964 35348 20992
rect 33459 20961 33471 20964
rect 33413 20955 33471 20961
rect 30653 20927 30711 20933
rect 30653 20924 30665 20927
rect 30484 20896 30665 20924
rect 30377 20859 30435 20865
rect 30377 20856 30389 20859
rect 30300 20828 30389 20856
rect 30116 20800 30144 20828
rect 30377 20825 30389 20828
rect 30423 20825 30435 20859
rect 30377 20819 30435 20825
rect 30484 20800 30512 20896
rect 30653 20893 30665 20896
rect 30699 20893 30711 20927
rect 30653 20887 30711 20893
rect 31389 20927 31447 20933
rect 31389 20893 31401 20927
rect 31435 20924 31447 20927
rect 32030 20924 32036 20936
rect 31435 20896 32036 20924
rect 31435 20893 31447 20896
rect 31389 20887 31447 20893
rect 32030 20884 32036 20896
rect 32088 20884 32094 20936
rect 33870 20884 33876 20936
rect 33928 20884 33934 20936
rect 35268 20933 35296 20964
rect 35342 20952 35348 20964
rect 35400 20952 35406 21004
rect 35434 20952 35440 21004
rect 35492 20992 35498 21004
rect 35529 20995 35587 21001
rect 35529 20992 35541 20995
rect 35492 20964 35541 20992
rect 35492 20952 35498 20964
rect 35529 20961 35541 20964
rect 35575 20961 35587 20995
rect 35529 20955 35587 20961
rect 33965 20927 34023 20933
rect 33965 20893 33977 20927
rect 34011 20893 34023 20927
rect 33965 20887 34023 20893
rect 34149 20927 34207 20933
rect 34149 20893 34161 20927
rect 34195 20924 34207 20927
rect 34425 20927 34483 20933
rect 34425 20924 34437 20927
rect 34195 20896 34437 20924
rect 34195 20893 34207 20896
rect 34149 20887 34207 20893
rect 34425 20893 34437 20896
rect 34471 20893 34483 20927
rect 34425 20887 34483 20893
rect 35069 20927 35127 20933
rect 35069 20893 35081 20927
rect 35115 20893 35127 20927
rect 35069 20887 35127 20893
rect 35253 20927 35311 20933
rect 35253 20893 35265 20927
rect 35299 20924 35311 20927
rect 35299 20896 35572 20924
rect 35299 20893 35311 20896
rect 35253 20887 35311 20893
rect 31656 20859 31714 20865
rect 31656 20825 31668 20859
rect 31702 20856 31714 20859
rect 32122 20856 32128 20868
rect 31702 20828 32128 20856
rect 31702 20825 31714 20828
rect 31656 20819 31714 20825
rect 32122 20816 32128 20828
rect 32180 20816 32186 20868
rect 33980 20856 34008 20887
rect 34885 20859 34943 20865
rect 34885 20856 34897 20859
rect 33980 20828 34897 20856
rect 34885 20825 34897 20828
rect 34931 20825 34943 20859
rect 34885 20819 34943 20825
rect 35084 20800 35112 20887
rect 35544 20868 35572 20896
rect 37182 20884 37188 20936
rect 37240 20884 37246 20936
rect 38565 20927 38623 20933
rect 38565 20893 38577 20927
rect 38611 20924 38623 20927
rect 38654 20924 38660 20936
rect 38611 20896 38660 20924
rect 38611 20893 38623 20896
rect 38565 20887 38623 20893
rect 35161 20859 35219 20865
rect 35161 20825 35173 20859
rect 35207 20825 35219 20859
rect 35161 20819 35219 20825
rect 29733 20791 29791 20797
rect 29733 20788 29745 20791
rect 29328 20760 29745 20788
rect 29328 20748 29334 20760
rect 29733 20757 29745 20760
rect 29779 20757 29791 20791
rect 29733 20751 29791 20757
rect 30009 20791 30067 20797
rect 30009 20757 30021 20791
rect 30055 20757 30067 20791
rect 30009 20751 30067 20757
rect 30098 20748 30104 20800
rect 30156 20748 30162 20800
rect 30466 20748 30472 20800
rect 30524 20748 30530 20800
rect 30558 20748 30564 20800
rect 30616 20748 30622 20800
rect 32858 20748 32864 20800
rect 32916 20748 32922 20800
rect 35066 20748 35072 20800
rect 35124 20748 35130 20800
rect 35176 20788 35204 20819
rect 35342 20816 35348 20868
rect 35400 20865 35406 20868
rect 35400 20859 35429 20865
rect 35417 20825 35429 20859
rect 35400 20819 35429 20825
rect 35400 20816 35406 20819
rect 35526 20816 35532 20868
rect 35584 20816 35590 20868
rect 35710 20856 35716 20868
rect 35636 20828 35716 20856
rect 35636 20788 35664 20828
rect 35710 20816 35716 20828
rect 35768 20856 35774 20868
rect 38580 20856 38608 20887
rect 38654 20884 38660 20896
rect 38712 20884 38718 20936
rect 35768 20828 38608 20856
rect 35768 20816 35774 20828
rect 35176 20760 35664 20788
rect 37826 20748 37832 20800
rect 37884 20748 37890 20800
rect 37918 20748 37924 20800
rect 37976 20748 37982 20800
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11054 20584 11060 20596
rect 11011 20556 11060 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 11333 20587 11391 20593
rect 11333 20553 11345 20587
rect 11379 20584 11391 20587
rect 11422 20584 11428 20596
rect 11379 20556 11428 20584
rect 11379 20553 11391 20556
rect 11333 20547 11391 20553
rect 11422 20544 11428 20556
rect 11480 20544 11486 20596
rect 11698 20544 11704 20596
rect 11756 20544 11762 20596
rect 12066 20544 12072 20596
rect 12124 20584 12130 20596
rect 12345 20587 12403 20593
rect 12345 20584 12357 20587
rect 12124 20556 12357 20584
rect 12124 20544 12130 20556
rect 12345 20553 12357 20556
rect 12391 20553 12403 20587
rect 12345 20547 12403 20553
rect 14737 20587 14795 20593
rect 14737 20553 14749 20587
rect 14783 20584 14795 20587
rect 14826 20584 14832 20596
rect 14783 20556 14832 20584
rect 14783 20553 14795 20556
rect 14737 20547 14795 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 14918 20544 14924 20596
rect 14976 20584 14982 20596
rect 14976 20556 16804 20584
rect 14976 20544 14982 20556
rect 8205 20519 8263 20525
rect 8205 20485 8217 20519
rect 8251 20516 8263 20519
rect 8478 20516 8484 20528
rect 8251 20488 8484 20516
rect 8251 20485 8263 20488
rect 8205 20479 8263 20485
rect 8478 20476 8484 20488
rect 8536 20476 8542 20528
rect 8662 20476 8668 20528
rect 8720 20476 8726 20528
rect 9953 20519 10011 20525
rect 9953 20485 9965 20519
rect 9999 20516 10011 20519
rect 9999 20488 11100 20516
rect 9999 20485 10011 20488
rect 9953 20479 10011 20485
rect 11072 20460 11100 20488
rect 11238 20476 11244 20528
rect 11296 20516 11302 20528
rect 11296 20488 11836 20516
rect 11296 20476 11302 20488
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 10413 20451 10471 20457
rect 10413 20448 10425 20451
rect 10376 20420 10425 20448
rect 10376 20408 10382 20420
rect 10413 20417 10425 20420
rect 10459 20417 10471 20451
rect 10413 20411 10471 20417
rect 7926 20340 7932 20392
rect 7984 20340 7990 20392
rect 10428 20380 10456 20411
rect 11054 20408 11060 20460
rect 11112 20408 11118 20460
rect 11333 20451 11391 20457
rect 11333 20448 11345 20451
rect 11164 20420 11345 20448
rect 11164 20380 11192 20420
rect 11333 20417 11345 20420
rect 11379 20417 11391 20451
rect 11333 20411 11391 20417
rect 11609 20451 11667 20457
rect 11609 20417 11621 20451
rect 11655 20448 11667 20451
rect 11698 20448 11704 20460
rect 11655 20420 11704 20448
rect 11655 20417 11667 20420
rect 11609 20411 11667 20417
rect 10428 20352 11192 20380
rect 11054 20272 11060 20324
rect 11112 20312 11118 20324
rect 11624 20312 11652 20411
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 11808 20457 11836 20488
rect 12618 20476 12624 20528
rect 12676 20516 12682 20528
rect 12676 20488 13492 20516
rect 12676 20476 12682 20488
rect 11793 20451 11851 20457
rect 11793 20417 11805 20451
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 12437 20451 12495 20457
rect 12437 20417 12449 20451
rect 12483 20448 12495 20451
rect 12989 20451 13047 20457
rect 12483 20420 12572 20448
rect 12483 20417 12495 20420
rect 12437 20411 12495 20417
rect 11112 20284 11652 20312
rect 11112 20272 11118 20284
rect 11808 20244 11836 20411
rect 11882 20340 11888 20392
rect 11940 20380 11946 20392
rect 12544 20389 12572 20420
rect 12989 20417 13001 20451
rect 13035 20448 13047 20451
rect 13262 20448 13268 20460
rect 13035 20420 13268 20448
rect 13035 20417 13047 20420
rect 12989 20411 13047 20417
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13464 20457 13492 20488
rect 14016 20488 15240 20516
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 13906 20408 13912 20460
rect 13964 20408 13970 20460
rect 14016 20457 14044 20488
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20417 14059 20451
rect 14001 20411 14059 20417
rect 14645 20451 14703 20457
rect 14645 20417 14657 20451
rect 14691 20417 14703 20451
rect 14645 20411 14703 20417
rect 11977 20383 12035 20389
rect 11977 20380 11989 20383
rect 11940 20352 11989 20380
rect 11940 20340 11946 20352
rect 11977 20349 11989 20352
rect 12023 20349 12035 20383
rect 11977 20343 12035 20349
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 13633 20383 13691 20389
rect 13633 20380 13645 20383
rect 12529 20343 12587 20349
rect 13004 20352 13645 20380
rect 12161 20315 12219 20321
rect 12161 20281 12173 20315
rect 12207 20312 12219 20315
rect 13004 20312 13032 20352
rect 13633 20349 13645 20352
rect 13679 20349 13691 20383
rect 13633 20343 13691 20349
rect 13725 20383 13783 20389
rect 13725 20349 13737 20383
rect 13771 20380 13783 20383
rect 14016 20380 14044 20411
rect 13771 20352 14044 20380
rect 13771 20349 13783 20352
rect 13725 20343 13783 20349
rect 12207 20284 13032 20312
rect 12207 20281 12219 20284
rect 12161 20275 12219 20281
rect 14660 20256 14688 20411
rect 15212 20312 15240 20488
rect 15396 20457 15424 20556
rect 16301 20519 16359 20525
rect 16301 20516 16313 20519
rect 15672 20488 16313 20516
rect 15672 20457 15700 20488
rect 16301 20485 16313 20488
rect 16347 20485 16359 20519
rect 16301 20479 16359 20485
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20417 15439 20451
rect 15381 20411 15439 20417
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 15930 20408 15936 20460
rect 15988 20408 15994 20460
rect 16022 20408 16028 20460
rect 16080 20448 16086 20460
rect 16209 20451 16267 20457
rect 16209 20448 16221 20451
rect 16080 20420 16221 20448
rect 16080 20408 16086 20420
rect 16209 20417 16221 20420
rect 16255 20417 16267 20451
rect 16209 20411 16267 20417
rect 16393 20451 16451 20457
rect 16393 20417 16405 20451
rect 16439 20448 16451 20451
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 16439 20420 16681 20448
rect 16439 20417 16451 20420
rect 16393 20411 16451 20417
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16776 20448 16804 20556
rect 17586 20544 17592 20596
rect 17644 20544 17650 20596
rect 18046 20544 18052 20596
rect 18104 20584 18110 20596
rect 18233 20587 18291 20593
rect 18233 20584 18245 20587
rect 18104 20556 18245 20584
rect 18104 20544 18110 20556
rect 18233 20553 18245 20556
rect 18279 20553 18291 20587
rect 18233 20547 18291 20553
rect 19981 20587 20039 20593
rect 19981 20553 19993 20587
rect 20027 20584 20039 20587
rect 20714 20584 20720 20596
rect 20027 20556 20720 20584
rect 20027 20553 20039 20556
rect 19981 20547 20039 20553
rect 20714 20544 20720 20556
rect 20772 20544 20778 20596
rect 22370 20544 22376 20596
rect 22428 20544 22434 20596
rect 23017 20587 23075 20593
rect 23017 20553 23029 20587
rect 23063 20584 23075 20587
rect 23106 20584 23112 20596
rect 23063 20556 23112 20584
rect 23063 20553 23075 20556
rect 23017 20547 23075 20553
rect 23106 20544 23112 20556
rect 23164 20544 23170 20596
rect 24670 20544 24676 20596
rect 24728 20544 24734 20596
rect 26145 20587 26203 20593
rect 26145 20553 26157 20587
rect 26191 20584 26203 20587
rect 26418 20584 26424 20596
rect 26191 20556 26424 20584
rect 26191 20553 26203 20556
rect 26145 20547 26203 20553
rect 26418 20544 26424 20556
rect 26476 20544 26482 20596
rect 27706 20544 27712 20596
rect 27764 20544 27770 20596
rect 29178 20544 29184 20596
rect 29236 20584 29242 20596
rect 30009 20587 30067 20593
rect 30009 20584 30021 20587
rect 29236 20556 30021 20584
rect 29236 20544 29242 20556
rect 30009 20553 30021 20556
rect 30055 20584 30067 20587
rect 30055 20556 31524 20584
rect 30055 20553 30067 20556
rect 30009 20547 30067 20553
rect 17310 20476 17316 20528
rect 17368 20516 17374 20528
rect 17604 20516 17632 20544
rect 17773 20519 17831 20525
rect 17773 20516 17785 20519
rect 17368 20488 17785 20516
rect 17368 20476 17374 20488
rect 17773 20485 17785 20488
rect 17819 20485 17831 20519
rect 17773 20479 17831 20485
rect 17589 20451 17647 20457
rect 17589 20448 17601 20451
rect 16776 20420 17601 20448
rect 16669 20411 16727 20417
rect 17589 20417 17601 20420
rect 17635 20417 17647 20451
rect 17589 20411 17647 20417
rect 17865 20451 17923 20457
rect 17865 20417 17877 20451
rect 17911 20417 17923 20451
rect 17865 20411 17923 20417
rect 15286 20340 15292 20392
rect 15344 20380 15350 20392
rect 15948 20380 15976 20408
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 15344 20352 17233 20380
rect 15344 20340 15350 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 17221 20343 17279 20349
rect 15212 20284 15884 20312
rect 12250 20244 12256 20256
rect 11808 20216 12256 20244
rect 12250 20204 12256 20216
rect 12308 20244 12314 20256
rect 12713 20247 12771 20253
rect 12713 20244 12725 20247
rect 12308 20216 12725 20244
rect 12308 20204 12314 20216
rect 12713 20213 12725 20216
rect 12759 20213 12771 20247
rect 12713 20207 12771 20213
rect 13262 20204 13268 20256
rect 13320 20204 13326 20256
rect 14090 20204 14096 20256
rect 14148 20204 14154 20256
rect 14642 20204 14648 20256
rect 14700 20204 14706 20256
rect 15194 20204 15200 20256
rect 15252 20204 15258 20256
rect 15565 20247 15623 20253
rect 15565 20213 15577 20247
rect 15611 20244 15623 20247
rect 15749 20247 15807 20253
rect 15749 20244 15761 20247
rect 15611 20216 15761 20244
rect 15611 20213 15623 20216
rect 15565 20207 15623 20213
rect 15749 20213 15761 20216
rect 15795 20213 15807 20247
rect 15856 20244 15884 20284
rect 17880 20244 17908 20411
rect 17954 20408 17960 20460
rect 18012 20408 18018 20460
rect 18417 20451 18475 20457
rect 18417 20448 18429 20451
rect 18156 20420 18429 20448
rect 18156 20321 18184 20420
rect 18417 20417 18429 20420
rect 18463 20417 18475 20451
rect 18417 20411 18475 20417
rect 18598 20408 18604 20460
rect 18656 20408 18662 20460
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 20254 20448 20260 20460
rect 19392 20420 20260 20448
rect 19392 20408 19398 20420
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20448 20867 20451
rect 20898 20448 20904 20460
rect 20855 20420 20904 20448
rect 20855 20417 20867 20420
rect 20809 20411 20867 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20448 22339 20451
rect 22388 20448 22416 20544
rect 22922 20476 22928 20528
rect 22980 20516 22986 20528
rect 26234 20516 26240 20528
rect 22980 20488 26240 20516
rect 22980 20476 22986 20488
rect 22327 20420 22416 20448
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 23382 20408 23388 20460
rect 23440 20408 23446 20460
rect 23474 20408 23480 20460
rect 23532 20408 23538 20460
rect 23753 20451 23811 20457
rect 23753 20417 23765 20451
rect 23799 20448 23811 20451
rect 24394 20448 24400 20460
rect 23799 20420 24400 20448
rect 23799 20417 23811 20420
rect 23753 20411 23811 20417
rect 24394 20408 24400 20420
rect 24452 20408 24458 20460
rect 24780 20457 24808 20488
rect 26234 20476 26240 20488
rect 26292 20476 26298 20528
rect 28442 20476 28448 20528
rect 28500 20476 28506 20528
rect 29288 20488 30880 20516
rect 29288 20460 29316 20488
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20417 24823 20451
rect 25021 20451 25079 20457
rect 25021 20448 25033 20451
rect 24765 20411 24823 20417
rect 24872 20420 25033 20448
rect 20165 20383 20223 20389
rect 20165 20349 20177 20383
rect 20211 20349 20223 20383
rect 20165 20343 20223 20349
rect 20625 20383 20683 20389
rect 20625 20349 20637 20383
rect 20671 20380 20683 20383
rect 21174 20380 21180 20392
rect 20671 20352 21180 20380
rect 20671 20349 20683 20352
rect 20625 20343 20683 20349
rect 18141 20315 18199 20321
rect 18141 20281 18153 20315
rect 18187 20281 18199 20315
rect 20180 20312 20208 20343
rect 21174 20340 21180 20352
rect 21232 20340 21238 20392
rect 23201 20383 23259 20389
rect 23201 20349 23213 20383
rect 23247 20349 23259 20383
rect 23201 20343 23259 20349
rect 24121 20383 24179 20389
rect 24121 20349 24133 20383
rect 24167 20380 24179 20383
rect 24210 20380 24216 20392
rect 24167 20352 24216 20380
rect 24167 20349 24179 20352
rect 24121 20343 24179 20349
rect 21358 20312 21364 20324
rect 20180 20284 21364 20312
rect 18141 20275 18199 20281
rect 21358 20272 21364 20284
rect 21416 20272 21422 20324
rect 22370 20272 22376 20324
rect 22428 20312 22434 20324
rect 23216 20312 23244 20343
rect 24210 20340 24216 20352
rect 24268 20340 24274 20392
rect 24872 20380 24900 20420
rect 25021 20417 25033 20420
rect 25067 20417 25079 20451
rect 25021 20411 25079 20417
rect 27890 20408 27896 20460
rect 27948 20448 27954 20460
rect 28261 20451 28319 20457
rect 28261 20448 28273 20451
rect 27948 20420 28273 20448
rect 27948 20408 27954 20420
rect 28261 20417 28273 20420
rect 28307 20417 28319 20451
rect 28261 20411 28319 20417
rect 28721 20451 28779 20457
rect 28721 20417 28733 20451
rect 28767 20417 28779 20451
rect 28721 20411 28779 20417
rect 24780 20352 24900 20380
rect 28736 20380 28764 20411
rect 29270 20408 29276 20460
rect 29328 20408 29334 20460
rect 29917 20451 29975 20457
rect 29917 20417 29929 20451
rect 29963 20417 29975 20451
rect 29917 20411 29975 20417
rect 28810 20380 28816 20392
rect 28736 20352 28816 20380
rect 22428 20284 23244 20312
rect 22428 20272 22434 20284
rect 18506 20244 18512 20256
rect 15856 20216 18512 20244
rect 15749 20207 15807 20213
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 22186 20204 22192 20256
rect 22244 20244 22250 20256
rect 22465 20247 22523 20253
rect 22465 20244 22477 20247
rect 22244 20216 22477 20244
rect 22244 20204 22250 20216
rect 22465 20213 22477 20216
rect 22511 20244 22523 20247
rect 22830 20244 22836 20256
rect 22511 20216 22836 20244
rect 22511 20213 22523 20216
rect 22465 20207 22523 20213
rect 22830 20204 22836 20216
rect 22888 20204 22894 20256
rect 23216 20244 23244 20284
rect 23937 20315 23995 20321
rect 23937 20281 23949 20315
rect 23983 20312 23995 20315
rect 24780 20312 24808 20352
rect 28810 20340 28816 20352
rect 28868 20340 28874 20392
rect 29932 20380 29960 20411
rect 30098 20408 30104 20460
rect 30156 20408 30162 20460
rect 30558 20408 30564 20460
rect 30616 20408 30622 20460
rect 30852 20457 30880 20488
rect 30837 20451 30895 20457
rect 30837 20417 30849 20451
rect 30883 20417 30895 20451
rect 31021 20451 31079 20457
rect 31021 20448 31033 20451
rect 30837 20411 30895 20417
rect 30944 20420 31033 20448
rect 30576 20380 30604 20408
rect 29932 20352 30604 20380
rect 23983 20284 24808 20312
rect 28629 20315 28687 20321
rect 23983 20281 23995 20284
rect 23937 20275 23995 20281
rect 28629 20281 28641 20315
rect 28675 20312 28687 20315
rect 28675 20284 29132 20312
rect 28675 20281 28687 20284
rect 28629 20275 28687 20281
rect 29104 20256 29132 20284
rect 30466 20272 30472 20324
rect 30524 20312 30530 20324
rect 30944 20312 30972 20420
rect 31021 20417 31033 20420
rect 31067 20417 31079 20451
rect 31021 20411 31079 20417
rect 31386 20408 31392 20460
rect 31444 20408 31450 20460
rect 31496 20448 31524 20556
rect 32122 20544 32128 20596
rect 32180 20544 32186 20596
rect 35161 20587 35219 20593
rect 35161 20553 35173 20587
rect 35207 20584 35219 20587
rect 35342 20584 35348 20596
rect 35207 20556 35348 20584
rect 35207 20553 35219 20556
rect 35161 20547 35219 20553
rect 35342 20544 35348 20556
rect 35400 20544 35406 20596
rect 35434 20544 35440 20596
rect 35492 20584 35498 20596
rect 35897 20587 35955 20593
rect 35897 20584 35909 20587
rect 35492 20556 35909 20584
rect 35492 20544 35498 20556
rect 35897 20553 35909 20556
rect 35943 20553 35955 20587
rect 35897 20547 35955 20553
rect 36817 20587 36875 20593
rect 36817 20553 36829 20587
rect 36863 20584 36875 20587
rect 37182 20584 37188 20596
rect 36863 20556 37188 20584
rect 36863 20553 36875 20556
rect 36817 20547 36875 20553
rect 37182 20544 37188 20556
rect 37240 20544 37246 20596
rect 38654 20544 38660 20596
rect 38712 20544 38718 20596
rect 33134 20476 33140 20528
rect 33192 20516 33198 20528
rect 35618 20516 35624 20528
rect 33192 20488 33916 20516
rect 33192 20476 33198 20488
rect 31573 20451 31631 20457
rect 31573 20448 31585 20451
rect 31496 20420 31585 20448
rect 31573 20417 31585 20420
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31665 20451 31723 20457
rect 31665 20417 31677 20451
rect 31711 20448 31723 20451
rect 32858 20448 32864 20460
rect 31711 20420 32864 20448
rect 31711 20417 31723 20420
rect 31665 20411 31723 20417
rect 32858 20408 32864 20420
rect 32916 20408 32922 20460
rect 33888 20457 33916 20488
rect 35176 20488 35624 20516
rect 33689 20451 33747 20457
rect 33689 20448 33701 20451
rect 32968 20420 33701 20448
rect 31849 20383 31907 20389
rect 31849 20349 31861 20383
rect 31895 20380 31907 20383
rect 32677 20383 32735 20389
rect 32677 20380 32689 20383
rect 31895 20352 32689 20380
rect 31895 20349 31907 20352
rect 31849 20343 31907 20349
rect 32677 20349 32689 20352
rect 32723 20349 32735 20383
rect 32677 20343 32735 20349
rect 30524 20284 30972 20312
rect 31021 20315 31079 20321
rect 30524 20272 30530 20284
rect 31021 20281 31033 20315
rect 31067 20312 31079 20315
rect 31481 20315 31539 20321
rect 31481 20312 31493 20315
rect 31067 20284 31493 20312
rect 31067 20281 31079 20284
rect 31021 20275 31079 20281
rect 31481 20281 31493 20284
rect 31527 20281 31539 20315
rect 32968 20312 32996 20420
rect 33689 20417 33701 20420
rect 33735 20417 33747 20451
rect 33689 20411 33747 20417
rect 33873 20451 33931 20457
rect 33873 20417 33885 20451
rect 33919 20448 33931 20451
rect 34514 20448 34520 20460
rect 33919 20420 34520 20448
rect 33919 20417 33931 20420
rect 33873 20411 33931 20417
rect 34514 20408 34520 20420
rect 34572 20408 34578 20460
rect 35066 20408 35072 20460
rect 35124 20457 35130 20460
rect 35124 20448 35135 20457
rect 35176 20448 35204 20488
rect 35618 20476 35624 20488
rect 35676 20516 35682 20528
rect 37544 20519 37602 20525
rect 35676 20488 35756 20516
rect 35676 20476 35682 20488
rect 35124 20420 35204 20448
rect 35253 20451 35311 20457
rect 35124 20411 35135 20420
rect 35253 20417 35265 20451
rect 35299 20448 35311 20451
rect 35342 20448 35348 20460
rect 35299 20420 35348 20448
rect 35299 20417 35311 20420
rect 35253 20411 35311 20417
rect 35124 20408 35130 20411
rect 35342 20408 35348 20420
rect 35400 20408 35406 20460
rect 35526 20408 35532 20460
rect 35584 20408 35590 20460
rect 35728 20457 35756 20488
rect 36372 20488 36860 20516
rect 35713 20451 35771 20457
rect 35713 20417 35725 20451
rect 35759 20446 35771 20451
rect 35802 20446 35808 20460
rect 35759 20418 35808 20446
rect 35759 20417 35771 20418
rect 35713 20411 35771 20417
rect 35802 20408 35808 20418
rect 35860 20448 35866 20460
rect 35860 20420 35953 20448
rect 35860 20408 35866 20420
rect 36078 20408 36084 20460
rect 36136 20408 36142 20460
rect 36170 20408 36176 20460
rect 36228 20408 36234 20460
rect 36372 20457 36400 20488
rect 36722 20457 36728 20460
rect 36321 20451 36400 20457
rect 36321 20417 36333 20451
rect 36367 20420 36400 20451
rect 36449 20451 36507 20457
rect 36367 20417 36379 20420
rect 36321 20411 36379 20417
rect 36449 20417 36461 20451
rect 36495 20417 36507 20451
rect 36449 20411 36507 20417
rect 36541 20451 36599 20457
rect 36541 20417 36553 20451
rect 36587 20417 36599 20451
rect 36541 20411 36599 20417
rect 36679 20451 36728 20457
rect 36679 20417 36691 20451
rect 36725 20417 36728 20451
rect 36679 20411 36728 20417
rect 33965 20383 34023 20389
rect 33965 20380 33977 20383
rect 31481 20275 31539 20281
rect 32784 20284 32996 20312
rect 33704 20352 33977 20380
rect 23382 20244 23388 20256
rect 23216 20216 23388 20244
rect 23382 20204 23388 20216
rect 23440 20244 23446 20256
rect 23750 20244 23756 20256
rect 23440 20216 23756 20244
rect 23440 20204 23446 20216
rect 23750 20204 23756 20216
rect 23808 20244 23814 20256
rect 24302 20244 24308 20256
rect 23808 20216 24308 20244
rect 23808 20204 23814 20216
rect 24302 20204 24308 20216
rect 24360 20204 24366 20256
rect 28534 20204 28540 20256
rect 28592 20204 28598 20256
rect 29086 20204 29092 20256
rect 29144 20204 29150 20256
rect 32674 20204 32680 20256
rect 32732 20244 32738 20256
rect 32784 20244 32812 20284
rect 33704 20256 33732 20352
rect 33965 20349 33977 20352
rect 34011 20349 34023 20383
rect 33965 20343 34023 20349
rect 35621 20383 35679 20389
rect 35621 20349 35633 20383
rect 35667 20380 35679 20383
rect 36464 20380 36492 20411
rect 35667 20352 36492 20380
rect 35667 20349 35679 20352
rect 35621 20343 35679 20349
rect 36556 20312 36584 20411
rect 36722 20408 36728 20411
rect 36780 20408 36786 20460
rect 36832 20448 36860 20488
rect 37544 20485 37556 20519
rect 37590 20516 37602 20519
rect 37826 20516 37832 20528
rect 37590 20488 37832 20516
rect 37590 20485 37602 20488
rect 37544 20479 37602 20485
rect 37826 20476 37832 20488
rect 37884 20476 37890 20528
rect 37918 20448 37924 20460
rect 36832 20420 37924 20448
rect 37918 20408 37924 20420
rect 37976 20408 37982 20460
rect 37274 20340 37280 20392
rect 37332 20340 37338 20392
rect 35912 20284 36584 20312
rect 35912 20256 35940 20284
rect 32732 20216 32812 20244
rect 32732 20204 32738 20216
rect 32858 20204 32864 20256
rect 32916 20244 32922 20256
rect 33505 20247 33563 20253
rect 33505 20244 33517 20247
rect 32916 20216 33517 20244
rect 32916 20204 32922 20216
rect 33505 20213 33517 20216
rect 33551 20213 33563 20247
rect 33505 20207 33563 20213
rect 33686 20204 33692 20256
rect 33744 20204 33750 20256
rect 35894 20204 35900 20256
rect 35952 20204 35958 20256
rect 36081 20247 36139 20253
rect 36081 20213 36093 20247
rect 36127 20244 36139 20247
rect 37182 20244 37188 20256
rect 36127 20216 37188 20244
rect 36127 20213 36139 20216
rect 36081 20207 36139 20213
rect 37182 20204 37188 20216
rect 37240 20204 37246 20256
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 9582 20000 9588 20052
rect 9640 20000 9646 20052
rect 15194 20000 15200 20052
rect 15252 20000 15258 20052
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 17037 20043 17095 20049
rect 17037 20040 17049 20043
rect 16080 20012 17049 20040
rect 16080 20000 16086 20012
rect 17037 20009 17049 20012
rect 17083 20040 17095 20043
rect 20070 20040 20076 20052
rect 17083 20012 20076 20040
rect 17083 20009 17095 20012
rect 17037 20003 17095 20009
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 21358 20000 21364 20052
rect 21416 20000 21422 20052
rect 22462 20000 22468 20052
rect 22520 20000 22526 20052
rect 22554 20000 22560 20052
rect 22612 20000 22618 20052
rect 23014 20000 23020 20052
rect 23072 20000 23078 20052
rect 23753 20043 23811 20049
rect 23753 20009 23765 20043
rect 23799 20040 23811 20043
rect 23934 20040 23940 20052
rect 23799 20012 23940 20040
rect 23799 20009 23811 20012
rect 23753 20003 23811 20009
rect 23934 20000 23940 20012
rect 23992 20000 23998 20052
rect 28534 20000 28540 20052
rect 28592 20000 28598 20052
rect 29086 20000 29092 20052
rect 29144 20000 29150 20052
rect 29362 20000 29368 20052
rect 29420 20040 29426 20052
rect 30466 20040 30472 20052
rect 29420 20012 30472 20040
rect 29420 20000 29426 20012
rect 30466 20000 30472 20012
rect 30524 20000 30530 20052
rect 32766 20000 32772 20052
rect 32824 20040 32830 20052
rect 35253 20043 35311 20049
rect 32824 20012 35204 20040
rect 32824 20000 32830 20012
rect 15212 19972 15240 20000
rect 15212 19944 15424 19972
rect 10597 19907 10655 19913
rect 10597 19873 10609 19907
rect 10643 19904 10655 19907
rect 10870 19904 10876 19916
rect 10643 19876 10876 19904
rect 10643 19873 10655 19876
rect 10597 19867 10655 19873
rect 10870 19864 10876 19876
rect 10928 19904 10934 19916
rect 12526 19904 12532 19916
rect 10928 19876 12532 19904
rect 10928 19864 10934 19876
rect 12526 19864 12532 19876
rect 12584 19904 12590 19916
rect 15289 19907 15347 19913
rect 15289 19904 15301 19907
rect 12584 19876 15301 19904
rect 12584 19864 12590 19876
rect 15289 19873 15301 19876
rect 15335 19873 15347 19907
rect 15396 19904 15424 19944
rect 15565 19907 15623 19913
rect 15565 19904 15577 19907
rect 15396 19876 15577 19904
rect 15289 19867 15347 19873
rect 15565 19873 15577 19876
rect 15611 19873 15623 19907
rect 21376 19904 21404 20000
rect 22278 19932 22284 19984
rect 22336 19932 22342 19984
rect 24026 19972 24032 19984
rect 23124 19944 24032 19972
rect 21821 19907 21879 19913
rect 21821 19904 21833 19907
rect 21376 19876 21833 19904
rect 15565 19867 15623 19873
rect 21821 19873 21833 19876
rect 21867 19873 21879 19907
rect 22296 19904 22324 19932
rect 22296 19876 22876 19904
rect 21821 19867 21879 19873
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 12250 19796 12256 19848
rect 12308 19836 12314 19848
rect 12621 19839 12679 19845
rect 12621 19836 12633 19839
rect 12308 19808 12633 19836
rect 12308 19796 12314 19808
rect 12621 19805 12633 19808
rect 12667 19805 12679 19839
rect 12621 19799 12679 19805
rect 20254 19796 20260 19848
rect 20312 19836 20318 19848
rect 20533 19839 20591 19845
rect 20533 19836 20545 19839
rect 20312 19808 20545 19836
rect 20312 19796 20318 19808
rect 20533 19805 20545 19808
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 20714 19796 20720 19848
rect 20772 19796 20778 19848
rect 21082 19836 21088 19848
rect 20824 19808 21088 19836
rect 10873 19771 10931 19777
rect 2746 19740 9720 19768
rect 1762 19660 1768 19712
rect 1820 19700 1826 19712
rect 2746 19700 2774 19740
rect 1820 19672 2774 19700
rect 9692 19700 9720 19740
rect 10873 19737 10885 19771
rect 10919 19768 10931 19771
rect 11146 19768 11152 19780
rect 10919 19740 11152 19768
rect 10919 19737 10931 19740
rect 10873 19731 10931 19737
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 11606 19728 11612 19780
rect 11664 19728 11670 19780
rect 12805 19771 12863 19777
rect 12805 19737 12817 19771
rect 12851 19737 12863 19771
rect 12805 19731 12863 19737
rect 12820 19700 12848 19731
rect 12986 19728 12992 19780
rect 13044 19728 13050 19780
rect 14090 19728 14096 19780
rect 14148 19768 14154 19780
rect 15562 19768 15568 19780
rect 14148 19740 15568 19768
rect 14148 19728 14154 19740
rect 15562 19728 15568 19740
rect 15620 19728 15626 19780
rect 16298 19728 16304 19780
rect 16356 19728 16362 19780
rect 19978 19768 19984 19780
rect 16960 19740 19984 19768
rect 9692 19672 12848 19700
rect 1820 19660 1826 19672
rect 16206 19660 16212 19712
rect 16264 19700 16270 19712
rect 16960 19700 16988 19740
rect 19978 19728 19984 19740
rect 20036 19768 20042 19780
rect 20824 19768 20852 19808
rect 21082 19796 21088 19808
rect 21140 19796 21146 19848
rect 22186 19796 22192 19848
rect 22244 19796 22250 19848
rect 22281 19839 22339 19845
rect 22281 19805 22293 19839
rect 22327 19836 22339 19839
rect 22370 19836 22376 19848
rect 22327 19808 22376 19836
rect 22327 19805 22339 19808
rect 22281 19799 22339 19805
rect 22370 19796 22376 19808
rect 22428 19796 22434 19848
rect 22462 19796 22468 19848
rect 22520 19836 22526 19848
rect 22848 19845 22876 19876
rect 23124 19845 23152 19944
rect 24026 19932 24032 19944
rect 24084 19932 24090 19984
rect 23845 19907 23903 19913
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 24673 19907 24731 19913
rect 24673 19904 24685 19907
rect 23891 19876 24685 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 24673 19873 24685 19876
rect 24719 19873 24731 19907
rect 24673 19867 24731 19873
rect 25222 19864 25228 19916
rect 25280 19864 25286 19916
rect 26234 19864 26240 19916
rect 26292 19904 26298 19916
rect 27522 19904 27528 19916
rect 26292 19876 27528 19904
rect 26292 19864 26298 19876
rect 27522 19864 27528 19876
rect 27580 19864 27586 19916
rect 22741 19839 22799 19845
rect 22741 19836 22753 19839
rect 22520 19808 22753 19836
rect 22520 19796 22526 19808
rect 22741 19805 22753 19808
rect 22787 19805 22799 19839
rect 22741 19799 22799 19805
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19805 22891 19839
rect 22833 19799 22891 19805
rect 23109 19839 23167 19845
rect 23109 19805 23121 19839
rect 23155 19805 23167 19839
rect 23109 19799 23167 19805
rect 23290 19796 23296 19848
rect 23348 19796 23354 19848
rect 23566 19796 23572 19848
rect 23624 19796 23630 19848
rect 23750 19796 23756 19848
rect 23808 19796 23814 19848
rect 23934 19796 23940 19848
rect 23992 19836 23998 19848
rect 24029 19839 24087 19845
rect 24029 19836 24041 19839
rect 23992 19808 24041 19836
rect 23992 19796 23998 19808
rect 24029 19805 24041 19808
rect 24075 19805 24087 19839
rect 24029 19799 24087 19805
rect 24213 19839 24271 19845
rect 24213 19805 24225 19839
rect 24259 19836 24271 19839
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 24259 19808 24409 19836
rect 24259 19805 24271 19808
rect 24213 19799 24271 19805
rect 24397 19805 24409 19808
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 27792 19839 27850 19845
rect 27792 19805 27804 19839
rect 27838 19836 27850 19839
rect 28552 19836 28580 20000
rect 28905 19975 28963 19981
rect 28905 19941 28917 19975
rect 28951 19972 28963 19975
rect 29730 19972 29736 19984
rect 28951 19944 29736 19972
rect 28951 19941 28963 19944
rect 28905 19935 28963 19941
rect 29730 19932 29736 19944
rect 29788 19972 29794 19984
rect 29788 19944 30144 19972
rect 29788 19932 29794 19944
rect 30116 19913 30144 19944
rect 30101 19907 30159 19913
rect 29288 19876 30052 19904
rect 29288 19848 29316 19876
rect 27838 19808 28580 19836
rect 27838 19805 27850 19808
rect 27792 19799 27850 19805
rect 29270 19796 29276 19848
rect 29328 19796 29334 19848
rect 29362 19796 29368 19848
rect 29420 19796 29426 19848
rect 30024 19836 30052 19876
rect 30101 19873 30113 19907
rect 30147 19904 30159 19907
rect 30285 19907 30343 19913
rect 30285 19904 30297 19907
rect 30147 19876 30297 19904
rect 30147 19873 30159 19876
rect 30101 19867 30159 19873
rect 30285 19873 30297 19876
rect 30331 19873 30343 19907
rect 30484 19904 30512 20000
rect 35176 19904 35204 20012
rect 35253 20009 35265 20043
rect 35299 20040 35311 20043
rect 35342 20040 35348 20052
rect 35299 20012 35348 20040
rect 35299 20009 35311 20012
rect 35253 20003 35311 20009
rect 35342 20000 35348 20012
rect 35400 20000 35406 20052
rect 35434 20000 35440 20052
rect 35492 20040 35498 20052
rect 35529 20043 35587 20049
rect 35529 20040 35541 20043
rect 35492 20012 35541 20040
rect 35492 20000 35498 20012
rect 35529 20009 35541 20012
rect 35575 20009 35587 20043
rect 35529 20003 35587 20009
rect 35897 20043 35955 20049
rect 35897 20009 35909 20043
rect 35943 20040 35955 20043
rect 36078 20040 36084 20052
rect 35943 20012 36084 20040
rect 35943 20009 35955 20012
rect 35897 20003 35955 20009
rect 36078 20000 36084 20012
rect 36136 20000 36142 20052
rect 37182 20000 37188 20052
rect 37240 20000 37246 20052
rect 35250 19904 35256 19916
rect 30484 19876 30604 19904
rect 35176 19876 35256 19904
rect 30285 19867 30343 19873
rect 30576 19845 30604 19876
rect 35250 19864 35256 19876
rect 35308 19904 35314 19916
rect 36170 19904 36176 19916
rect 35308 19876 36176 19904
rect 35308 19864 35314 19876
rect 36170 19864 36176 19876
rect 36228 19904 36234 19916
rect 36998 19904 37004 19916
rect 36228 19876 37004 19904
rect 36228 19864 36234 19876
rect 36998 19864 37004 19876
rect 37056 19864 37062 19916
rect 37200 19913 37228 20000
rect 37185 19907 37243 19913
rect 37185 19873 37197 19907
rect 37231 19873 37243 19907
rect 37185 19867 37243 19873
rect 30469 19839 30527 19845
rect 30469 19836 30481 19839
rect 30024 19808 30481 19836
rect 30469 19805 30481 19808
rect 30515 19805 30527 19839
rect 30469 19799 30527 19805
rect 30561 19839 30619 19845
rect 30561 19805 30573 19839
rect 30607 19805 30619 19839
rect 30561 19799 30619 19805
rect 32030 19796 32036 19848
rect 32088 19836 32094 19848
rect 34333 19839 34391 19845
rect 32088 19808 32996 19836
rect 32088 19796 32094 19808
rect 21959 19771 22017 19777
rect 21959 19768 21971 19771
rect 20036 19740 20852 19768
rect 20916 19740 21971 19768
rect 20036 19728 20042 19740
rect 20916 19712 20944 19740
rect 21959 19737 21971 19740
rect 22005 19737 22017 19771
rect 21959 19731 22017 19737
rect 22097 19771 22155 19777
rect 22097 19737 22109 19771
rect 22143 19768 22155 19771
rect 22646 19768 22652 19780
rect 22143 19740 22652 19768
rect 22143 19737 22155 19740
rect 22097 19731 22155 19737
rect 22646 19728 22652 19740
rect 22704 19768 22710 19780
rect 23308 19768 23336 19796
rect 32968 19780 32996 19808
rect 34333 19805 34345 19839
rect 34379 19805 34391 19839
rect 34333 19799 34391 19805
rect 35069 19839 35127 19845
rect 35069 19805 35081 19839
rect 35115 19836 35127 19839
rect 35894 19836 35900 19848
rect 35115 19808 35900 19836
rect 35115 19805 35127 19808
rect 35069 19799 35127 19805
rect 22704 19740 23336 19768
rect 29089 19771 29147 19777
rect 22704 19728 22710 19740
rect 29089 19737 29101 19771
rect 29135 19768 29147 19771
rect 29549 19771 29607 19777
rect 29549 19768 29561 19771
rect 29135 19740 29561 19768
rect 29135 19737 29147 19740
rect 29089 19731 29147 19737
rect 29549 19737 29561 19740
rect 29595 19737 29607 19771
rect 30653 19771 30711 19777
rect 30653 19768 30665 19771
rect 29549 19731 29607 19737
rect 30116 19740 30665 19768
rect 30116 19712 30144 19740
rect 30653 19737 30665 19740
rect 30699 19737 30711 19771
rect 30653 19731 30711 19737
rect 32300 19771 32358 19777
rect 32300 19737 32312 19771
rect 32346 19768 32358 19771
rect 32858 19768 32864 19780
rect 32346 19740 32864 19768
rect 32346 19737 32358 19740
rect 32300 19731 32358 19737
rect 32858 19728 32864 19740
rect 32916 19728 32922 19780
rect 32950 19728 32956 19780
rect 33008 19728 33014 19780
rect 33686 19768 33692 19780
rect 33336 19740 33692 19768
rect 16264 19672 16988 19700
rect 20625 19703 20683 19709
rect 16264 19660 16270 19672
rect 20625 19669 20637 19703
rect 20671 19700 20683 19703
rect 20898 19700 20904 19712
rect 20671 19672 20904 19700
rect 20671 19669 20683 19672
rect 20625 19663 20683 19669
rect 20898 19660 20904 19672
rect 20956 19660 20962 19712
rect 24578 19660 24584 19712
rect 24636 19660 24642 19712
rect 30098 19660 30104 19712
rect 30156 19660 30162 19712
rect 30558 19660 30564 19712
rect 30616 19700 30622 19712
rect 30837 19703 30895 19709
rect 30837 19700 30849 19703
rect 30616 19672 30849 19700
rect 30616 19660 30622 19672
rect 30837 19669 30849 19672
rect 30883 19669 30895 19703
rect 30837 19663 30895 19669
rect 32766 19660 32772 19712
rect 32824 19700 32830 19712
rect 33336 19700 33364 19740
rect 33686 19728 33692 19740
rect 33744 19728 33750 19780
rect 32824 19672 33364 19700
rect 32824 19660 32830 19672
rect 33410 19660 33416 19712
rect 33468 19700 33474 19712
rect 34348 19700 34376 19799
rect 35894 19796 35900 19808
rect 35952 19796 35958 19848
rect 36541 19839 36599 19845
rect 36541 19805 36553 19839
rect 36587 19836 36599 19839
rect 36587 19808 37044 19836
rect 36587 19805 36599 19808
rect 36541 19799 36599 19805
rect 34606 19728 34612 19780
rect 34664 19768 34670 19780
rect 34701 19771 34759 19777
rect 34701 19768 34713 19771
rect 34664 19740 34713 19768
rect 34664 19728 34670 19740
rect 34701 19737 34713 19740
rect 34747 19737 34759 19771
rect 34701 19731 34759 19737
rect 34977 19771 35035 19777
rect 34977 19737 34989 19771
rect 35023 19768 35035 19771
rect 35713 19771 35771 19777
rect 35713 19768 35725 19771
rect 35023 19740 35725 19768
rect 35023 19737 35035 19740
rect 34977 19731 35035 19737
rect 35713 19737 35725 19740
rect 35759 19768 35771 19771
rect 36556 19768 36584 19799
rect 35759 19740 36584 19768
rect 35759 19737 35771 19740
rect 35713 19731 35771 19737
rect 37016 19712 37044 19808
rect 34882 19700 34888 19712
rect 33468 19672 34888 19700
rect 33468 19660 33474 19672
rect 34882 19660 34888 19672
rect 34940 19660 34946 19712
rect 35158 19660 35164 19712
rect 35216 19700 35222 19712
rect 35526 19709 35532 19712
rect 35345 19703 35403 19709
rect 35345 19700 35357 19703
rect 35216 19672 35357 19700
rect 35216 19660 35222 19672
rect 35345 19669 35357 19672
rect 35391 19669 35403 19703
rect 35345 19663 35403 19669
rect 35513 19703 35532 19709
rect 35513 19669 35525 19703
rect 35513 19663 35532 19669
rect 35526 19660 35532 19663
rect 35584 19660 35590 19712
rect 35618 19660 35624 19712
rect 35676 19700 35682 19712
rect 36633 19703 36691 19709
rect 36633 19700 36645 19703
rect 35676 19672 36645 19700
rect 35676 19660 35682 19672
rect 36633 19669 36645 19672
rect 36679 19669 36691 19703
rect 36633 19663 36691 19669
rect 36998 19660 37004 19712
rect 37056 19660 37062 19712
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11664 19468 11713 19496
rect 11664 19456 11670 19468
rect 11701 19465 11713 19468
rect 11747 19465 11759 19499
rect 11701 19459 11759 19465
rect 12986 19456 12992 19508
rect 13044 19496 13050 19508
rect 13081 19499 13139 19505
rect 13081 19496 13093 19499
rect 13044 19468 13093 19496
rect 13044 19456 13050 19468
rect 13081 19465 13093 19468
rect 13127 19465 13139 19499
rect 16206 19496 16212 19508
rect 13081 19459 13139 19465
rect 15580 19468 16212 19496
rect 14642 19428 14648 19440
rect 11624 19400 14648 19428
rect 11624 19369 11652 19400
rect 14642 19388 14648 19400
rect 14700 19428 14706 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 14700 19400 15393 19428
rect 14700 19388 14706 19400
rect 15381 19397 15393 19400
rect 15427 19397 15439 19431
rect 15381 19391 15439 19397
rect 11609 19363 11667 19369
rect 11609 19360 11621 19363
rect 11072 19332 11621 19360
rect 11072 19304 11100 19332
rect 11609 19329 11621 19332
rect 11655 19329 11667 19363
rect 11609 19323 11667 19329
rect 13446 19320 13452 19372
rect 13504 19320 13510 19372
rect 13541 19363 13599 19369
rect 13541 19329 13553 19363
rect 13587 19360 13599 19363
rect 14274 19360 14280 19372
rect 13587 19332 14280 19360
rect 13587 19329 13599 19332
rect 13541 19323 13599 19329
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 15580 19360 15608 19468
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 16298 19456 16304 19508
rect 16356 19496 16362 19508
rect 16393 19499 16451 19505
rect 16393 19496 16405 19499
rect 16356 19468 16405 19496
rect 16356 19456 16362 19468
rect 16393 19465 16405 19468
rect 16439 19465 16451 19499
rect 16393 19459 16451 19465
rect 18506 19456 18512 19508
rect 18564 19456 18570 19508
rect 20990 19496 20996 19508
rect 19444 19468 20996 19496
rect 19444 19428 19472 19468
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21361 19499 21419 19505
rect 21361 19465 21373 19499
rect 21407 19496 21419 19499
rect 23201 19499 23259 19505
rect 23201 19496 23213 19499
rect 21407 19468 22094 19496
rect 21407 19465 21419 19468
rect 21361 19459 21419 19465
rect 21542 19428 21548 19440
rect 15672 19400 19472 19428
rect 19904 19400 21548 19428
rect 15672 19369 15700 19400
rect 14507 19332 15608 19360
rect 15657 19363 15715 19369
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 15657 19329 15669 19363
rect 15703 19329 15715 19363
rect 15657 19323 15715 19329
rect 16298 19320 16304 19372
rect 16356 19320 16362 19372
rect 17310 19369 17316 19372
rect 17304 19323 17316 19369
rect 17310 19320 17316 19323
rect 17368 19320 17374 19372
rect 19633 19363 19691 19369
rect 19633 19329 19645 19363
rect 19679 19360 19691 19363
rect 19794 19360 19800 19372
rect 19679 19332 19800 19360
rect 19679 19329 19691 19332
rect 19633 19323 19691 19329
rect 19794 19320 19800 19332
rect 19852 19320 19858 19372
rect 19904 19369 19932 19400
rect 21542 19388 21548 19400
rect 21600 19428 21606 19440
rect 22066 19437 22094 19468
rect 22296 19468 23213 19496
rect 22296 19440 22324 19468
rect 23201 19465 23213 19468
rect 23247 19465 23259 19499
rect 23201 19459 23259 19465
rect 29730 19456 29736 19508
rect 29788 19456 29794 19508
rect 30650 19456 30656 19508
rect 30708 19496 30714 19508
rect 31846 19496 31852 19508
rect 30708 19468 31852 19496
rect 30708 19456 30714 19468
rect 31846 19456 31852 19468
rect 31904 19456 31910 19508
rect 32766 19456 32772 19508
rect 32824 19456 32830 19508
rect 32950 19456 32956 19508
rect 33008 19496 33014 19508
rect 33008 19468 35664 19496
rect 33008 19456 33014 19468
rect 22066 19431 22124 19437
rect 21600 19400 21864 19428
rect 21600 19388 21606 19400
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 19978 19320 19984 19372
rect 20036 19360 20042 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 20036 19332 20269 19360
rect 20036 19320 20042 19332
rect 20257 19329 20269 19332
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 11054 19252 11060 19304
rect 11112 19252 11118 19304
rect 13725 19295 13783 19301
rect 13725 19261 13737 19295
rect 13771 19292 13783 19295
rect 14090 19292 14096 19304
rect 13771 19264 14096 19292
rect 13771 19261 13783 19264
rect 13725 19255 13783 19261
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 17037 19295 17095 19301
rect 17037 19261 17049 19295
rect 17083 19261 17095 19295
rect 17037 19255 17095 19261
rect 14369 19159 14427 19165
rect 14369 19125 14381 19159
rect 14415 19156 14427 19159
rect 14458 19156 14464 19168
rect 14415 19128 14464 19156
rect 14415 19125 14427 19128
rect 14369 19119 14427 19125
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 17052 19156 17080 19255
rect 20548 19224 20576 19323
rect 20622 19320 20628 19372
rect 20680 19360 20686 19372
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20680 19332 20821 19360
rect 20680 19320 20686 19332
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 20898 19320 20904 19372
rect 20956 19360 20962 19372
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20956 19332 21005 19360
rect 20956 19320 20962 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 21100 19292 21128 19323
rect 21174 19320 21180 19372
rect 21232 19320 21238 19372
rect 21266 19320 21272 19372
rect 21324 19360 21330 19372
rect 21453 19363 21511 19369
rect 21453 19360 21465 19363
rect 21324 19332 21465 19360
rect 21324 19320 21330 19332
rect 21453 19329 21465 19332
rect 21499 19329 21511 19363
rect 21453 19323 21511 19329
rect 21634 19320 21640 19372
rect 21692 19320 21698 19372
rect 21836 19369 21864 19400
rect 22066 19397 22078 19431
rect 22112 19397 22124 19431
rect 22066 19391 22124 19397
rect 22278 19388 22284 19440
rect 22336 19388 22342 19440
rect 22940 19400 25360 19428
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 22296 19360 22324 19388
rect 22940 19372 22968 19400
rect 21821 19323 21879 19329
rect 21928 19332 22324 19360
rect 21928 19292 21956 19332
rect 22922 19320 22928 19372
rect 22980 19320 22986 19372
rect 23290 19320 23296 19372
rect 23348 19360 23354 19372
rect 23477 19363 23535 19369
rect 23477 19360 23489 19363
rect 23348 19332 23489 19360
rect 23348 19320 23354 19332
rect 23477 19329 23489 19332
rect 23523 19329 23535 19363
rect 23477 19323 23535 19329
rect 24578 19320 24584 19372
rect 24636 19360 24642 19372
rect 25332 19369 25360 19400
rect 26510 19388 26516 19440
rect 26568 19428 26574 19440
rect 27065 19431 27123 19437
rect 27065 19428 27077 19431
rect 26568 19400 27077 19428
rect 26568 19388 26574 19400
rect 27065 19397 27077 19400
rect 27111 19397 27123 19431
rect 27065 19391 27123 19397
rect 27617 19431 27675 19437
rect 27617 19397 27629 19431
rect 27663 19428 27675 19431
rect 28074 19428 28080 19440
rect 27663 19400 28080 19428
rect 27663 19397 27675 19400
rect 27617 19391 27675 19397
rect 28074 19388 28080 19400
rect 28132 19388 28138 19440
rect 25682 19369 25688 19372
rect 25050 19363 25108 19369
rect 25050 19360 25062 19363
rect 24636 19332 25062 19360
rect 24636 19320 24642 19332
rect 25050 19329 25062 19332
rect 25096 19329 25108 19363
rect 25050 19323 25108 19329
rect 25317 19363 25375 19369
rect 25317 19329 25329 19363
rect 25363 19360 25375 19363
rect 25409 19363 25467 19369
rect 25409 19360 25421 19363
rect 25363 19332 25421 19360
rect 25363 19329 25375 19332
rect 25317 19323 25375 19329
rect 25409 19329 25421 19332
rect 25455 19329 25467 19363
rect 25409 19323 25467 19329
rect 25676 19323 25688 19369
rect 25682 19320 25688 19323
rect 25740 19320 25746 19372
rect 29748 19369 29776 19456
rect 31386 19428 31392 19440
rect 30392 19400 31392 19428
rect 29733 19363 29791 19369
rect 29733 19329 29745 19363
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29914 19320 29920 19372
rect 29972 19320 29978 19372
rect 30193 19363 30251 19369
rect 30193 19329 30205 19363
rect 30239 19360 30251 19363
rect 30282 19360 30288 19372
rect 30239 19332 30288 19360
rect 30239 19329 30251 19332
rect 30193 19323 30251 19329
rect 30282 19320 30288 19332
rect 30340 19320 30346 19372
rect 21100 19264 21956 19292
rect 30098 19252 30104 19304
rect 30156 19252 30162 19304
rect 20714 19224 20720 19236
rect 20548 19196 20720 19224
rect 20714 19184 20720 19196
rect 20772 19224 20778 19236
rect 20772 19196 20944 19224
rect 20772 19184 20778 19196
rect 20916 19168 20944 19196
rect 21174 19184 21180 19236
rect 21232 19224 21238 19236
rect 21637 19227 21695 19233
rect 21637 19224 21649 19227
rect 21232 19196 21649 19224
rect 21232 19184 21238 19196
rect 21637 19193 21649 19196
rect 21683 19193 21695 19227
rect 21637 19187 21695 19193
rect 27246 19184 27252 19236
rect 27304 19224 27310 19236
rect 30392 19224 30420 19400
rect 31386 19388 31392 19400
rect 31444 19388 31450 19440
rect 31662 19388 31668 19440
rect 31720 19437 31726 19440
rect 31720 19431 31743 19437
rect 31731 19397 31743 19431
rect 31720 19391 31743 19397
rect 31720 19388 31726 19391
rect 30469 19363 30527 19369
rect 30469 19329 30481 19363
rect 30515 19360 30527 19363
rect 30515 19332 30604 19360
rect 30515 19329 30527 19332
rect 30469 19323 30527 19329
rect 27304 19196 30420 19224
rect 27304 19184 27310 19196
rect 17402 19156 17408 19168
rect 17052 19128 17408 19156
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 18414 19116 18420 19168
rect 18472 19116 18478 19168
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 21266 19156 21272 19168
rect 20956 19128 21272 19156
rect 20956 19116 20962 19128
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 23474 19116 23480 19168
rect 23532 19156 23538 19168
rect 23569 19159 23627 19165
rect 23569 19156 23581 19159
rect 23532 19128 23581 19156
rect 23532 19116 23538 19128
rect 23569 19125 23581 19128
rect 23615 19125 23627 19159
rect 23569 19119 23627 19125
rect 23934 19116 23940 19168
rect 23992 19116 23998 19168
rect 26050 19116 26056 19168
rect 26108 19156 26114 19168
rect 26789 19159 26847 19165
rect 26789 19156 26801 19159
rect 26108 19128 26801 19156
rect 26108 19116 26114 19128
rect 26789 19125 26801 19128
rect 26835 19125 26847 19159
rect 26789 19119 26847 19125
rect 26878 19116 26884 19168
rect 26936 19156 26942 19168
rect 27157 19159 27215 19165
rect 27157 19156 27169 19159
rect 26936 19128 27169 19156
rect 26936 19116 26942 19128
rect 27157 19125 27169 19128
rect 27203 19125 27215 19159
rect 27157 19119 27215 19125
rect 27706 19116 27712 19168
rect 27764 19116 27770 19168
rect 30576 19165 30604 19332
rect 31864 19292 31892 19456
rect 32968 19428 32996 19456
rect 31956 19400 32996 19428
rect 33045 19431 33103 19437
rect 31956 19372 31984 19400
rect 33045 19397 33057 19431
rect 33091 19428 33103 19431
rect 33410 19428 33416 19440
rect 33091 19400 33416 19428
rect 33091 19397 33103 19400
rect 33045 19391 33103 19397
rect 33410 19388 33416 19400
rect 33468 19388 33474 19440
rect 34514 19388 34520 19440
rect 34572 19428 34578 19440
rect 34945 19431 35003 19437
rect 34945 19428 34957 19431
rect 34572 19400 34957 19428
rect 34572 19388 34578 19400
rect 34945 19397 34957 19400
rect 34991 19428 35003 19431
rect 35066 19428 35072 19440
rect 34991 19400 35072 19428
rect 34991 19397 35003 19400
rect 34945 19391 35003 19397
rect 35066 19388 35072 19400
rect 35124 19388 35130 19440
rect 35161 19431 35219 19437
rect 35161 19397 35173 19431
rect 35207 19397 35219 19431
rect 35161 19391 35219 19397
rect 31938 19320 31944 19372
rect 31996 19320 32002 19372
rect 32585 19363 32643 19369
rect 32585 19360 32597 19363
rect 32048 19332 32597 19360
rect 32048 19292 32076 19332
rect 32585 19329 32597 19332
rect 32631 19329 32643 19363
rect 32585 19323 32643 19329
rect 32674 19320 32680 19372
rect 32732 19320 32738 19372
rect 32861 19363 32919 19369
rect 32861 19329 32873 19363
rect 32907 19360 32919 19363
rect 32953 19363 33011 19369
rect 32953 19360 32965 19363
rect 32907 19332 32965 19360
rect 32907 19329 32919 19332
rect 32861 19323 32919 19329
rect 32953 19329 32965 19332
rect 32999 19360 33011 19363
rect 33134 19360 33140 19372
rect 32999 19332 33140 19360
rect 32999 19329 33011 19332
rect 32953 19323 33011 19329
rect 33134 19320 33140 19332
rect 33192 19320 33198 19372
rect 33229 19363 33287 19369
rect 33229 19329 33241 19363
rect 33275 19360 33287 19363
rect 34057 19363 34115 19369
rect 34057 19360 34069 19363
rect 33275 19332 34069 19360
rect 33275 19329 33287 19332
rect 33229 19323 33287 19329
rect 34057 19329 34069 19332
rect 34103 19329 34115 19363
rect 35176 19360 35204 19391
rect 35250 19388 35256 19440
rect 35308 19388 35314 19440
rect 35636 19428 35664 19468
rect 36998 19456 37004 19508
rect 37056 19456 37062 19508
rect 35636 19400 37320 19428
rect 34057 19323 34115 19329
rect 34624 19332 35204 19360
rect 31864 19264 32076 19292
rect 32585 19227 32643 19233
rect 32585 19193 32597 19227
rect 32631 19224 32643 19227
rect 32692 19224 32720 19320
rect 34624 19304 34652 19332
rect 35526 19320 35532 19372
rect 35584 19320 35590 19372
rect 35636 19369 35664 19400
rect 37292 19372 37320 19400
rect 35621 19363 35679 19369
rect 35621 19329 35633 19363
rect 35667 19329 35679 19363
rect 35877 19363 35935 19369
rect 35877 19360 35889 19363
rect 35621 19323 35679 19329
rect 35728 19332 35889 19360
rect 33873 19295 33931 19301
rect 33873 19261 33885 19295
rect 33919 19261 33931 19295
rect 33873 19255 33931 19261
rect 32631 19196 32720 19224
rect 33229 19227 33287 19233
rect 32631 19193 32643 19196
rect 32585 19187 32643 19193
rect 33229 19193 33241 19227
rect 33275 19224 33287 19227
rect 33888 19224 33916 19255
rect 34606 19252 34612 19304
rect 34664 19252 34670 19304
rect 35066 19252 35072 19304
rect 35124 19252 35130 19304
rect 35728 19292 35756 19332
rect 35877 19329 35889 19332
rect 35923 19329 35935 19363
rect 35877 19323 35935 19329
rect 37274 19320 37280 19372
rect 37332 19320 37338 19372
rect 35544 19264 35756 19292
rect 33275 19196 33916 19224
rect 35084 19224 35112 19252
rect 35544 19233 35572 19264
rect 35437 19227 35495 19233
rect 35437 19224 35449 19227
rect 35084 19196 35449 19224
rect 33275 19193 33287 19196
rect 33229 19187 33287 19193
rect 35437 19193 35449 19196
rect 35483 19193 35495 19227
rect 35437 19187 35495 19193
rect 35529 19227 35587 19233
rect 35529 19193 35541 19227
rect 35575 19193 35587 19227
rect 35529 19187 35587 19193
rect 30561 19159 30619 19165
rect 30561 19125 30573 19159
rect 30607 19156 30619 19159
rect 30742 19156 30748 19168
rect 30607 19128 30748 19156
rect 30607 19125 30619 19128
rect 30561 19119 30619 19125
rect 30742 19116 30748 19128
rect 30800 19116 30806 19168
rect 32674 19116 32680 19168
rect 32732 19156 32738 19168
rect 33321 19159 33379 19165
rect 33321 19156 33333 19159
rect 32732 19128 33333 19156
rect 32732 19116 32738 19128
rect 33321 19125 33333 19128
rect 33367 19125 33379 19159
rect 33321 19119 33379 19125
rect 34790 19116 34796 19168
rect 34848 19116 34854 19168
rect 34882 19116 34888 19168
rect 34940 19156 34946 19168
rect 34977 19159 35035 19165
rect 34977 19156 34989 19159
rect 34940 19128 34989 19156
rect 34940 19116 34946 19128
rect 34977 19125 34989 19128
rect 35023 19125 35035 19159
rect 34977 19119 35035 19125
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 13004 18924 13952 18952
rect 12618 18776 12624 18828
rect 12676 18816 12682 18828
rect 12713 18819 12771 18825
rect 12713 18816 12725 18819
rect 12676 18788 12725 18816
rect 12676 18776 12682 18788
rect 12713 18785 12725 18788
rect 12759 18816 12771 18819
rect 13004 18816 13032 18924
rect 13725 18887 13783 18893
rect 13725 18853 13737 18887
rect 13771 18853 13783 18887
rect 13725 18847 13783 18853
rect 12759 18788 13032 18816
rect 13081 18819 13139 18825
rect 12759 18785 12771 18788
rect 12713 18779 12771 18785
rect 13081 18785 13093 18819
rect 13127 18816 13139 18819
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 13127 18788 13553 18816
rect 13127 18785 13139 18788
rect 13081 18779 13139 18785
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 13541 18779 13599 18785
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18816 13691 18819
rect 13740 18816 13768 18847
rect 13679 18788 13768 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9548 18720 9597 18748
rect 9548 18708 9554 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 9600 18680 9628 18711
rect 10594 18708 10600 18760
rect 10652 18708 10658 18760
rect 11054 18708 11060 18760
rect 11112 18708 11118 18760
rect 11514 18708 11520 18760
rect 11572 18708 11578 18760
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18748 12955 18751
rect 12943 18720 13124 18748
rect 12943 18717 12955 18720
rect 12897 18711 12955 18717
rect 11072 18680 11100 18708
rect 9600 18652 11100 18680
rect 13096 18680 13124 18720
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 13924 18757 13952 18924
rect 14274 18912 14280 18964
rect 14332 18952 14338 18964
rect 14921 18955 14979 18961
rect 14921 18952 14933 18955
rect 14332 18924 14933 18952
rect 14332 18912 14338 18924
rect 14921 18921 14933 18924
rect 14967 18921 14979 18955
rect 18598 18952 18604 18964
rect 14921 18915 14979 18921
rect 16500 18924 18604 18952
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 16500 18884 16528 18924
rect 18598 18912 18604 18924
rect 18656 18912 18662 18964
rect 19794 18912 19800 18964
rect 19852 18952 19858 18964
rect 19981 18955 20039 18961
rect 19981 18952 19993 18955
rect 19852 18924 19993 18952
rect 19852 18912 19858 18924
rect 19981 18921 19993 18924
rect 20027 18921 20039 18955
rect 19981 18915 20039 18921
rect 21910 18912 21916 18964
rect 21968 18952 21974 18964
rect 23566 18952 23572 18964
rect 21968 18924 23572 18952
rect 21968 18912 21974 18924
rect 23566 18912 23572 18924
rect 23624 18912 23630 18964
rect 23658 18912 23664 18964
rect 23716 18952 23722 18964
rect 25590 18952 25596 18964
rect 23716 18924 25596 18952
rect 23716 18912 23722 18924
rect 21637 18887 21695 18893
rect 21637 18884 21649 18887
rect 14148 18856 16528 18884
rect 18340 18856 21649 18884
rect 14148 18844 14154 18856
rect 15562 18776 15568 18828
rect 15620 18776 15626 18828
rect 18340 18816 18368 18856
rect 21637 18853 21649 18856
rect 21683 18853 21695 18887
rect 21637 18847 21695 18853
rect 22112 18856 23980 18884
rect 22112 18828 22140 18856
rect 17328 18788 18368 18816
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18717 13783 18751
rect 13725 18711 13783 18717
rect 13909 18751 13967 18757
rect 13909 18717 13921 18751
rect 13955 18717 13967 18751
rect 13909 18711 13967 18717
rect 13446 18680 13452 18692
rect 13096 18652 13452 18680
rect 13096 18624 13124 18652
rect 13446 18640 13452 18652
rect 13504 18680 13510 18692
rect 13740 18680 13768 18711
rect 13504 18652 13768 18680
rect 13504 18640 13510 18652
rect 9490 18572 9496 18624
rect 9548 18572 9554 18624
rect 10134 18572 10140 18624
rect 10192 18612 10198 18624
rect 10413 18615 10471 18621
rect 10413 18612 10425 18615
rect 10192 18584 10425 18612
rect 10192 18572 10198 18584
rect 10413 18581 10425 18584
rect 10459 18581 10471 18615
rect 10413 18575 10471 18581
rect 10962 18572 10968 18624
rect 11020 18572 11026 18624
rect 12158 18572 12164 18624
rect 12216 18572 12222 18624
rect 13078 18572 13084 18624
rect 13136 18572 13142 18624
rect 13170 18572 13176 18624
rect 13228 18572 13234 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 13924 18612 13952 18711
rect 15286 18708 15292 18760
rect 15344 18708 15350 18760
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18748 15439 18751
rect 17328 18748 17356 18788
rect 18414 18776 18420 18828
rect 18472 18816 18478 18828
rect 18877 18819 18935 18825
rect 18877 18816 18889 18819
rect 18472 18788 18889 18816
rect 18472 18776 18478 18788
rect 18877 18785 18889 18788
rect 18923 18785 18935 18819
rect 18877 18779 18935 18785
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18816 19947 18819
rect 20438 18816 20444 18828
rect 19935 18788 20444 18816
rect 19935 18785 19947 18788
rect 19889 18779 19947 18785
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 20548 18788 20852 18816
rect 15427 18720 17356 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 17862 18748 17868 18760
rect 17460 18720 17868 18748
rect 17460 18708 17466 18720
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 18046 18708 18052 18760
rect 18104 18708 18110 18760
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18564 18720 19257 18748
rect 18564 18708 18570 18720
rect 19245 18717 19257 18720
rect 19291 18748 19303 18751
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 19291 18720 20177 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 20165 18717 20177 18720
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 20254 18708 20260 18760
rect 20312 18708 20318 18760
rect 20346 18708 20352 18760
rect 20404 18748 20410 18760
rect 20548 18748 20576 18788
rect 20404 18720 20576 18748
rect 20625 18751 20683 18757
rect 20404 18708 20410 18720
rect 20625 18717 20637 18751
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 17160 18683 17218 18689
rect 17160 18649 17172 18683
rect 17206 18680 17218 18683
rect 17497 18683 17555 18689
rect 17497 18680 17509 18683
rect 17206 18652 17509 18680
rect 17206 18649 17218 18652
rect 17160 18643 17218 18649
rect 17497 18649 17509 18652
rect 17543 18649 17555 18683
rect 17497 18643 17555 18649
rect 17972 18652 20300 18680
rect 17972 18624 18000 18652
rect 13780 18584 13952 18612
rect 13780 18572 13786 18584
rect 16022 18572 16028 18624
rect 16080 18572 16086 18624
rect 17954 18572 17960 18624
rect 18012 18572 18018 18624
rect 18322 18572 18328 18624
rect 18380 18572 18386 18624
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 20162 18612 20168 18624
rect 19392 18584 20168 18612
rect 19392 18572 19398 18584
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 20272 18612 20300 18652
rect 20438 18640 20444 18692
rect 20496 18689 20502 18692
rect 20496 18683 20525 18689
rect 20513 18649 20525 18683
rect 20496 18643 20525 18649
rect 20496 18640 20502 18643
rect 20640 18612 20668 18711
rect 20714 18708 20720 18760
rect 20772 18708 20778 18760
rect 20824 18680 20852 18788
rect 22094 18776 22100 18828
rect 22152 18776 22158 18828
rect 22278 18776 22284 18828
rect 22336 18776 22342 18828
rect 20898 18708 20904 18760
rect 20956 18708 20962 18760
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18748 22063 18751
rect 22830 18748 22836 18760
rect 22051 18720 22836 18748
rect 22051 18717 22063 18720
rect 22005 18711 22063 18717
rect 22830 18708 22836 18720
rect 22888 18708 22894 18760
rect 23124 18757 23152 18856
rect 23569 18819 23627 18825
rect 23569 18785 23581 18819
rect 23615 18816 23627 18819
rect 23753 18819 23811 18825
rect 23753 18816 23765 18819
rect 23615 18788 23765 18816
rect 23615 18785 23627 18788
rect 23569 18779 23627 18785
rect 23753 18785 23765 18788
rect 23799 18785 23811 18819
rect 23753 18779 23811 18785
rect 22925 18751 22983 18757
rect 22925 18717 22937 18751
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 23109 18751 23167 18757
rect 23109 18717 23121 18751
rect 23155 18717 23167 18751
rect 23109 18711 23167 18717
rect 22646 18680 22652 18692
rect 20824 18652 22652 18680
rect 22646 18640 22652 18652
rect 22704 18640 22710 18692
rect 20809 18615 20867 18621
rect 20809 18612 20821 18615
rect 20272 18584 20821 18612
rect 20809 18581 20821 18584
rect 20855 18581 20867 18615
rect 20809 18575 20867 18581
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22940 18612 22968 18711
rect 23198 18708 23204 18760
rect 23256 18708 23262 18760
rect 23382 18708 23388 18760
rect 23440 18708 23446 18760
rect 23952 18757 23980 18856
rect 24121 18819 24179 18825
rect 24121 18785 24133 18819
rect 24167 18816 24179 18819
rect 25038 18816 25044 18828
rect 24167 18788 25044 18816
rect 24167 18785 24179 18788
rect 24121 18779 24179 18785
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18717 23719 18751
rect 23661 18711 23719 18717
rect 23937 18751 23995 18757
rect 23937 18717 23949 18751
rect 23983 18717 23995 18751
rect 23937 18711 23995 18717
rect 23017 18683 23075 18689
rect 23017 18649 23029 18683
rect 23063 18680 23075 18683
rect 23676 18680 23704 18711
rect 23063 18652 23704 18680
rect 23063 18649 23075 18652
rect 23017 18643 23075 18649
rect 24136 18612 24164 18779
rect 25038 18776 25044 18788
rect 25096 18776 25102 18828
rect 25148 18748 25176 18924
rect 25590 18912 25596 18924
rect 25648 18912 25654 18964
rect 25682 18912 25688 18964
rect 25740 18952 25746 18964
rect 25961 18955 26019 18961
rect 25961 18952 25973 18955
rect 25740 18924 25973 18952
rect 25740 18912 25746 18924
rect 25961 18921 25973 18924
rect 26007 18921 26019 18955
rect 25961 18915 26019 18921
rect 29914 18912 29920 18964
rect 29972 18952 29978 18964
rect 30469 18955 30527 18961
rect 30469 18952 30481 18955
rect 29972 18924 30481 18952
rect 29972 18912 29978 18924
rect 28718 18844 28724 18896
rect 28776 18844 28782 18896
rect 27706 18776 27712 18828
rect 27764 18816 27770 18828
rect 28353 18819 28411 18825
rect 28353 18816 28365 18819
rect 27764 18788 28365 18816
rect 27764 18776 27770 18788
rect 28353 18785 28365 18788
rect 28399 18785 28411 18819
rect 28353 18779 28411 18785
rect 28537 18819 28595 18825
rect 28537 18785 28549 18819
rect 28583 18816 28595 18819
rect 28810 18816 28816 18828
rect 28583 18788 28816 18816
rect 28583 18785 28595 18788
rect 28537 18779 28595 18785
rect 28810 18776 28816 18788
rect 28868 18816 28874 18828
rect 28868 18788 29040 18816
rect 28868 18776 28874 18788
rect 25590 18748 25596 18760
rect 25148 18720 25596 18748
rect 25590 18708 25596 18720
rect 25648 18748 25654 18760
rect 25777 18751 25835 18757
rect 25777 18748 25789 18751
rect 25648 18720 25789 18748
rect 25648 18708 25654 18720
rect 25777 18717 25789 18720
rect 25823 18717 25835 18751
rect 25777 18711 25835 18717
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18748 26019 18751
rect 26053 18751 26111 18757
rect 26053 18748 26065 18751
rect 26007 18720 26065 18748
rect 26007 18717 26019 18720
rect 25961 18711 26019 18717
rect 26053 18717 26065 18720
rect 26099 18717 26111 18751
rect 26053 18711 26111 18717
rect 26602 18708 26608 18760
rect 26660 18708 26666 18760
rect 26881 18751 26939 18757
rect 26881 18717 26893 18751
rect 26927 18748 26939 18751
rect 28074 18748 28080 18760
rect 26927 18720 28080 18748
rect 26927 18717 26939 18720
rect 26881 18711 26939 18717
rect 25866 18640 25872 18692
rect 25924 18680 25930 18692
rect 26896 18680 26924 18711
rect 28074 18708 28080 18720
rect 28132 18708 28138 18760
rect 29012 18757 29040 18788
rect 28629 18751 28687 18757
rect 28629 18717 28641 18751
rect 28675 18748 28687 18751
rect 28997 18751 29055 18757
rect 28675 18720 28948 18748
rect 28675 18717 28687 18720
rect 28629 18711 28687 18717
rect 25924 18652 26924 18680
rect 28353 18683 28411 18689
rect 25924 18640 25930 18652
rect 28353 18649 28365 18683
rect 28399 18680 28411 18683
rect 28721 18683 28779 18689
rect 28721 18680 28733 18683
rect 28399 18652 28733 18680
rect 28399 18649 28411 18652
rect 28353 18643 28411 18649
rect 28721 18649 28733 18652
rect 28767 18649 28779 18683
rect 28721 18643 28779 18649
rect 22152 18584 24164 18612
rect 26973 18615 27031 18621
rect 22152 18572 22158 18584
rect 26973 18581 26985 18615
rect 27019 18612 27031 18615
rect 27062 18612 27068 18624
rect 27019 18584 27068 18612
rect 27019 18581 27031 18584
rect 26973 18575 27031 18581
rect 27062 18572 27068 18584
rect 27120 18572 27126 18624
rect 28920 18621 28948 18720
rect 28997 18717 29009 18751
rect 29043 18717 29055 18751
rect 28997 18711 29055 18717
rect 29012 18680 29040 18711
rect 29178 18708 29184 18760
rect 29236 18748 29242 18760
rect 30116 18757 30144 18924
rect 30469 18921 30481 18924
rect 30515 18921 30527 18955
rect 30469 18915 30527 18921
rect 31386 18912 31392 18964
rect 31444 18952 31450 18964
rect 31444 18924 31708 18952
rect 31444 18912 31450 18924
rect 30558 18884 30564 18896
rect 30208 18856 30564 18884
rect 30101 18751 30159 18757
rect 30101 18748 30113 18751
rect 29236 18720 30113 18748
rect 29236 18708 29242 18720
rect 30101 18717 30113 18720
rect 30147 18717 30159 18751
rect 30101 18711 30159 18717
rect 29638 18680 29644 18692
rect 29012 18652 29644 18680
rect 29638 18640 29644 18652
rect 29696 18680 29702 18692
rect 30208 18680 30236 18856
rect 30558 18844 30564 18856
rect 30616 18844 30622 18896
rect 30653 18887 30711 18893
rect 30653 18853 30665 18887
rect 30699 18884 30711 18887
rect 30834 18884 30840 18896
rect 30699 18856 30840 18884
rect 30699 18853 30711 18856
rect 30653 18847 30711 18853
rect 30834 18844 30840 18856
rect 30892 18884 30898 18896
rect 31573 18887 31631 18893
rect 31573 18884 31585 18887
rect 30892 18856 31585 18884
rect 30892 18844 30898 18856
rect 31573 18853 31585 18856
rect 31619 18853 31631 18887
rect 31573 18847 31631 18853
rect 31680 18828 31708 18924
rect 31754 18912 31760 18964
rect 31812 18952 31818 18964
rect 31941 18955 31999 18961
rect 31941 18952 31953 18955
rect 31812 18924 31953 18952
rect 31812 18912 31818 18924
rect 31941 18921 31953 18924
rect 31987 18921 31999 18955
rect 33962 18952 33968 18964
rect 31941 18915 31999 18921
rect 32784 18924 33968 18952
rect 32784 18893 32812 18924
rect 33962 18912 33968 18924
rect 34020 18952 34026 18964
rect 34333 18955 34391 18961
rect 34020 18924 34284 18952
rect 34020 18912 34026 18924
rect 32769 18887 32827 18893
rect 32769 18853 32781 18887
rect 32815 18853 32827 18887
rect 34256 18884 34284 18924
rect 34333 18921 34345 18955
rect 34379 18952 34391 18955
rect 34606 18952 34612 18964
rect 34379 18924 34612 18952
rect 34379 18921 34391 18924
rect 34333 18915 34391 18921
rect 34606 18912 34612 18924
rect 34664 18912 34670 18964
rect 34974 18884 34980 18896
rect 34256 18856 34980 18884
rect 32769 18847 32827 18853
rect 34974 18844 34980 18856
rect 35032 18884 35038 18896
rect 36722 18884 36728 18896
rect 35032 18856 36728 18884
rect 35032 18844 35038 18856
rect 36722 18844 36728 18856
rect 36780 18844 36786 18896
rect 30742 18776 30748 18828
rect 30800 18776 30806 18828
rect 31662 18776 31668 18828
rect 31720 18816 31726 18828
rect 31720 18788 31800 18816
rect 31720 18776 31726 18788
rect 31772 18757 31800 18788
rect 32582 18776 32588 18828
rect 32640 18776 32646 18828
rect 32950 18776 32956 18828
rect 33008 18776 33014 18828
rect 31389 18751 31447 18757
rect 31389 18717 31401 18751
rect 31435 18748 31447 18751
rect 31481 18751 31539 18757
rect 31481 18748 31493 18751
rect 31435 18720 31493 18748
rect 31435 18717 31447 18720
rect 31389 18711 31447 18717
rect 31481 18717 31493 18720
rect 31527 18717 31539 18751
rect 31481 18711 31539 18717
rect 31757 18751 31815 18757
rect 31757 18717 31769 18751
rect 31803 18717 31815 18751
rect 31757 18711 31815 18717
rect 32674 18708 32680 18760
rect 32732 18708 32738 18760
rect 32861 18751 32919 18757
rect 32861 18717 32873 18751
rect 32907 18717 32919 18751
rect 32861 18711 32919 18717
rect 29696 18652 30236 18680
rect 29696 18640 29702 18652
rect 28905 18615 28963 18621
rect 28905 18581 28917 18615
rect 28951 18612 28963 18615
rect 29549 18615 29607 18621
rect 29549 18612 29561 18615
rect 28951 18584 29561 18612
rect 28951 18581 28963 18584
rect 28905 18575 28963 18581
rect 29549 18581 29561 18584
rect 29595 18612 29607 18615
rect 29730 18612 29736 18624
rect 29595 18584 29736 18612
rect 29595 18581 29607 18584
rect 29549 18575 29607 18581
rect 29730 18572 29736 18584
rect 29788 18572 29794 18624
rect 30208 18612 30236 18652
rect 30282 18640 30288 18692
rect 30340 18640 30346 18692
rect 32692 18680 32720 18708
rect 32876 18680 32904 18711
rect 34790 18708 34796 18760
rect 34848 18708 34854 18760
rect 37182 18708 37188 18760
rect 37240 18708 37246 18760
rect 37461 18751 37519 18757
rect 37461 18717 37473 18751
rect 37507 18717 37519 18751
rect 37461 18711 37519 18717
rect 37645 18751 37703 18757
rect 37645 18717 37657 18751
rect 37691 18748 37703 18751
rect 37921 18751 37979 18757
rect 37921 18748 37933 18751
rect 37691 18720 37933 18748
rect 37691 18717 37703 18720
rect 37645 18711 37703 18717
rect 37921 18717 37933 18720
rect 37967 18717 37979 18751
rect 37921 18711 37979 18717
rect 38473 18751 38531 18757
rect 38473 18717 38485 18751
rect 38519 18717 38531 18751
rect 38473 18711 38531 18717
rect 32692 18652 32904 18680
rect 33198 18683 33256 18689
rect 33198 18649 33210 18683
rect 33244 18649 33256 18683
rect 37476 18680 37504 18711
rect 38286 18680 38292 18692
rect 33198 18643 33256 18649
rect 36648 18652 38292 18680
rect 30485 18615 30543 18621
rect 30485 18612 30497 18615
rect 30208 18584 30497 18612
rect 30485 18581 30497 18584
rect 30531 18581 30543 18615
rect 30485 18575 30543 18581
rect 32861 18615 32919 18621
rect 32861 18581 32873 18615
rect 32907 18612 32919 18615
rect 33213 18612 33241 18643
rect 36648 18624 36676 18652
rect 38286 18640 38292 18652
rect 38344 18640 38350 18692
rect 38488 18624 38516 18711
rect 32907 18584 33241 18612
rect 32907 18581 32919 18584
rect 32861 18575 32919 18581
rect 36630 18572 36636 18624
rect 36688 18572 36694 18624
rect 36998 18572 37004 18624
rect 37056 18572 37062 18624
rect 38470 18572 38476 18624
rect 38528 18572 38534 18624
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 7926 18408 7932 18420
rect 7760 18380 7932 18408
rect 7760 18284 7788 18380
rect 7926 18368 7932 18380
rect 7984 18408 7990 18420
rect 10870 18408 10876 18420
rect 7984 18380 10876 18408
rect 7984 18368 7990 18380
rect 9490 18340 9496 18352
rect 9246 18312 9496 18340
rect 9490 18300 9496 18312
rect 9548 18300 9554 18352
rect 7742 18232 7748 18284
rect 7800 18232 7806 18284
rect 9600 18281 9628 18380
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 11333 18411 11391 18417
rect 11333 18377 11345 18411
rect 11379 18408 11391 18411
rect 11514 18408 11520 18420
rect 11379 18380 11520 18408
rect 11379 18377 11391 18380
rect 11333 18371 11391 18377
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 12158 18368 12164 18420
rect 12216 18368 12222 18420
rect 13170 18368 13176 18420
rect 13228 18408 13234 18420
rect 13228 18380 13492 18408
rect 13228 18368 13234 18380
rect 9861 18343 9919 18349
rect 9861 18309 9873 18343
rect 9907 18340 9919 18343
rect 10134 18340 10140 18352
rect 9907 18312 10140 18340
rect 9907 18309 9919 18312
rect 9861 18303 9919 18309
rect 10134 18300 10140 18312
rect 10192 18300 10198 18352
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 10962 18232 10968 18284
rect 11020 18232 11026 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18272 11759 18275
rect 12176 18272 12204 18368
rect 13354 18340 13360 18352
rect 11747 18244 12204 18272
rect 12406 18312 13360 18340
rect 11747 18241 11759 18244
rect 11701 18235 11759 18241
rect 8021 18207 8079 18213
rect 8021 18173 8033 18207
rect 8067 18204 8079 18207
rect 8478 18204 8484 18216
rect 8067 18176 8484 18204
rect 8067 18173 8079 18176
rect 8021 18167 8079 18173
rect 8478 18164 8484 18176
rect 8536 18164 8542 18216
rect 11532 18204 11560 18235
rect 12406 18204 12434 18312
rect 13354 18300 13360 18312
rect 13412 18300 13418 18352
rect 13464 18349 13492 18380
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 13780 18380 15240 18408
rect 13780 18368 13786 18380
rect 13449 18343 13507 18349
rect 13449 18309 13461 18343
rect 13495 18309 13507 18343
rect 13449 18303 13507 18309
rect 14458 18300 14464 18352
rect 14516 18300 14522 18352
rect 15212 18349 15240 18380
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 15528 18380 17172 18408
rect 15528 18368 15534 18380
rect 15197 18343 15255 18349
rect 15197 18309 15209 18343
rect 15243 18340 15255 18343
rect 15243 18312 17080 18340
rect 15243 18309 15255 18312
rect 15197 18303 15255 18309
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 13170 18272 13176 18284
rect 12584 18244 13176 18272
rect 12584 18232 12590 18244
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 11532 18176 12434 18204
rect 11808 18080 11836 18176
rect 15562 18096 15568 18148
rect 15620 18136 15626 18148
rect 17052 18136 17080 18312
rect 17144 18272 17172 18380
rect 17310 18368 17316 18420
rect 17368 18368 17374 18420
rect 17497 18411 17555 18417
rect 17497 18377 17509 18411
rect 17543 18408 17555 18411
rect 18046 18408 18052 18420
rect 17543 18380 18052 18408
rect 17543 18377 17555 18380
rect 17497 18371 17555 18377
rect 18046 18368 18052 18380
rect 18104 18368 18110 18420
rect 18322 18368 18328 18420
rect 18380 18368 18386 18420
rect 18598 18408 18604 18420
rect 18524 18380 18604 18408
rect 17328 18340 17356 18368
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 17328 18312 18245 18340
rect 18233 18309 18245 18312
rect 18279 18309 18291 18343
rect 18233 18303 18291 18309
rect 17494 18272 17500 18284
rect 17144 18244 17500 18272
rect 17494 18232 17500 18244
rect 17552 18272 17558 18284
rect 17681 18275 17739 18281
rect 17681 18272 17693 18275
rect 17552 18244 17693 18272
rect 17552 18232 17558 18244
rect 17681 18241 17693 18244
rect 17727 18241 17739 18275
rect 17681 18235 17739 18241
rect 17770 18232 17776 18284
rect 17828 18232 17834 18284
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18241 17923 18275
rect 17865 18235 17923 18241
rect 17218 18164 17224 18216
rect 17276 18164 17282 18216
rect 17880 18204 17908 18235
rect 17954 18232 17960 18284
rect 18012 18281 18018 18284
rect 18012 18275 18041 18281
rect 18029 18241 18041 18275
rect 18012 18235 18041 18241
rect 18141 18275 18199 18281
rect 18141 18241 18153 18275
rect 18187 18272 18199 18275
rect 18340 18272 18368 18368
rect 18524 18281 18552 18380
rect 18598 18368 18604 18380
rect 18656 18408 18662 18420
rect 19426 18408 19432 18420
rect 18656 18380 19432 18408
rect 18656 18368 18662 18380
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 19521 18411 19579 18417
rect 19521 18377 19533 18411
rect 19567 18408 19579 18411
rect 20438 18408 20444 18420
rect 19567 18380 20444 18408
rect 19567 18377 19579 18380
rect 19521 18371 19579 18377
rect 19334 18340 19340 18352
rect 18616 18312 19340 18340
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 18187 18244 18429 18272
rect 18187 18241 18199 18244
rect 18141 18235 18199 18241
rect 18417 18241 18429 18244
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 18509 18275 18567 18281
rect 18509 18241 18521 18275
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 18012 18232 18018 18235
rect 18616 18204 18644 18312
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 18690 18232 18696 18284
rect 18748 18232 18754 18284
rect 18785 18275 18843 18281
rect 18785 18241 18797 18275
rect 18831 18272 18843 18275
rect 19536 18272 19564 18371
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 22646 18368 22652 18420
rect 22704 18368 22710 18420
rect 23198 18368 23204 18420
rect 23256 18408 23262 18420
rect 23256 18380 23336 18408
rect 23256 18368 23262 18380
rect 20073 18343 20131 18349
rect 20073 18309 20085 18343
rect 20119 18340 20131 18343
rect 20714 18340 20720 18352
rect 20119 18312 20720 18340
rect 20119 18309 20131 18312
rect 20073 18303 20131 18309
rect 20714 18300 20720 18312
rect 20772 18300 20778 18352
rect 20806 18300 20812 18352
rect 20864 18340 20870 18352
rect 23308 18349 23336 18380
rect 28718 18368 28724 18420
rect 28776 18368 28782 18420
rect 29178 18368 29184 18420
rect 29236 18368 29242 18420
rect 29549 18411 29607 18417
rect 29549 18377 29561 18411
rect 29595 18408 29607 18411
rect 30282 18408 30288 18420
rect 29595 18380 30288 18408
rect 29595 18377 29607 18380
rect 29549 18371 29607 18377
rect 30282 18368 30288 18380
rect 30340 18368 30346 18420
rect 36722 18368 36728 18420
rect 36780 18368 36786 18420
rect 36998 18368 37004 18420
rect 37056 18368 37062 18420
rect 21177 18343 21235 18349
rect 21177 18340 21189 18343
rect 20864 18312 21189 18340
rect 20864 18300 20870 18312
rect 21177 18309 21189 18312
rect 21223 18309 21235 18343
rect 21177 18303 21235 18309
rect 23293 18343 23351 18349
rect 23293 18309 23305 18343
rect 23339 18309 23351 18343
rect 23293 18303 23351 18309
rect 25038 18300 25044 18352
rect 25096 18300 25102 18352
rect 28068 18343 28126 18349
rect 28068 18309 28080 18343
rect 28114 18340 28126 18343
rect 28736 18340 28764 18368
rect 28114 18312 28764 18340
rect 30684 18343 30742 18349
rect 28114 18309 28126 18312
rect 28068 18303 28126 18309
rect 30684 18309 30696 18343
rect 30730 18340 30742 18343
rect 31021 18343 31079 18349
rect 31021 18340 31033 18343
rect 30730 18312 31033 18340
rect 30730 18309 30742 18312
rect 30684 18303 30742 18309
rect 31021 18309 31033 18312
rect 31067 18309 31079 18343
rect 31021 18303 31079 18309
rect 34974 18300 34980 18352
rect 35032 18300 35038 18352
rect 35452 18312 36400 18340
rect 18831 18244 19564 18272
rect 19981 18275 20039 18281
rect 18831 18241 18843 18244
rect 18785 18235 18843 18241
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20441 18275 20499 18281
rect 20027 18244 20116 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20088 18216 20116 18244
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 21453 18275 21511 18281
rect 21453 18272 21465 18275
rect 20441 18235 20499 18241
rect 21008 18244 21465 18272
rect 17880 18176 18644 18204
rect 18966 18164 18972 18216
rect 19024 18164 19030 18216
rect 19334 18164 19340 18216
rect 19392 18164 19398 18216
rect 20070 18164 20076 18216
rect 20128 18164 20134 18216
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 19352 18136 19380 18164
rect 15620 18108 16896 18136
rect 17052 18108 19380 18136
rect 15620 18096 15626 18108
rect 9493 18071 9551 18077
rect 9493 18037 9505 18071
rect 9539 18068 9551 18071
rect 9858 18068 9864 18080
rect 9539 18040 9864 18068
rect 9539 18037 9551 18040
rect 9493 18031 9551 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 11606 18028 11612 18080
rect 11664 18028 11670 18080
rect 11790 18028 11796 18080
rect 11848 18028 11854 18080
rect 13446 18028 13452 18080
rect 13504 18068 13510 18080
rect 15470 18068 15476 18080
rect 13504 18040 15476 18068
rect 13504 18028 13510 18040
rect 15470 18028 15476 18040
rect 15528 18028 15534 18080
rect 16669 18071 16727 18077
rect 16669 18037 16681 18071
rect 16715 18068 16727 18071
rect 16758 18068 16764 18080
rect 16715 18040 16764 18068
rect 16715 18037 16727 18040
rect 16669 18031 16727 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 16868 18068 16896 18108
rect 19426 18096 19432 18148
rect 19484 18136 19490 18148
rect 19613 18139 19671 18145
rect 19613 18136 19625 18139
rect 19484 18108 19625 18136
rect 19484 18096 19490 18108
rect 19613 18105 19625 18108
rect 19659 18105 19671 18139
rect 19613 18099 19671 18105
rect 18138 18068 18144 18080
rect 16868 18040 18144 18068
rect 18138 18028 18144 18040
rect 18196 18068 18202 18080
rect 20180 18068 20208 18167
rect 20456 18136 20484 18235
rect 21008 18216 21036 18244
rect 21453 18241 21465 18244
rect 21499 18272 21511 18275
rect 21910 18272 21916 18284
rect 21499 18244 21916 18272
rect 21499 18241 21511 18244
rect 21453 18235 21511 18241
rect 21910 18232 21916 18244
rect 21968 18232 21974 18284
rect 22557 18275 22615 18281
rect 22557 18241 22569 18275
rect 22603 18241 22615 18275
rect 22557 18235 22615 18241
rect 20990 18164 20996 18216
rect 21048 18164 21054 18216
rect 21545 18207 21603 18213
rect 21545 18173 21557 18207
rect 21591 18204 21603 18207
rect 21818 18204 21824 18216
rect 21591 18176 21824 18204
rect 21591 18173 21603 18176
rect 21545 18167 21603 18173
rect 21818 18164 21824 18176
rect 21876 18204 21882 18216
rect 22572 18204 22600 18235
rect 22922 18232 22928 18284
rect 22980 18272 22986 18284
rect 23017 18275 23075 18281
rect 23017 18272 23029 18275
rect 22980 18244 23029 18272
rect 22980 18232 22986 18244
rect 23017 18241 23029 18244
rect 23063 18241 23075 18275
rect 23017 18235 23075 18241
rect 24394 18232 24400 18284
rect 24452 18232 24458 18284
rect 25498 18232 25504 18284
rect 25556 18232 25562 18284
rect 25682 18232 25688 18284
rect 25740 18272 25746 18284
rect 25777 18275 25835 18281
rect 25777 18272 25789 18275
rect 25740 18244 25789 18272
rect 25740 18232 25746 18244
rect 25777 18241 25789 18244
rect 25823 18241 25835 18275
rect 25777 18235 25835 18241
rect 25869 18275 25927 18281
rect 25869 18241 25881 18275
rect 25915 18272 25927 18275
rect 25958 18272 25964 18284
rect 25915 18244 25964 18272
rect 25915 18241 25927 18244
rect 25869 18235 25927 18241
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 26053 18275 26111 18281
rect 26053 18241 26065 18275
rect 26099 18272 26111 18275
rect 26973 18275 27031 18281
rect 26973 18272 26985 18275
rect 26099 18244 26985 18272
rect 26099 18241 26111 18244
rect 26053 18235 26111 18241
rect 26973 18241 26985 18244
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 27522 18232 27528 18284
rect 27580 18272 27586 18284
rect 27801 18275 27859 18281
rect 27801 18272 27813 18275
rect 27580 18244 27813 18272
rect 27580 18232 27586 18244
rect 27801 18241 27813 18244
rect 27847 18241 27859 18275
rect 27801 18235 27859 18241
rect 30929 18275 30987 18281
rect 30929 18241 30941 18275
rect 30975 18272 30987 18275
rect 31938 18272 31944 18284
rect 30975 18244 31944 18272
rect 30975 18241 30987 18244
rect 30929 18235 30987 18241
rect 31938 18232 31944 18244
rect 31996 18232 32002 18284
rect 34992 18272 35020 18300
rect 35069 18275 35127 18281
rect 35069 18272 35081 18275
rect 34992 18244 35081 18272
rect 35069 18241 35081 18244
rect 35115 18241 35127 18275
rect 35069 18235 35127 18241
rect 35161 18275 35219 18281
rect 35161 18241 35173 18275
rect 35207 18241 35219 18275
rect 35161 18235 35219 18241
rect 21876 18176 24348 18204
rect 21876 18164 21882 18176
rect 20898 18136 20904 18148
rect 20456 18108 20904 18136
rect 20898 18096 20904 18108
rect 20956 18136 20962 18148
rect 24320 18136 24348 18176
rect 26602 18164 26608 18216
rect 26660 18164 26666 18216
rect 27614 18164 27620 18216
rect 27672 18164 27678 18216
rect 31202 18164 31208 18216
rect 31260 18204 31266 18216
rect 31573 18207 31631 18213
rect 31573 18204 31585 18207
rect 31260 18176 31585 18204
rect 31260 18164 31266 18176
rect 31573 18173 31585 18176
rect 31619 18173 31631 18207
rect 35176 18204 35204 18235
rect 35342 18232 35348 18284
rect 35400 18232 35406 18284
rect 35452 18281 35480 18312
rect 36372 18284 36400 18312
rect 36630 18300 36636 18352
rect 36688 18300 36694 18352
rect 36740 18340 36768 18368
rect 37016 18340 37044 18368
rect 37522 18343 37580 18349
rect 37522 18340 37534 18343
rect 36740 18312 36865 18340
rect 37016 18312 37534 18340
rect 35437 18275 35495 18281
rect 35437 18241 35449 18275
rect 35483 18241 35495 18275
rect 35437 18235 35495 18241
rect 36078 18232 36084 18284
rect 36136 18232 36142 18284
rect 36354 18232 36360 18284
rect 36412 18232 36418 18284
rect 36446 18232 36452 18284
rect 36504 18272 36510 18284
rect 36504 18244 36676 18272
rect 36504 18232 36510 18244
rect 36096 18204 36124 18232
rect 35176 18176 36124 18204
rect 31573 18167 31631 18173
rect 25866 18136 25872 18148
rect 20956 18108 22232 18136
rect 24320 18108 25872 18136
rect 20956 18096 20962 18108
rect 22204 18077 22232 18108
rect 25866 18096 25872 18108
rect 25924 18096 25930 18148
rect 26053 18139 26111 18145
rect 26053 18105 26065 18139
rect 26099 18136 26111 18139
rect 26620 18136 26648 18164
rect 26099 18108 26648 18136
rect 26099 18105 26111 18108
rect 26053 18099 26111 18105
rect 18196 18040 20208 18068
rect 22189 18071 22247 18077
rect 18196 18028 18202 18040
rect 22189 18037 22201 18071
rect 22235 18068 22247 18071
rect 23290 18068 23296 18080
rect 22235 18040 23296 18068
rect 22235 18037 22247 18040
rect 22189 18031 22247 18037
rect 23290 18028 23296 18040
rect 23348 18028 23354 18080
rect 25317 18071 25375 18077
rect 25317 18037 25329 18071
rect 25363 18068 25375 18071
rect 25406 18068 25412 18080
rect 25363 18040 25412 18068
rect 25363 18037 25375 18040
rect 25317 18031 25375 18037
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 25590 18028 25596 18080
rect 25648 18068 25654 18080
rect 31018 18068 31024 18080
rect 25648 18040 31024 18068
rect 25648 18028 25654 18040
rect 31018 18028 31024 18040
rect 31076 18028 31082 18080
rect 34790 18028 34796 18080
rect 34848 18068 34854 18080
rect 34885 18071 34943 18077
rect 34885 18068 34897 18071
rect 34848 18040 34897 18068
rect 34848 18028 34854 18040
rect 34885 18037 34897 18040
rect 34931 18037 34943 18071
rect 36648 18068 36676 18244
rect 36722 18232 36728 18284
rect 36780 18232 36786 18284
rect 36837 18281 36865 18312
rect 37522 18309 37534 18312
rect 37568 18309 37580 18343
rect 37522 18303 37580 18309
rect 36906 18281 36912 18284
rect 36837 18275 36912 18281
rect 36837 18244 36873 18275
rect 36861 18241 36873 18244
rect 36907 18241 36912 18275
rect 36861 18235 36912 18241
rect 36906 18232 36912 18235
rect 36964 18232 36970 18284
rect 37182 18232 37188 18284
rect 37240 18232 37246 18284
rect 37274 18232 37280 18284
rect 37332 18232 37338 18284
rect 37001 18139 37059 18145
rect 37001 18105 37013 18139
rect 37047 18136 37059 18139
rect 37200 18136 37228 18232
rect 37047 18108 37228 18136
rect 37047 18105 37059 18108
rect 37001 18099 37059 18105
rect 38470 18068 38476 18080
rect 36648 18040 38476 18068
rect 34885 18031 34943 18037
rect 38470 18028 38476 18040
rect 38528 18068 38534 18080
rect 38657 18071 38715 18077
rect 38657 18068 38669 18071
rect 38528 18040 38669 18068
rect 38528 18028 38534 18040
rect 38657 18037 38669 18040
rect 38703 18037 38715 18071
rect 38657 18031 38715 18037
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 8478 17824 8484 17876
rect 8536 17864 8542 17876
rect 8941 17867 8999 17873
rect 8941 17864 8953 17867
rect 8536 17836 8953 17864
rect 8536 17824 8542 17836
rect 8941 17833 8953 17836
rect 8987 17833 8999 17867
rect 8941 17827 8999 17833
rect 10505 17867 10563 17873
rect 10505 17833 10517 17867
rect 10551 17864 10563 17867
rect 10594 17864 10600 17876
rect 10551 17836 10600 17864
rect 10551 17833 10563 17836
rect 10505 17827 10563 17833
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 10870 17824 10876 17876
rect 10928 17864 10934 17876
rect 10928 17836 11376 17864
rect 10928 17824 10934 17836
rect 11348 17737 11376 17836
rect 13078 17824 13084 17876
rect 13136 17873 13142 17876
rect 13136 17867 13185 17873
rect 13136 17833 13139 17867
rect 13173 17833 13185 17867
rect 13136 17827 13185 17833
rect 13136 17824 13142 17827
rect 20714 17824 20720 17876
rect 20772 17824 20778 17876
rect 22278 17864 22284 17876
rect 21376 17836 22284 17864
rect 19889 17799 19947 17805
rect 19889 17765 19901 17799
rect 19935 17796 19947 17799
rect 20346 17796 20352 17808
rect 19935 17768 20352 17796
rect 19935 17765 19947 17768
rect 19889 17759 19947 17765
rect 20346 17756 20352 17768
rect 20404 17756 20410 17808
rect 11149 17731 11207 17737
rect 11149 17697 11161 17731
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17697 11391 17731
rect 11333 17691 11391 17697
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 11164 17660 11192 17691
rect 11514 17688 11520 17740
rect 11572 17688 11578 17740
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 11701 17731 11759 17737
rect 11701 17728 11713 17731
rect 11664 17700 11713 17728
rect 11664 17688 11670 17700
rect 11701 17697 11713 17700
rect 11747 17697 11759 17731
rect 11701 17691 11759 17697
rect 13170 17688 13176 17740
rect 13228 17728 13234 17740
rect 13722 17728 13728 17740
rect 13228 17700 13728 17728
rect 13228 17688 13234 17700
rect 13722 17688 13728 17700
rect 13780 17728 13786 17740
rect 15102 17728 15108 17740
rect 13780 17700 15108 17728
rect 13780 17688 13786 17700
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 21376 17737 21404 17836
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 24394 17824 24400 17876
rect 24452 17864 24458 17876
rect 24489 17867 24547 17873
rect 24489 17864 24501 17867
rect 24452 17836 24501 17864
rect 24452 17824 24458 17836
rect 24489 17833 24501 17836
rect 24535 17833 24547 17867
rect 26513 17867 26571 17873
rect 24489 17827 24547 17833
rect 25148 17836 26188 17864
rect 19429 17731 19487 17737
rect 19429 17728 19441 17731
rect 19392 17700 19441 17728
rect 19392 17688 19398 17700
rect 19429 17697 19441 17700
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 21361 17731 21419 17737
rect 21361 17697 21373 17731
rect 21407 17697 21419 17731
rect 21361 17691 21419 17697
rect 21634 17688 21640 17740
rect 21692 17688 21698 17740
rect 21818 17688 21824 17740
rect 21876 17688 21882 17740
rect 22925 17731 22983 17737
rect 22925 17728 22937 17731
rect 22020 17700 22937 17728
rect 11532 17660 11560 17688
rect 11164 17632 11560 17660
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 17957 17663 18015 17669
rect 17957 17660 17969 17663
rect 17920 17632 17969 17660
rect 17920 17620 17926 17632
rect 17957 17629 17969 17632
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 18230 17620 18236 17672
rect 18288 17620 18294 17672
rect 21652 17660 21680 17688
rect 22020 17669 22048 17700
rect 22925 17697 22937 17700
rect 22971 17697 22983 17731
rect 22925 17691 22983 17697
rect 23014 17688 23020 17740
rect 23072 17728 23078 17740
rect 23290 17728 23296 17740
rect 23072 17700 23296 17728
rect 23072 17688 23078 17700
rect 23290 17688 23296 17700
rect 23348 17728 23354 17740
rect 23569 17731 23627 17737
rect 23348 17700 23428 17728
rect 23348 17688 23354 17700
rect 22005 17663 22063 17669
rect 22005 17660 22017 17663
rect 21652 17632 22017 17660
rect 22005 17629 22017 17632
rect 22051 17629 22063 17663
rect 22465 17663 22523 17669
rect 22465 17660 22477 17663
rect 22005 17623 22063 17629
rect 22204 17632 22477 17660
rect 12710 17552 12716 17604
rect 12768 17552 12774 17604
rect 15378 17601 15384 17604
rect 15372 17555 15384 17601
rect 15378 17552 15384 17555
rect 15436 17552 15442 17604
rect 17712 17595 17770 17601
rect 17712 17561 17724 17595
rect 17758 17592 17770 17595
rect 17758 17564 18092 17592
rect 17758 17561 17770 17564
rect 17712 17555 17770 17561
rect 10870 17484 10876 17536
rect 10928 17484 10934 17536
rect 10965 17527 11023 17533
rect 10965 17493 10977 17527
rect 11011 17524 11023 17527
rect 11790 17524 11796 17536
rect 11011 17496 11796 17524
rect 11011 17493 11023 17496
rect 10965 17487 11023 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 16485 17527 16543 17533
rect 16485 17524 16497 17527
rect 15620 17496 16497 17524
rect 15620 17484 15626 17496
rect 16485 17493 16497 17496
rect 16531 17493 16543 17527
rect 16485 17487 16543 17493
rect 16574 17484 16580 17536
rect 16632 17484 16638 17536
rect 18064 17533 18092 17564
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19518 17592 19524 17604
rect 19392 17564 19524 17592
rect 19392 17552 19398 17564
rect 19518 17552 19524 17564
rect 19576 17592 19582 17604
rect 20622 17592 20628 17604
rect 19576 17564 20628 17592
rect 19576 17552 19582 17564
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 22204 17536 22232 17632
rect 22465 17629 22477 17632
rect 22511 17629 22523 17663
rect 22465 17623 22523 17629
rect 22833 17663 22891 17669
rect 22833 17629 22845 17663
rect 22879 17660 22891 17663
rect 23400 17660 23428 17700
rect 23569 17697 23581 17731
rect 23615 17728 23627 17731
rect 23934 17728 23940 17740
rect 23615 17700 23940 17728
rect 23615 17697 23627 17700
rect 23569 17691 23627 17697
rect 23934 17688 23940 17700
rect 23992 17688 23998 17740
rect 25148 17672 25176 17836
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 22879 17632 23336 17660
rect 23400 17632 23673 17660
rect 22879 17629 22891 17632
rect 22833 17623 22891 17629
rect 22370 17552 22376 17604
rect 22428 17592 22434 17604
rect 22557 17595 22615 17601
rect 22557 17592 22569 17595
rect 22428 17564 22569 17592
rect 22428 17552 22434 17564
rect 22557 17561 22569 17564
rect 22603 17561 22615 17595
rect 22557 17555 22615 17561
rect 22649 17595 22707 17601
rect 22649 17561 22661 17595
rect 22695 17592 22707 17595
rect 23198 17592 23204 17604
rect 22695 17564 23204 17592
rect 22695 17561 22707 17564
rect 22649 17555 22707 17561
rect 23198 17552 23204 17564
rect 23256 17552 23262 17604
rect 23308 17592 23336 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 23750 17620 23756 17672
rect 23808 17620 23814 17672
rect 24397 17663 24455 17669
rect 24397 17629 24409 17663
rect 24443 17629 24455 17663
rect 24397 17623 24455 17629
rect 23768 17592 23796 17620
rect 23308 17564 23796 17592
rect 23842 17552 23848 17604
rect 23900 17592 23906 17604
rect 23937 17595 23995 17601
rect 23937 17592 23949 17595
rect 23900 17564 23949 17592
rect 23900 17552 23906 17564
rect 23937 17561 23949 17564
rect 23983 17592 23995 17595
rect 24412 17592 24440 17623
rect 25130 17620 25136 17672
rect 25188 17620 25194 17672
rect 25406 17669 25412 17672
rect 25400 17623 25412 17669
rect 25464 17660 25470 17672
rect 26160 17660 26188 17836
rect 26513 17833 26525 17867
rect 26559 17864 26571 17867
rect 27614 17864 27620 17876
rect 26559 17836 27620 17864
rect 26559 17833 26571 17836
rect 26513 17827 26571 17833
rect 27614 17824 27620 17836
rect 27672 17824 27678 17876
rect 30837 17867 30895 17873
rect 30837 17833 30849 17867
rect 30883 17864 30895 17867
rect 31202 17864 31208 17876
rect 30883 17836 31208 17864
rect 30883 17833 30895 17836
rect 30837 17827 30895 17833
rect 31202 17824 31208 17836
rect 31260 17824 31266 17876
rect 33689 17867 33747 17873
rect 33689 17864 33701 17867
rect 31404 17836 33701 17864
rect 30282 17688 30288 17740
rect 30340 17728 30346 17740
rect 30377 17731 30435 17737
rect 30377 17728 30389 17731
rect 30340 17700 30389 17728
rect 30340 17688 30346 17700
rect 30377 17697 30389 17700
rect 30423 17697 30435 17731
rect 30377 17691 30435 17697
rect 30561 17731 30619 17737
rect 30561 17697 30573 17731
rect 30607 17728 30619 17731
rect 30650 17728 30656 17740
rect 30607 17700 30656 17728
rect 30607 17697 30619 17700
rect 30561 17691 30619 17697
rect 30650 17688 30656 17700
rect 30708 17688 30714 17740
rect 27982 17660 27988 17672
rect 25464 17632 25500 17660
rect 26160 17632 27988 17660
rect 25406 17620 25412 17623
rect 25464 17620 25470 17632
rect 27982 17620 27988 17632
rect 28040 17620 28046 17672
rect 28258 17620 28264 17672
rect 28316 17620 28322 17672
rect 30742 17620 30748 17672
rect 30800 17620 30806 17672
rect 30834 17620 30840 17672
rect 30892 17620 30898 17672
rect 31018 17620 31024 17672
rect 31076 17660 31082 17672
rect 31404 17669 31432 17836
rect 33689 17833 33701 17836
rect 33735 17833 33747 17867
rect 35342 17864 35348 17876
rect 33689 17827 33747 17833
rect 33888 17836 35348 17864
rect 32861 17799 32919 17805
rect 32861 17765 32873 17799
rect 32907 17765 32919 17799
rect 32861 17759 32919 17765
rect 32876 17728 32904 17759
rect 32953 17731 33011 17737
rect 32953 17728 32965 17731
rect 32876 17700 32965 17728
rect 32953 17697 32965 17700
rect 32999 17697 33011 17731
rect 32953 17691 33011 17697
rect 31205 17663 31263 17669
rect 31205 17660 31217 17663
rect 31076 17632 31217 17660
rect 31076 17620 31082 17632
rect 31205 17629 31217 17632
rect 31251 17629 31263 17663
rect 31205 17623 31263 17629
rect 31389 17663 31447 17669
rect 31389 17629 31401 17663
rect 31435 17629 31447 17663
rect 31389 17623 31447 17629
rect 31478 17620 31484 17672
rect 31536 17620 31542 17672
rect 33888 17669 33916 17836
rect 35342 17824 35348 17836
rect 35400 17864 35406 17876
rect 35894 17864 35900 17876
rect 35400 17836 35900 17864
rect 35400 17824 35406 17836
rect 33962 17756 33968 17808
rect 34020 17756 34026 17808
rect 33980 17669 34008 17756
rect 33873 17663 33931 17669
rect 33873 17629 33885 17663
rect 33919 17629 33931 17663
rect 33873 17623 33931 17629
rect 33965 17663 34023 17669
rect 33965 17629 33977 17663
rect 34011 17629 34023 17663
rect 33965 17623 34023 17629
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 34701 17663 34759 17669
rect 34701 17660 34713 17663
rect 34572 17632 34713 17660
rect 34572 17620 34578 17632
rect 34701 17629 34713 17632
rect 34747 17629 34759 17663
rect 34701 17623 34759 17629
rect 23983 17564 24440 17592
rect 27740 17595 27798 17601
rect 23983 17561 23995 17564
rect 23937 17555 23995 17561
rect 27740 17561 27752 17595
rect 27786 17592 27798 17595
rect 31297 17595 31355 17601
rect 27786 17564 28120 17592
rect 27786 17561 27798 17564
rect 27740 17555 27798 17561
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17493 18107 17527
rect 18049 17487 18107 17493
rect 19426 17484 19432 17536
rect 19484 17484 19490 17536
rect 21082 17484 21088 17536
rect 21140 17484 21146 17536
rect 21177 17527 21235 17533
rect 21177 17493 21189 17527
rect 21223 17524 21235 17527
rect 22094 17524 22100 17536
rect 21223 17496 22100 17524
rect 21223 17493 21235 17496
rect 21177 17487 21235 17493
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 22186 17484 22192 17536
rect 22244 17484 22250 17536
rect 22278 17484 22284 17536
rect 22336 17484 22342 17536
rect 26510 17484 26516 17536
rect 26568 17524 26574 17536
rect 28092 17533 28120 17564
rect 31297 17561 31309 17595
rect 31343 17592 31355 17595
rect 31726 17595 31784 17601
rect 31726 17592 31738 17595
rect 31343 17564 31738 17592
rect 31343 17561 31355 17564
rect 31297 17555 31355 17561
rect 31726 17561 31738 17564
rect 31772 17561 31784 17595
rect 31726 17555 31784 17561
rect 33689 17595 33747 17601
rect 33689 17561 33701 17595
rect 33735 17561 33747 17595
rect 34946 17595 35004 17601
rect 34946 17592 34958 17595
rect 33689 17555 33747 17561
rect 34716 17564 34958 17592
rect 26605 17527 26663 17533
rect 26605 17524 26617 17527
rect 26568 17496 26617 17524
rect 26568 17484 26574 17496
rect 26605 17493 26617 17496
rect 26651 17493 26663 17527
rect 26605 17487 26663 17493
rect 28077 17527 28135 17533
rect 28077 17493 28089 17527
rect 28123 17493 28135 17527
rect 28077 17487 28135 17493
rect 29822 17484 29828 17536
rect 29880 17484 29886 17536
rect 33597 17527 33655 17533
rect 33597 17493 33609 17527
rect 33643 17524 33655 17527
rect 33704 17524 33732 17555
rect 34716 17536 34744 17564
rect 34946 17561 34958 17564
rect 34992 17561 35004 17595
rect 35728 17592 35756 17836
rect 35894 17824 35900 17836
rect 35952 17824 35958 17876
rect 38105 17867 38163 17873
rect 38105 17833 38117 17867
rect 38151 17833 38163 17867
rect 38105 17827 38163 17833
rect 36078 17756 36084 17808
rect 36136 17756 36142 17808
rect 36096 17728 36124 17756
rect 38120 17728 38148 17827
rect 38286 17824 38292 17876
rect 38344 17824 38350 17876
rect 36096 17700 38148 17728
rect 36832 17672 36860 17700
rect 36265 17663 36323 17669
rect 36265 17629 36277 17663
rect 36311 17660 36323 17663
rect 36446 17660 36452 17672
rect 36311 17632 36452 17660
rect 36311 17629 36323 17632
rect 36265 17623 36323 17629
rect 36446 17620 36452 17632
rect 36504 17620 36510 17672
rect 36814 17620 36820 17672
rect 36872 17620 36878 17672
rect 36906 17620 36912 17672
rect 36964 17620 36970 17672
rect 37093 17663 37151 17669
rect 37093 17629 37105 17663
rect 37139 17629 37151 17663
rect 37093 17623 37151 17629
rect 36541 17595 36599 17601
rect 36541 17592 36553 17595
rect 35728 17564 36553 17592
rect 34946 17555 35004 17561
rect 36541 17561 36553 17564
rect 36587 17592 36599 17595
rect 36722 17592 36728 17604
rect 36587 17564 36728 17592
rect 36587 17561 36599 17564
rect 36541 17555 36599 17561
rect 36722 17552 36728 17564
rect 36780 17552 36786 17604
rect 33778 17524 33784 17536
rect 33643 17496 33784 17524
rect 33643 17493 33655 17496
rect 33597 17487 33655 17493
rect 33778 17484 33784 17496
rect 33836 17484 33842 17536
rect 34698 17484 34704 17536
rect 34756 17484 34762 17536
rect 36924 17524 36952 17620
rect 37108 17592 37136 17623
rect 37182 17620 37188 17672
rect 37240 17620 37246 17672
rect 37826 17620 37832 17672
rect 37884 17620 37890 17672
rect 37918 17592 37924 17604
rect 37108 17564 37924 17592
rect 37918 17552 37924 17564
rect 37976 17552 37982 17604
rect 38121 17527 38179 17533
rect 38121 17524 38133 17527
rect 36924 17496 38133 17524
rect 38121 17493 38133 17496
rect 38167 17493 38179 17527
rect 38121 17487 38179 17493
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 4120 17292 12434 17320
rect 4120 17280 4126 17292
rect 7742 17252 7748 17264
rect 7484 17224 7748 17252
rect 7484 17193 7512 17224
rect 7742 17212 7748 17224
rect 7800 17212 7806 17264
rect 8478 17212 8484 17264
rect 8536 17212 8542 17264
rect 9122 17212 9128 17264
rect 9180 17212 9186 17264
rect 9861 17255 9919 17261
rect 9861 17221 9873 17255
rect 9907 17252 9919 17255
rect 9950 17252 9956 17264
rect 9907 17224 9956 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 9950 17212 9956 17224
rect 10008 17212 10014 17264
rect 10870 17212 10876 17264
rect 10928 17212 10934 17264
rect 12406 17252 12434 17292
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 13173 17323 13231 17329
rect 13173 17320 13185 17323
rect 12768 17292 13185 17320
rect 12768 17280 12774 17292
rect 13173 17289 13185 17292
rect 13219 17289 13231 17323
rect 13173 17283 13231 17289
rect 15289 17323 15347 17329
rect 15289 17289 15301 17323
rect 15335 17320 15347 17323
rect 15378 17320 15384 17332
rect 15335 17292 15384 17320
rect 15335 17289 15347 17292
rect 15289 17283 15347 17289
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15650 17323 15708 17329
rect 15650 17289 15662 17323
rect 15696 17320 15708 17323
rect 17218 17320 17224 17332
rect 15696 17292 17224 17320
rect 15696 17289 15708 17292
rect 15650 17283 15708 17289
rect 17218 17280 17224 17292
rect 17276 17280 17282 17332
rect 18966 17280 18972 17332
rect 19024 17280 19030 17332
rect 19058 17280 19064 17332
rect 19116 17280 19122 17332
rect 24581 17323 24639 17329
rect 19245 17289 19303 17295
rect 18874 17252 18880 17264
rect 12406 17224 18880 17252
rect 18874 17212 18880 17224
rect 18932 17212 18938 17264
rect 19150 17212 19156 17264
rect 19208 17252 19214 17264
rect 19245 17255 19257 17289
rect 19291 17255 19303 17289
rect 24581 17289 24593 17323
rect 24627 17320 24639 17323
rect 24670 17320 24676 17332
rect 24627 17292 24676 17320
rect 24627 17289 24639 17292
rect 24581 17283 24639 17289
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 25498 17280 25504 17332
rect 25556 17320 25562 17332
rect 25777 17323 25835 17329
rect 25777 17320 25789 17323
rect 25556 17292 25789 17320
rect 25556 17280 25562 17292
rect 25777 17289 25789 17292
rect 25823 17289 25835 17323
rect 26326 17320 26332 17332
rect 25777 17283 25835 17289
rect 25884 17292 26332 17320
rect 19245 17252 19303 17255
rect 19208 17249 19303 17252
rect 19208 17224 19288 17249
rect 19423 17224 23060 17252
rect 19208 17212 19214 17224
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 7745 17119 7803 17125
rect 7745 17085 7757 17119
rect 7791 17116 7803 17119
rect 8754 17116 8760 17128
rect 7791 17088 8760 17116
rect 7791 17085 7803 17088
rect 7745 17079 7803 17085
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 9140 17048 9168 17212
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9732 17156 9781 17184
rect 9732 17144 9738 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 10888 17184 10916 17212
rect 19423 17206 19451 17224
rect 12345 17187 12403 17193
rect 12345 17184 12357 17187
rect 10888 17156 12357 17184
rect 9769 17147 9827 17153
rect 12345 17153 12357 17156
rect 12391 17153 12403 17187
rect 12345 17147 12403 17153
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17184 13323 17187
rect 13814 17184 13820 17196
rect 13311 17156 13820 17184
rect 13311 17153 13323 17156
rect 13265 17147 13323 17153
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14849 17187 14907 17193
rect 14849 17153 14861 17187
rect 14895 17184 14907 17187
rect 15010 17184 15016 17196
rect 14895 17156 15016 17184
rect 14895 17153 14907 17156
rect 14849 17147 14907 17153
rect 15010 17144 15016 17156
rect 15068 17144 15074 17196
rect 15102 17144 15108 17196
rect 15160 17144 15166 17196
rect 15194 17144 15200 17196
rect 15252 17144 15258 17196
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9916 17088 9965 17116
rect 9916 17076 9922 17088
rect 9953 17085 9965 17088
rect 9999 17116 10011 17119
rect 10686 17116 10692 17128
rect 9999 17088 10692 17116
rect 9999 17085 10011 17088
rect 9953 17079 10011 17085
rect 10686 17076 10692 17088
rect 10744 17076 10750 17128
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17085 10839 17119
rect 10781 17079 10839 17085
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17085 13047 17119
rect 12989 17079 13047 17085
rect 9401 17051 9459 17057
rect 9401 17048 9413 17051
rect 9140 17020 9413 17048
rect 9401 17017 9413 17020
rect 9447 17017 9459 17051
rect 10796 17048 10824 17079
rect 9401 17011 9459 17017
rect 10060 17020 10824 17048
rect 13004 17048 13032 17079
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 13004 17020 13737 17048
rect 9217 16983 9275 16989
rect 9217 16949 9229 16983
rect 9263 16980 9275 16983
rect 9306 16980 9312 16992
rect 9263 16952 9312 16980
rect 9263 16949 9275 16952
rect 9217 16943 9275 16949
rect 9306 16940 9312 16952
rect 9364 16980 9370 16992
rect 10060 16980 10088 17020
rect 13725 17017 13737 17020
rect 13771 17017 13783 17051
rect 13725 17011 13783 17017
rect 9364 16952 10088 16980
rect 9364 16940 9370 16952
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 10192 16952 10241 16980
rect 10192 16940 10198 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10229 16943 10287 16949
rect 14918 16940 14924 16992
rect 14976 16980 14982 16992
rect 15212 16980 15240 17144
rect 15396 17048 15424 17147
rect 15470 17144 15476 17196
rect 15528 17144 15534 17196
rect 15562 17144 15568 17196
rect 15620 17144 15626 17196
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17184 15807 17187
rect 15795 17156 16528 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 15654 17076 15660 17128
rect 15712 17116 15718 17128
rect 16022 17116 16028 17128
rect 15712 17088 16028 17116
rect 15712 17076 15718 17088
rect 16022 17076 16028 17088
rect 16080 17116 16086 17128
rect 16393 17119 16451 17125
rect 16393 17116 16405 17119
rect 16080 17088 16405 17116
rect 16080 17076 16086 17088
rect 16393 17085 16405 17088
rect 16439 17085 16451 17119
rect 16500 17116 16528 17156
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 16632 17156 17233 17184
rect 16632 17144 16638 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17856 17187 17914 17193
rect 17856 17153 17868 17187
rect 17902 17184 17914 17187
rect 18138 17184 18144 17196
rect 17902 17156 18144 17184
rect 17902 17153 17914 17156
rect 17856 17147 17914 17153
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 18966 17144 18972 17196
rect 19024 17144 19030 17196
rect 19242 17187 19300 17193
rect 19242 17153 19254 17187
rect 19288 17182 19300 17187
rect 19352 17182 19451 17206
rect 20533 17187 20591 17193
rect 20533 17184 20545 17187
rect 19288 17178 19451 17182
rect 19288 17154 19380 17178
rect 19516 17156 20545 17184
rect 19288 17153 19300 17154
rect 19242 17147 19300 17153
rect 16669 17119 16727 17125
rect 16669 17116 16681 17119
rect 16500 17088 16681 17116
rect 16393 17079 16451 17085
rect 16669 17085 16681 17088
rect 16715 17085 16727 17119
rect 16669 17079 16727 17085
rect 16758 17076 16764 17128
rect 16816 17076 16822 17128
rect 17586 17076 17592 17128
rect 17644 17076 17650 17128
rect 16776 17048 16804 17076
rect 15396 17020 16804 17048
rect 14976 16952 15240 16980
rect 14976 16940 14982 16952
rect 15838 16940 15844 16992
rect 15896 16940 15902 16992
rect 16390 16940 16396 16992
rect 16448 16980 16454 16992
rect 18984 16980 19012 17144
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 19516 17116 19544 17156
rect 20533 17153 20545 17156
rect 20579 17153 20591 17187
rect 20533 17147 20591 17153
rect 21634 17144 21640 17196
rect 21692 17184 21698 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 21692 17156 21833 17184
rect 21692 17144 21698 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22278 17144 22284 17196
rect 22336 17184 22342 17196
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 22336 17156 22385 17184
rect 22336 17144 22342 17156
rect 22373 17153 22385 17156
rect 22419 17153 22431 17187
rect 23032 17184 23060 17224
rect 23106 17212 23112 17264
rect 23164 17212 23170 17264
rect 25593 17255 25651 17261
rect 25593 17221 25605 17255
rect 25639 17252 25651 17255
rect 25884 17252 25912 17292
rect 26326 17280 26332 17292
rect 26384 17280 26390 17332
rect 26694 17320 26700 17332
rect 26436 17292 26700 17320
rect 25639 17224 25912 17252
rect 25639 17221 25651 17224
rect 25593 17215 25651 17221
rect 25958 17212 25964 17264
rect 26016 17252 26022 17264
rect 26436 17252 26464 17292
rect 26694 17280 26700 17292
rect 26752 17280 26758 17332
rect 26789 17323 26847 17329
rect 26789 17289 26801 17323
rect 26835 17320 26847 17323
rect 28258 17320 28264 17332
rect 26835 17292 28264 17320
rect 26835 17289 26847 17292
rect 26789 17283 26847 17289
rect 28258 17280 28264 17292
rect 28316 17280 28322 17332
rect 29730 17280 29736 17332
rect 29788 17280 29794 17332
rect 29822 17280 29828 17332
rect 29880 17280 29886 17332
rect 32401 17323 32459 17329
rect 32401 17320 32413 17323
rect 31726 17292 32413 17320
rect 29840 17252 29868 17280
rect 29917 17255 29975 17261
rect 29917 17252 29929 17255
rect 26016 17224 26464 17252
rect 26528 17224 29776 17252
rect 29840 17224 29929 17252
rect 26016 17212 26022 17224
rect 26528 17184 26556 17224
rect 23032 17156 25544 17184
rect 22373 17147 22431 17153
rect 19116 17108 19196 17116
rect 19306 17108 19544 17116
rect 19116 17088 19544 17108
rect 19705 17119 19763 17125
rect 19116 17076 19122 17088
rect 19168 17080 19334 17088
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 20438 17116 20444 17128
rect 19751 17088 20444 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 20438 17076 20444 17088
rect 20496 17076 20502 17128
rect 21266 17076 21272 17128
rect 21324 17076 21330 17128
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17116 22155 17119
rect 23198 17116 23204 17128
rect 22143 17088 23204 17116
rect 22143 17085 22155 17088
rect 22097 17079 22155 17085
rect 23198 17076 23204 17088
rect 23256 17076 23262 17128
rect 25516 17116 25544 17156
rect 26344 17156 26556 17184
rect 26344 17116 26372 17156
rect 26602 17144 26608 17196
rect 26660 17144 26666 17196
rect 26694 17144 26700 17196
rect 26752 17184 26758 17196
rect 26973 17187 27031 17193
rect 26973 17184 26985 17187
rect 26752 17156 26985 17184
rect 26752 17144 26758 17156
rect 26973 17153 26985 17156
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 29638 17144 29644 17196
rect 29696 17144 29702 17196
rect 29748 17184 29776 17224
rect 29917 17221 29929 17224
rect 29963 17221 29975 17255
rect 29917 17215 29975 17221
rect 31726 17184 31754 17292
rect 32401 17289 32413 17292
rect 32447 17320 32459 17323
rect 34606 17320 34612 17332
rect 32447 17292 34612 17320
rect 32447 17289 32459 17292
rect 32401 17283 32459 17289
rect 34606 17280 34612 17292
rect 34664 17280 34670 17332
rect 34698 17280 34704 17332
rect 34756 17280 34762 17332
rect 34790 17280 34796 17332
rect 34848 17280 34854 17332
rect 35897 17323 35955 17329
rect 35897 17289 35909 17323
rect 35943 17320 35955 17323
rect 36814 17320 36820 17332
rect 35943 17292 36820 17320
rect 35943 17289 35955 17292
rect 35897 17283 35955 17289
rect 36814 17280 36820 17292
rect 36872 17280 36878 17332
rect 37826 17280 37832 17332
rect 37884 17320 37890 17332
rect 37884 17292 38240 17320
rect 37884 17280 37890 17292
rect 32217 17255 32275 17261
rect 32217 17221 32229 17255
rect 32263 17252 32275 17255
rect 32263 17224 32706 17252
rect 32263 17221 32275 17224
rect 32217 17215 32275 17221
rect 33778 17212 33784 17264
rect 33836 17252 33842 17264
rect 33873 17255 33931 17261
rect 33873 17252 33885 17255
rect 33836 17224 33885 17252
rect 33836 17212 33842 17224
rect 33873 17221 33885 17224
rect 33919 17221 33931 17255
rect 33873 17215 33931 17221
rect 33962 17212 33968 17264
rect 34020 17252 34026 17264
rect 34020 17224 34744 17252
rect 34020 17212 34026 17224
rect 29748 17156 31754 17184
rect 31846 17144 31852 17196
rect 31904 17184 31910 17196
rect 32125 17187 32183 17193
rect 32125 17184 32137 17187
rect 31904 17156 32137 17184
rect 31904 17144 31910 17156
rect 32125 17153 32137 17156
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 25516 17088 26372 17116
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17116 26479 17119
rect 27706 17116 27712 17128
rect 26467 17088 27712 17116
rect 26467 17085 26479 17088
rect 26421 17079 26479 17085
rect 27706 17076 27712 17088
rect 27764 17076 27770 17128
rect 27890 17076 27896 17128
rect 27948 17076 27954 17128
rect 30742 17076 30748 17128
rect 30800 17076 30806 17128
rect 34149 17119 34207 17125
rect 34149 17085 34161 17119
rect 34195 17116 34207 17119
rect 34514 17116 34520 17128
rect 34195 17088 34520 17116
rect 34195 17085 34207 17088
rect 34149 17079 34207 17085
rect 19518 17008 19524 17060
rect 19576 17048 19582 17060
rect 19981 17051 20039 17057
rect 19981 17048 19993 17051
rect 19576 17020 19993 17048
rect 19576 17008 19582 17020
rect 19981 17017 19993 17020
rect 20027 17017 20039 17051
rect 19981 17011 20039 17017
rect 21913 17051 21971 17057
rect 21913 17017 21925 17051
rect 21959 17048 21971 17051
rect 22646 17048 22652 17060
rect 21959 17020 22652 17048
rect 21959 17017 21971 17020
rect 21913 17011 21971 17017
rect 22646 17008 22652 17020
rect 22704 17008 22710 17060
rect 25222 17008 25228 17060
rect 25280 17048 25286 17060
rect 25682 17048 25688 17060
rect 25280 17020 25688 17048
rect 25280 17008 25286 17020
rect 25682 17008 25688 17020
rect 25740 17008 25746 17060
rect 29917 17051 29975 17057
rect 29917 17017 29929 17051
rect 29963 17048 29975 17051
rect 30760 17048 30788 17076
rect 29963 17020 30788 17048
rect 29963 17017 29975 17020
rect 29917 17011 29975 17017
rect 16448 16952 19012 16980
rect 16448 16940 16454 16952
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19613 16983 19671 16989
rect 19613 16980 19625 16983
rect 19484 16952 19625 16980
rect 19484 16940 19490 16952
rect 19613 16949 19625 16952
rect 19659 16949 19671 16983
rect 19613 16943 19671 16949
rect 20717 16983 20775 16989
rect 20717 16949 20729 16983
rect 20763 16980 20775 16983
rect 20806 16980 20812 16992
rect 20763 16952 20812 16980
rect 20763 16949 20775 16952
rect 20717 16943 20775 16949
rect 20806 16940 20812 16952
rect 20864 16940 20870 16992
rect 22005 16983 22063 16989
rect 22005 16949 22017 16983
rect 22051 16980 22063 16983
rect 22370 16980 22376 16992
rect 22051 16952 22376 16980
rect 22051 16949 22063 16952
rect 22005 16943 22063 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 23017 16983 23075 16989
rect 23017 16949 23029 16983
rect 23063 16980 23075 16983
rect 23106 16980 23112 16992
rect 23063 16952 23112 16980
rect 23063 16949 23075 16952
rect 23017 16943 23075 16949
rect 23106 16940 23112 16952
rect 23164 16940 23170 16992
rect 25593 16983 25651 16989
rect 25593 16949 25605 16983
rect 25639 16980 25651 16983
rect 25866 16980 25872 16992
rect 25639 16952 25872 16980
rect 25639 16949 25651 16952
rect 25593 16943 25651 16949
rect 25866 16940 25872 16952
rect 25924 16940 25930 16992
rect 27614 16940 27620 16992
rect 27672 16940 27678 16992
rect 28258 16940 28264 16992
rect 28316 16980 28322 16992
rect 28537 16983 28595 16989
rect 28537 16980 28549 16983
rect 28316 16952 28549 16980
rect 28316 16940 28322 16952
rect 28537 16949 28549 16952
rect 28583 16949 28595 16983
rect 28537 16943 28595 16949
rect 33410 16940 33416 16992
rect 33468 16980 33474 16992
rect 34164 16980 34192 17079
rect 34514 17076 34520 17088
rect 34572 17076 34578 17128
rect 34716 17116 34744 17224
rect 34808 17184 34836 17280
rect 35176 17224 35848 17252
rect 35176 17193 35204 17224
rect 35820 17193 35848 17224
rect 37090 17212 37096 17264
rect 37148 17252 37154 17264
rect 38013 17255 38071 17261
rect 38013 17252 38025 17255
rect 37148 17224 38025 17252
rect 37148 17212 37154 17224
rect 38013 17221 38025 17224
rect 38059 17221 38071 17255
rect 38013 17215 38071 17221
rect 38212 17193 38240 17292
rect 38286 17280 38292 17332
rect 38344 17280 38350 17332
rect 38304 17193 38332 17280
rect 34885 17187 34943 17193
rect 34885 17184 34897 17187
rect 34808 17156 34897 17184
rect 34885 17153 34897 17156
rect 34931 17153 34943 17187
rect 34885 17147 34943 17153
rect 35161 17187 35219 17193
rect 35161 17153 35173 17187
rect 35207 17153 35219 17187
rect 35161 17147 35219 17153
rect 35345 17187 35403 17193
rect 35345 17153 35357 17187
rect 35391 17153 35403 17187
rect 35345 17147 35403 17153
rect 35805 17187 35863 17193
rect 35805 17153 35817 17187
rect 35851 17153 35863 17187
rect 35805 17147 35863 17153
rect 36081 17187 36139 17193
rect 36081 17153 36093 17187
rect 36127 17184 36139 17187
rect 37277 17187 37335 17193
rect 37277 17184 37289 17187
rect 36127 17156 37289 17184
rect 36127 17153 36139 17156
rect 36081 17147 36139 17153
rect 37277 17153 37289 17156
rect 37323 17153 37335 17187
rect 37277 17147 37335 17153
rect 38197 17187 38255 17193
rect 38197 17153 38209 17187
rect 38243 17153 38255 17187
rect 38197 17147 38255 17153
rect 38289 17187 38347 17193
rect 38289 17153 38301 17187
rect 38335 17153 38347 17187
rect 38289 17147 38347 17153
rect 35176 17116 35204 17147
rect 34716 17088 35204 17116
rect 35360 17116 35388 17147
rect 36173 17119 36231 17125
rect 36173 17116 36185 17119
rect 35360 17088 36185 17116
rect 36173 17085 36185 17088
rect 36219 17085 36231 17119
rect 36173 17079 36231 17085
rect 36814 17076 36820 17128
rect 36872 17076 36878 17128
rect 37182 17076 37188 17128
rect 37240 17076 37246 17128
rect 37918 17076 37924 17128
rect 37976 17076 37982 17128
rect 36081 17051 36139 17057
rect 36081 17017 36093 17051
rect 36127 17048 36139 17051
rect 37200 17048 37228 17076
rect 36127 17020 37228 17048
rect 36127 17017 36139 17020
rect 36081 17011 36139 17017
rect 33468 16952 34192 16980
rect 33468 16940 33474 16952
rect 38102 16940 38108 16992
rect 38160 16940 38166 16992
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 8573 16779 8631 16785
rect 8573 16776 8585 16779
rect 8536 16748 8585 16776
rect 8536 16736 8542 16748
rect 8573 16745 8585 16748
rect 8619 16745 8631 16779
rect 8573 16739 8631 16745
rect 8754 16736 8760 16788
rect 8812 16776 8818 16788
rect 9585 16779 9643 16785
rect 9585 16776 9597 16779
rect 8812 16748 9597 16776
rect 8812 16736 8818 16748
rect 9585 16745 9597 16748
rect 9631 16745 9643 16779
rect 9585 16739 9643 16745
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 13780 16748 13952 16776
rect 13780 16736 13786 16748
rect 9493 16711 9551 16717
rect 9493 16677 9505 16711
rect 9539 16708 9551 16711
rect 9539 16680 9904 16708
rect 9539 16677 9551 16680
rect 9493 16671 9551 16677
rect 8662 16640 8668 16652
rect 8496 16612 8668 16640
rect 8496 16581 8524 16612
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16572 9275 16575
rect 9769 16575 9827 16581
rect 9263 16544 9444 16572
rect 9263 16541 9275 16544
rect 9217 16535 9275 16541
rect 9306 16396 9312 16448
rect 9364 16396 9370 16448
rect 9416 16436 9444 16544
rect 9769 16541 9781 16575
rect 9815 16572 9827 16575
rect 9876 16572 9904 16680
rect 10042 16668 10048 16720
rect 10100 16708 10106 16720
rect 11422 16708 11428 16720
rect 10100 16680 11428 16708
rect 10100 16668 10106 16680
rect 11422 16668 11428 16680
rect 11480 16708 11486 16720
rect 11480 16680 11744 16708
rect 11480 16668 11486 16680
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 11514 16640 11520 16652
rect 11287 16612 11520 16640
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 11716 16640 11744 16680
rect 12618 16640 12624 16652
rect 11716 16612 12624 16640
rect 9815 16544 10088 16572
rect 9815 16541 9827 16544
rect 9769 16535 9827 16541
rect 9490 16464 9496 16516
rect 9548 16464 9554 16516
rect 9858 16464 9864 16516
rect 9916 16464 9922 16516
rect 9950 16464 9956 16516
rect 10008 16464 10014 16516
rect 10060 16504 10088 16544
rect 10134 16532 10140 16584
rect 10192 16532 10198 16584
rect 11716 16581 11744 16612
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 13924 16649 13952 16748
rect 15010 16736 15016 16788
rect 15068 16776 15074 16788
rect 15197 16779 15255 16785
rect 15197 16776 15209 16779
rect 15068 16748 15209 16776
rect 15068 16736 15074 16748
rect 15197 16745 15209 16748
rect 15243 16745 15255 16779
rect 15197 16739 15255 16745
rect 17957 16779 18015 16785
rect 17957 16745 17969 16779
rect 18003 16776 18015 16779
rect 18138 16776 18144 16788
rect 18003 16748 18144 16776
rect 18003 16745 18015 16748
rect 17957 16739 18015 16745
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 18966 16736 18972 16788
rect 19024 16736 19030 16788
rect 19978 16776 19984 16788
rect 19812 16748 19984 16776
rect 16390 16708 16396 16720
rect 14936 16680 16396 16708
rect 13909 16643 13967 16649
rect 13909 16609 13921 16643
rect 13955 16609 13967 16643
rect 13909 16603 13967 16609
rect 11882 16581 11888 16584
rect 11425 16575 11483 16581
rect 11425 16541 11437 16575
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 11701 16575 11759 16581
rect 11701 16541 11713 16575
rect 11747 16541 11759 16575
rect 11878 16572 11888 16581
rect 11843 16544 11888 16572
rect 11701 16535 11759 16541
rect 11878 16535 11888 16544
rect 10229 16507 10287 16513
rect 10229 16504 10241 16507
rect 10060 16476 10241 16504
rect 10229 16473 10241 16476
rect 10275 16473 10287 16507
rect 10229 16467 10287 16473
rect 10410 16464 10416 16516
rect 10468 16504 10474 16516
rect 10468 16476 11008 16504
rect 10468 16464 10474 16476
rect 9876 16436 9904 16464
rect 9416 16408 9904 16436
rect 9968 16436 9996 16464
rect 10597 16439 10655 16445
rect 10597 16436 10609 16439
rect 9968 16408 10609 16436
rect 10597 16405 10609 16408
rect 10643 16405 10655 16439
rect 10980 16436 11008 16476
rect 11054 16464 11060 16516
rect 11112 16504 11118 16516
rect 11440 16504 11468 16535
rect 11882 16532 11888 16535
rect 11940 16532 11946 16584
rect 12250 16532 12256 16584
rect 12308 16532 12314 16584
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13096 16544 14105 16572
rect 11793 16507 11851 16513
rect 11793 16504 11805 16507
rect 11112 16476 11805 16504
rect 11112 16464 11118 16476
rect 11793 16473 11805 16476
rect 11839 16473 11851 16507
rect 11793 16467 11851 16473
rect 13096 16448 13124 16544
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14734 16532 14740 16584
rect 14792 16532 14798 16584
rect 14936 16581 14964 16680
rect 16390 16668 16396 16680
rect 16448 16668 16454 16720
rect 18984 16708 19012 16736
rect 16859 16680 19012 16708
rect 19337 16711 19395 16717
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 16577 16643 16635 16649
rect 16577 16640 16589 16643
rect 15620 16612 16589 16640
rect 15620 16600 15626 16612
rect 16577 16609 16589 16612
rect 16623 16640 16635 16643
rect 16761 16643 16819 16649
rect 16761 16640 16773 16643
rect 16623 16612 16773 16640
rect 16623 16609 16635 16612
rect 16577 16603 16635 16609
rect 16761 16609 16773 16612
rect 16807 16609 16819 16643
rect 16761 16603 16819 16609
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 15197 16575 15255 16581
rect 15197 16541 15209 16575
rect 15243 16572 15255 16575
rect 15289 16575 15347 16581
rect 15289 16572 15301 16575
rect 15243 16544 15301 16572
rect 15243 16541 15255 16544
rect 15197 16535 15255 16541
rect 15289 16541 15301 16544
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 15930 16532 15936 16584
rect 15988 16532 15994 16584
rect 13664 16507 13722 16513
rect 13664 16473 13676 16507
rect 13710 16504 13722 16507
rect 15028 16504 15056 16532
rect 16859 16504 16887 16680
rect 17865 16643 17923 16649
rect 17865 16609 17877 16643
rect 17911 16640 17923 16643
rect 17911 16612 18184 16640
rect 17911 16609 17923 16612
rect 17865 16603 17923 16609
rect 18156 16581 18184 16612
rect 18892 16581 18920 16680
rect 19337 16677 19349 16711
rect 19383 16708 19395 16711
rect 19426 16708 19432 16720
rect 19383 16680 19432 16708
rect 19383 16677 19395 16680
rect 19337 16671 19395 16677
rect 19426 16668 19432 16680
rect 19484 16668 19490 16720
rect 19518 16668 19524 16720
rect 19576 16668 19582 16720
rect 18969 16643 19027 16649
rect 18969 16609 18981 16643
rect 19015 16640 19027 16643
rect 19536 16640 19564 16668
rect 19812 16649 19840 16748
rect 19978 16736 19984 16748
rect 20036 16776 20042 16788
rect 26329 16779 26387 16785
rect 20036 16748 21404 16776
rect 20036 16736 20042 16748
rect 19705 16643 19763 16649
rect 19705 16640 19717 16643
rect 19015 16612 19472 16640
rect 19536 16612 19717 16640
rect 19015 16609 19027 16612
rect 18969 16603 19027 16609
rect 17405 16575 17463 16581
rect 17405 16541 17417 16575
rect 17451 16572 17463 16575
rect 17497 16575 17555 16581
rect 17497 16572 17509 16575
rect 17451 16544 17509 16572
rect 17451 16541 17463 16544
rect 17405 16535 17463 16541
rect 17497 16541 17509 16544
rect 17543 16541 17555 16575
rect 17497 16535 17555 16541
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16541 17739 16575
rect 17681 16535 17739 16541
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16541 18199 16575
rect 18141 16535 18199 16541
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 19061 16575 19119 16581
rect 19061 16541 19073 16575
rect 19107 16572 19119 16575
rect 19334 16572 19340 16584
rect 19107 16544 19340 16572
rect 19107 16541 19119 16544
rect 19061 16535 19119 16541
rect 13710 16476 14320 16504
rect 15028 16476 16887 16504
rect 13710 16473 13722 16476
rect 13664 16467 13722 16473
rect 11609 16439 11667 16445
rect 11609 16436 11621 16439
rect 10980 16408 11621 16436
rect 10597 16399 10655 16405
rect 11609 16405 11621 16408
rect 11655 16405 11667 16439
rect 11609 16399 11667 16405
rect 12434 16396 12440 16448
rect 12492 16396 12498 16448
rect 12529 16439 12587 16445
rect 12529 16405 12541 16439
rect 12575 16436 12587 16439
rect 13078 16436 13084 16448
rect 12575 16408 13084 16436
rect 12575 16405 12587 16408
rect 12529 16399 12587 16405
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 14182 16396 14188 16448
rect 14240 16396 14246 16448
rect 14292 16436 14320 16476
rect 17696 16448 17724 16535
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 19444 16504 19472 16612
rect 19705 16609 19717 16612
rect 19751 16609 19763 16643
rect 19705 16603 19763 16609
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 21376 16581 21404 16748
rect 26329 16745 26341 16779
rect 26375 16776 26387 16779
rect 27890 16776 27896 16788
rect 26375 16748 27896 16776
rect 26375 16745 26387 16748
rect 26329 16739 26387 16745
rect 27890 16736 27896 16748
rect 27948 16736 27954 16788
rect 30650 16776 30656 16788
rect 29840 16748 30656 16776
rect 25222 16708 25228 16720
rect 25148 16680 25228 16708
rect 25038 16600 25044 16652
rect 25096 16600 25102 16652
rect 25148 16649 25176 16680
rect 25222 16668 25228 16680
rect 25280 16668 25286 16720
rect 25133 16643 25191 16649
rect 25133 16609 25145 16643
rect 25179 16609 25191 16643
rect 25133 16603 25191 16609
rect 25317 16643 25375 16649
rect 25317 16609 25329 16643
rect 25363 16640 25375 16643
rect 25406 16640 25412 16652
rect 25363 16612 25412 16640
rect 25363 16609 25375 16612
rect 25317 16603 25375 16609
rect 25406 16600 25412 16612
rect 25464 16640 25470 16652
rect 25464 16612 27660 16640
rect 25464 16600 25470 16612
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16572 19579 16575
rect 21361 16575 21419 16581
rect 19567 16544 20576 16572
rect 19567 16541 19579 16544
rect 19521 16535 19579 16541
rect 20548 16516 20576 16544
rect 21361 16541 21373 16575
rect 21407 16572 21419 16575
rect 22094 16572 22100 16584
rect 21407 16544 22100 16572
rect 21407 16541 21419 16544
rect 21361 16535 21419 16541
rect 22094 16532 22100 16544
rect 22152 16572 22158 16584
rect 23106 16581 23112 16584
rect 22833 16575 22891 16581
rect 22833 16572 22845 16575
rect 22152 16544 22845 16572
rect 22152 16532 22158 16544
rect 22833 16541 22845 16544
rect 22879 16541 22891 16575
rect 23100 16572 23112 16581
rect 23067 16544 23112 16572
rect 22833 16535 22891 16541
rect 23100 16535 23112 16544
rect 23106 16532 23112 16535
rect 23164 16532 23170 16584
rect 25056 16572 25084 16600
rect 27632 16584 27660 16612
rect 27982 16600 27988 16652
rect 28040 16600 28046 16652
rect 29840 16640 29868 16748
rect 30650 16736 30656 16748
rect 30708 16736 30714 16788
rect 31478 16736 31484 16788
rect 31536 16736 31542 16788
rect 37553 16779 37611 16785
rect 37553 16745 37565 16779
rect 37599 16776 37611 16779
rect 37918 16776 37924 16788
rect 37599 16748 37924 16776
rect 37599 16745 37611 16748
rect 37553 16739 37611 16745
rect 37918 16736 37924 16748
rect 37976 16736 37982 16788
rect 29917 16711 29975 16717
rect 29917 16677 29929 16711
rect 29963 16677 29975 16711
rect 29917 16671 29975 16677
rect 29656 16612 29868 16640
rect 29932 16640 29960 16671
rect 31389 16643 31447 16649
rect 29932 16612 30420 16640
rect 25225 16575 25283 16581
rect 25225 16572 25237 16575
rect 25056 16544 25237 16572
rect 25225 16541 25237 16544
rect 25271 16541 25283 16575
rect 25225 16535 25283 16541
rect 25774 16532 25780 16584
rect 25832 16532 25838 16584
rect 25866 16532 25872 16584
rect 25924 16532 25930 16584
rect 26053 16575 26111 16581
rect 26053 16541 26065 16575
rect 26099 16541 26111 16575
rect 26053 16535 26111 16541
rect 26145 16575 26203 16581
rect 26145 16541 26157 16575
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 20042 16507 20100 16513
rect 20042 16504 20054 16507
rect 19444 16476 20054 16504
rect 20042 16473 20054 16476
rect 20088 16473 20100 16507
rect 20042 16467 20100 16473
rect 20530 16464 20536 16516
rect 20588 16464 20594 16516
rect 21628 16507 21686 16513
rect 21628 16473 21640 16507
rect 21674 16504 21686 16507
rect 21818 16504 21824 16516
rect 21674 16476 21824 16504
rect 21674 16473 21686 16476
rect 21628 16467 21686 16473
rect 21818 16464 21824 16476
rect 21876 16464 21882 16516
rect 14829 16439 14887 16445
rect 14829 16436 14841 16439
rect 14292 16408 14841 16436
rect 14829 16405 14841 16408
rect 14875 16405 14887 16439
rect 14829 16399 14887 16405
rect 16022 16396 16028 16448
rect 16080 16396 16086 16448
rect 17678 16396 17684 16448
rect 17736 16396 17742 16448
rect 18966 16396 18972 16448
rect 19024 16436 19030 16448
rect 21174 16436 21180 16448
rect 19024 16408 21180 16436
rect 19024 16396 19030 16408
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 22738 16396 22744 16448
rect 22796 16396 22802 16448
rect 23750 16396 23756 16448
rect 23808 16436 23814 16448
rect 24213 16439 24271 16445
rect 24213 16436 24225 16439
rect 23808 16408 24225 16436
rect 23808 16396 23814 16408
rect 24213 16405 24225 16408
rect 24259 16405 24271 16439
rect 24213 16399 24271 16405
rect 24946 16396 24952 16448
rect 25004 16396 25010 16448
rect 26068 16436 26096 16535
rect 26160 16504 26188 16535
rect 26510 16532 26516 16584
rect 26568 16572 26574 16584
rect 26973 16575 27031 16581
rect 26973 16572 26985 16575
rect 26568 16544 26985 16572
rect 26568 16532 26574 16544
rect 26973 16541 26985 16544
rect 27019 16541 27031 16575
rect 26973 16535 27031 16541
rect 27614 16532 27620 16584
rect 27672 16532 27678 16584
rect 27798 16532 27804 16584
rect 27856 16532 27862 16584
rect 29656 16581 29684 16612
rect 29641 16575 29699 16581
rect 29641 16541 29653 16575
rect 29687 16541 29699 16575
rect 29641 16535 29699 16541
rect 29825 16575 29883 16581
rect 29825 16541 29837 16575
rect 29871 16541 29883 16575
rect 29825 16535 29883 16541
rect 27249 16507 27307 16513
rect 27249 16504 27261 16507
rect 26160 16476 27261 16504
rect 27249 16473 27261 16476
rect 27295 16473 27307 16507
rect 27249 16467 27307 16473
rect 28252 16507 28310 16513
rect 28252 16473 28264 16507
rect 28298 16504 28310 16507
rect 28534 16504 28540 16516
rect 28298 16476 28540 16504
rect 28298 16473 28310 16476
rect 28252 16467 28310 16473
rect 28534 16464 28540 16476
rect 28592 16464 28598 16516
rect 29840 16504 29868 16535
rect 29914 16532 29920 16584
rect 29972 16532 29978 16584
rect 30098 16532 30104 16584
rect 30156 16532 30162 16584
rect 30392 16572 30420 16612
rect 31389 16609 31401 16643
rect 31435 16640 31447 16643
rect 31496 16640 31524 16736
rect 31435 16612 31524 16640
rect 31435 16609 31447 16612
rect 31389 16603 31447 16609
rect 31846 16600 31852 16652
rect 31904 16640 31910 16652
rect 32309 16643 32367 16649
rect 32309 16640 32321 16643
rect 31904 16612 32321 16640
rect 31904 16600 31910 16612
rect 32309 16609 32321 16612
rect 32355 16609 32367 16643
rect 32309 16603 32367 16609
rect 34514 16600 34520 16652
rect 34572 16640 34578 16652
rect 36173 16643 36231 16649
rect 36173 16640 36185 16643
rect 34572 16612 36185 16640
rect 34572 16600 34578 16612
rect 36173 16609 36185 16612
rect 36219 16609 36231 16643
rect 36173 16603 36231 16609
rect 31122 16575 31180 16581
rect 31122 16572 31134 16575
rect 30392 16544 31134 16572
rect 31122 16541 31134 16544
rect 31168 16541 31180 16575
rect 31122 16535 31180 16541
rect 36440 16575 36498 16581
rect 36440 16541 36452 16575
rect 36486 16572 36498 16575
rect 38102 16572 38108 16584
rect 36486 16544 38108 16572
rect 36486 16541 36498 16544
rect 36440 16535 36498 16541
rect 38102 16532 38108 16544
rect 38160 16532 38166 16584
rect 30116 16504 30144 16532
rect 29840 16476 30144 16504
rect 30742 16464 30748 16516
rect 30800 16504 30806 16516
rect 33137 16507 33195 16513
rect 33137 16504 33149 16507
rect 30800 16476 33149 16504
rect 30800 16464 30806 16476
rect 33137 16473 33149 16476
rect 33183 16473 33195 16507
rect 33137 16467 33195 16473
rect 26142 16436 26148 16448
rect 26068 16408 26148 16436
rect 26142 16396 26148 16408
rect 26200 16396 26206 16448
rect 26418 16396 26424 16448
rect 26476 16396 26482 16448
rect 29365 16439 29423 16445
rect 29365 16405 29377 16439
rect 29411 16436 29423 16439
rect 29822 16436 29828 16448
rect 29411 16408 29828 16436
rect 29411 16405 29423 16408
rect 29365 16399 29423 16405
rect 29822 16396 29828 16408
rect 29880 16396 29886 16448
rect 30009 16439 30067 16445
rect 30009 16405 30021 16439
rect 30055 16436 30067 16439
rect 30834 16436 30840 16448
rect 30055 16408 30840 16436
rect 30055 16405 30067 16408
rect 30009 16399 30067 16405
rect 30834 16396 30840 16408
rect 30892 16396 30898 16448
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 9674 16192 9680 16244
rect 9732 16192 9738 16244
rect 10686 16192 10692 16244
rect 10744 16192 10750 16244
rect 11977 16235 12035 16241
rect 11977 16201 11989 16235
rect 12023 16232 12035 16235
rect 12250 16232 12256 16244
rect 12023 16204 12256 16232
rect 12023 16201 12035 16204
rect 11977 16195 12035 16201
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12492 16204 12572 16232
rect 12492 16192 12498 16204
rect 9858 16173 9864 16176
rect 9829 16167 9864 16173
rect 9829 16164 9841 16167
rect 9692 16136 9841 16164
rect 9692 16040 9720 16136
rect 9829 16133 9841 16136
rect 9829 16127 9864 16133
rect 9858 16124 9864 16127
rect 9916 16124 9922 16176
rect 10042 16124 10048 16176
rect 10100 16124 10106 16176
rect 10704 16164 10732 16192
rect 10704 16136 11008 16164
rect 10704 16096 10732 16136
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 10704 16068 10793 16096
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 9674 15988 9680 16040
rect 9732 15988 9738 16040
rect 10888 15960 10916 16059
rect 10980 16028 11008 16136
rect 11072 16136 11560 16164
rect 11072 16105 11100 16136
rect 11532 16108 11560 16136
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11238 16096 11244 16108
rect 11195 16068 11244 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11514 16056 11520 16108
rect 11572 16056 11578 16108
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16065 12311 16099
rect 12253 16059 12311 16065
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16096 12403 16099
rect 12434 16096 12440 16108
rect 12391 16068 12440 16096
rect 12391 16065 12403 16068
rect 12345 16059 12403 16065
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 10980 16000 12081 16028
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 11977 15963 12035 15969
rect 11977 15960 11989 15963
rect 10888 15932 11989 15960
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 9861 15895 9919 15901
rect 9861 15892 9873 15895
rect 9364 15864 9873 15892
rect 9364 15852 9370 15864
rect 9861 15861 9873 15864
rect 9907 15892 9919 15895
rect 10888 15892 10916 15932
rect 11977 15929 11989 15932
rect 12023 15929 12035 15963
rect 12268 15960 12296 16059
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 12544 16105 12572 16204
rect 13078 16192 13084 16244
rect 13136 16192 13142 16244
rect 15105 16235 15163 16241
rect 15105 16201 15117 16235
rect 15151 16232 15163 16235
rect 15746 16232 15752 16244
rect 15151 16204 15752 16232
rect 15151 16201 15163 16204
rect 15105 16195 15163 16201
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 15838 16192 15844 16244
rect 15896 16192 15902 16244
rect 16485 16235 16543 16241
rect 16485 16201 16497 16235
rect 16531 16232 16543 16235
rect 18230 16232 18236 16244
rect 16531 16204 18236 16232
rect 16531 16201 16543 16204
rect 16485 16195 16543 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 18966 16192 18972 16244
rect 19024 16192 19030 16244
rect 19794 16232 19800 16244
rect 19076 16204 19800 16232
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 13096 16096 13124 16192
rect 13173 16099 13231 16105
rect 13173 16096 13185 16099
rect 13096 16068 13185 16096
rect 13173 16065 13185 16068
rect 13219 16065 13231 16099
rect 13173 16059 13231 16065
rect 13262 16056 13268 16108
rect 13320 16056 13326 16108
rect 15105 16099 15163 16105
rect 15105 16065 15117 16099
rect 15151 16096 15163 16099
rect 15856 16096 15884 16192
rect 17678 16164 17684 16176
rect 17604 16136 17684 16164
rect 17604 16105 17632 16136
rect 17678 16124 17684 16136
rect 17736 16164 17742 16176
rect 17957 16167 18015 16173
rect 17957 16164 17969 16167
rect 17736 16136 17969 16164
rect 17736 16124 17742 16136
rect 17957 16133 17969 16136
rect 18003 16133 18015 16167
rect 19076 16164 19104 16204
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 20625 16235 20683 16241
rect 20625 16201 20637 16235
rect 20671 16232 20683 16235
rect 21266 16232 21272 16244
rect 20671 16204 21272 16232
rect 20671 16201 20683 16204
rect 20625 16195 20683 16201
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 21818 16192 21824 16244
rect 21876 16192 21882 16244
rect 22738 16192 22744 16244
rect 22796 16192 22802 16244
rect 24946 16192 24952 16244
rect 25004 16192 25010 16244
rect 26973 16235 27031 16241
rect 26973 16201 26985 16235
rect 27019 16232 27031 16235
rect 27798 16232 27804 16244
rect 27019 16204 27804 16232
rect 27019 16201 27031 16204
rect 26973 16195 27031 16201
rect 27798 16192 27804 16204
rect 27856 16192 27862 16244
rect 27908 16204 28488 16232
rect 17957 16127 18015 16133
rect 18892 16136 19104 16164
rect 19153 16167 19211 16173
rect 15151 16068 15884 16096
rect 16301 16099 16359 16105
rect 15151 16065 15163 16068
rect 15105 16059 15163 16065
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 17589 16099 17647 16105
rect 17589 16096 17601 16099
rect 16347 16068 17601 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 17589 16065 17601 16068
rect 17635 16065 17647 16099
rect 17589 16059 17647 16065
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18414 16096 18420 16108
rect 18095 16068 18420 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 14550 15988 14556 16040
rect 14608 16028 14614 16040
rect 14829 16031 14887 16037
rect 14829 16028 14841 16031
rect 14608 16000 14841 16028
rect 14608 15988 14614 16000
rect 14829 15997 14841 16000
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 15286 15988 15292 16040
rect 15344 16028 15350 16040
rect 15749 16031 15807 16037
rect 15749 16028 15761 16031
rect 15344 16000 15761 16028
rect 15344 15988 15350 16000
rect 15749 15997 15761 16000
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 16117 16031 16175 16037
rect 16117 15997 16129 16031
rect 16163 16028 16175 16031
rect 16574 16028 16580 16040
rect 16163 16000 16580 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 16574 15988 16580 16000
rect 16632 16028 16638 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 16632 16000 16681 16028
rect 16632 15988 16638 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 17770 16028 17776 16040
rect 16669 15991 16727 15997
rect 16776 16000 17776 16028
rect 12526 15960 12532 15972
rect 12268 15932 12532 15960
rect 11977 15923 12035 15929
rect 12526 15920 12532 15932
rect 12584 15920 12590 15972
rect 15013 15963 15071 15969
rect 15013 15929 15025 15963
rect 15059 15960 15071 15963
rect 16022 15960 16028 15972
rect 15059 15932 16028 15960
rect 15059 15929 15071 15932
rect 15013 15923 15071 15929
rect 16022 15920 16028 15932
rect 16080 15920 16086 15972
rect 9907 15864 10916 15892
rect 9907 15861 9919 15864
rect 9861 15855 9919 15861
rect 11330 15852 11336 15904
rect 11388 15852 11394 15904
rect 12158 15852 12164 15904
rect 12216 15852 12222 15904
rect 13722 15852 13728 15904
rect 13780 15852 13786 15904
rect 15194 15852 15200 15904
rect 15252 15852 15258 15904
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 16776 15892 16804 16000
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 16850 15920 16856 15972
rect 16908 15960 16914 15972
rect 17494 15960 17500 15972
rect 16908 15932 17500 15960
rect 16908 15920 16914 15932
rect 17494 15920 17500 15932
rect 17552 15960 17558 15972
rect 17880 15960 17908 16059
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 18892 16105 18920 16136
rect 19153 16133 19165 16167
rect 19199 16164 19211 16167
rect 20806 16164 20812 16176
rect 19199 16136 20812 16164
rect 19199 16133 19211 16136
rect 19153 16127 19211 16133
rect 20806 16124 20812 16136
rect 20864 16124 20870 16176
rect 18877 16099 18935 16105
rect 18877 16065 18889 16099
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 18966 16056 18972 16108
rect 19024 16096 19030 16108
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 19024 16068 19257 16096
rect 19024 16056 19030 16068
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19501 16099 19559 16105
rect 19501 16096 19513 16099
rect 19392 16068 19513 16096
rect 19392 16056 19398 16068
rect 19501 16065 19513 16068
rect 19547 16065 19559 16099
rect 19501 16059 19559 16065
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 20714 16096 20720 16108
rect 19852 16068 20720 16096
rect 19852 16056 19858 16068
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 20990 16096 20996 16108
rect 20947 16068 20996 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 18432 16028 18460 16056
rect 20916 16028 20944 16059
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 21174 16056 21180 16108
rect 21232 16096 21238 16108
rect 21545 16099 21603 16105
rect 21545 16096 21557 16099
rect 21232 16068 21557 16096
rect 21232 16056 21238 16068
rect 21545 16065 21557 16068
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 22756 16096 22784 16192
rect 24964 16164 24992 16192
rect 25102 16167 25160 16173
rect 25102 16164 25114 16167
rect 24964 16136 25114 16164
rect 25102 16133 25114 16136
rect 25148 16133 25160 16167
rect 25102 16127 25160 16133
rect 25222 16124 25228 16176
rect 25280 16124 25286 16176
rect 23109 16099 23167 16105
rect 23109 16096 23121 16099
rect 22756 16068 23121 16096
rect 23109 16065 23121 16068
rect 23155 16096 23167 16099
rect 23290 16096 23296 16108
rect 23155 16068 23296 16096
rect 23155 16065 23167 16068
rect 23109 16059 23167 16065
rect 23290 16056 23296 16068
rect 23348 16056 23354 16108
rect 25240 16096 25268 16124
rect 24872 16068 25268 16096
rect 18432 16000 19288 16028
rect 17552 15932 17908 15960
rect 17552 15920 17558 15932
rect 19058 15920 19064 15972
rect 19116 15960 19122 15972
rect 19153 15963 19211 15969
rect 19153 15960 19165 15963
rect 19116 15932 19165 15960
rect 19116 15920 19122 15932
rect 19153 15929 19165 15932
rect 19199 15929 19211 15963
rect 19153 15923 19211 15929
rect 15712 15864 16804 15892
rect 15712 15852 15718 15864
rect 17310 15852 17316 15904
rect 17368 15852 17374 15904
rect 17402 15852 17408 15904
rect 17460 15852 17466 15904
rect 19260 15892 19288 16000
rect 20364 16000 20944 16028
rect 20364 15892 20392 16000
rect 23934 15988 23940 16040
rect 23992 15988 23998 16040
rect 24872 16037 24900 16068
rect 26878 16056 26884 16108
rect 26936 16096 26942 16108
rect 27908 16096 27936 16204
rect 27982 16124 27988 16176
rect 28040 16164 28046 16176
rect 28040 16136 28396 16164
rect 28040 16124 28046 16136
rect 26936 16068 27936 16096
rect 28097 16099 28155 16105
rect 26936 16056 26942 16068
rect 28097 16065 28109 16099
rect 28143 16096 28155 16099
rect 28258 16096 28264 16108
rect 28143 16068 28264 16096
rect 28143 16065 28155 16068
rect 28097 16059 28155 16065
rect 28258 16056 28264 16068
rect 28316 16056 28322 16108
rect 28368 16105 28396 16136
rect 28460 16105 28488 16204
rect 28534 16192 28540 16244
rect 28592 16192 28598 16244
rect 29914 16192 29920 16244
rect 29972 16192 29978 16244
rect 34790 16232 34796 16244
rect 30116 16204 30692 16232
rect 28353 16099 28411 16105
rect 28353 16065 28365 16099
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 28445 16099 28503 16105
rect 28445 16065 28457 16099
rect 28491 16065 28503 16099
rect 28445 16059 28503 16065
rect 28629 16099 28687 16105
rect 28629 16065 28641 16099
rect 28675 16065 28687 16099
rect 29932 16096 29960 16192
rect 30116 16176 30144 16204
rect 30098 16124 30104 16176
rect 30156 16124 30162 16176
rect 30285 16167 30343 16173
rect 30285 16133 30297 16167
rect 30331 16164 30343 16167
rect 30561 16167 30619 16173
rect 30561 16164 30573 16167
rect 30331 16136 30573 16164
rect 30331 16133 30343 16136
rect 30285 16127 30343 16133
rect 30561 16133 30573 16136
rect 30607 16133 30619 16167
rect 30561 16127 30619 16133
rect 30664 16105 30692 16204
rect 31726 16204 34796 16232
rect 31726 16164 31754 16204
rect 34790 16192 34796 16204
rect 34848 16192 34854 16244
rect 35342 16192 35348 16244
rect 35400 16192 35406 16244
rect 31036 16136 31754 16164
rect 30377 16099 30435 16105
rect 30377 16096 30389 16099
rect 29932 16068 30389 16096
rect 28629 16059 28687 16065
rect 30377 16065 30389 16068
rect 30423 16065 30435 16099
rect 30377 16059 30435 16065
rect 30653 16099 30711 16105
rect 30653 16065 30665 16099
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 30745 16099 30803 16105
rect 30745 16065 30757 16099
rect 30791 16065 30803 16099
rect 30745 16059 30803 16065
rect 30929 16099 30987 16105
rect 30929 16065 30941 16099
rect 30975 16065 30987 16099
rect 30929 16059 30987 16065
rect 24857 16031 24915 16037
rect 24857 15997 24869 16031
rect 24903 15997 24915 16031
rect 24857 15991 24915 15997
rect 20438 15920 20444 15972
rect 20496 15960 20502 15972
rect 20993 15963 21051 15969
rect 20993 15960 21005 15963
rect 20496 15932 21005 15960
rect 20496 15920 20502 15932
rect 20993 15929 21005 15932
rect 21039 15929 21051 15963
rect 28644 15960 28672 16059
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 16028 29791 16031
rect 29822 16028 29828 16040
rect 29779 16000 29828 16028
rect 29779 15997 29791 16000
rect 29733 15991 29791 15997
rect 29822 15988 29828 16000
rect 29880 16028 29886 16040
rect 30760 16028 30788 16059
rect 29880 16000 30788 16028
rect 29880 15988 29886 16000
rect 30834 15988 30840 16040
rect 30892 16028 30898 16040
rect 30944 16028 30972 16059
rect 30892 16000 30972 16028
rect 30892 15988 30898 16000
rect 30377 15963 30435 15969
rect 30377 15960 30389 15963
rect 28644 15932 30389 15960
rect 20993 15923 21051 15929
rect 30377 15929 30389 15932
rect 30423 15929 30435 15963
rect 31036 15960 31064 16136
rect 31754 16056 31760 16108
rect 31812 16096 31818 16108
rect 32309 16099 32367 16105
rect 32309 16096 32321 16099
rect 31812 16068 32321 16096
rect 31812 16056 31818 16068
rect 32309 16065 32321 16068
rect 32355 16065 32367 16099
rect 33410 16096 33416 16108
rect 32309 16059 32367 16065
rect 32508 16068 33416 16096
rect 31478 15988 31484 16040
rect 31536 16028 31542 16040
rect 32508 16028 32536 16068
rect 33410 16056 33416 16068
rect 33468 16056 33474 16108
rect 33680 16099 33738 16105
rect 33680 16065 33692 16099
rect 33726 16096 33738 16099
rect 34054 16096 34060 16108
rect 33726 16068 34060 16096
rect 33726 16065 33738 16068
rect 33680 16059 33738 16065
rect 34054 16056 34060 16068
rect 34112 16056 34118 16108
rect 34606 16056 34612 16108
rect 34664 16096 34670 16108
rect 34885 16099 34943 16105
rect 34885 16096 34897 16099
rect 34664 16068 34897 16096
rect 34664 16056 34670 16068
rect 34885 16065 34897 16068
rect 34931 16065 34943 16099
rect 34885 16059 34943 16065
rect 35404 16099 35462 16105
rect 35404 16065 35416 16099
rect 35450 16096 35462 16099
rect 35450 16068 37412 16096
rect 35450 16065 35462 16068
rect 35404 16059 35462 16065
rect 31536 16000 32536 16028
rect 32585 16031 32643 16037
rect 31536 15988 31542 16000
rect 32585 15997 32597 16031
rect 32631 16028 32643 16031
rect 32677 16031 32735 16037
rect 32677 16028 32689 16031
rect 32631 16000 32689 16028
rect 32631 15997 32643 16000
rect 32585 15991 32643 15997
rect 32677 15997 32689 16000
rect 32723 15997 32735 16031
rect 32677 15991 32735 15997
rect 33321 16031 33379 16037
rect 33321 15997 33333 16031
rect 33367 15997 33379 16031
rect 33321 15991 33379 15997
rect 30377 15923 30435 15929
rect 30484 15932 31064 15960
rect 19260 15864 20392 15892
rect 20530 15852 20536 15904
rect 20588 15892 20594 15904
rect 20717 15895 20775 15901
rect 20717 15892 20729 15895
rect 20588 15864 20729 15892
rect 20588 15852 20594 15864
rect 20717 15861 20729 15864
rect 20763 15861 20775 15895
rect 20717 15855 20775 15861
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 21450 15892 21456 15904
rect 20864 15864 21456 15892
rect 20864 15852 20870 15864
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 22554 15852 22560 15904
rect 22612 15852 22618 15904
rect 23382 15852 23388 15904
rect 23440 15852 23446 15904
rect 25866 15852 25872 15904
rect 25924 15892 25930 15904
rect 26237 15895 26295 15901
rect 26237 15892 26249 15895
rect 25924 15864 26249 15892
rect 25924 15852 25930 15864
rect 26237 15861 26249 15864
rect 26283 15892 26295 15895
rect 26970 15892 26976 15904
rect 26283 15864 26976 15892
rect 26283 15861 26295 15864
rect 26237 15855 26295 15861
rect 26970 15852 26976 15864
rect 27028 15852 27034 15904
rect 27154 15852 27160 15904
rect 27212 15892 27218 15904
rect 30484 15892 30512 15932
rect 33336 15904 33364 15991
rect 34698 15920 34704 15972
rect 34756 15960 34762 15972
rect 35529 15963 35587 15969
rect 35529 15960 35541 15963
rect 34756 15932 35541 15960
rect 34756 15920 34762 15932
rect 35529 15929 35541 15932
rect 35575 15929 35587 15963
rect 35529 15923 35587 15929
rect 37384 15904 37412 16068
rect 27212 15864 30512 15892
rect 27212 15852 27218 15864
rect 30742 15852 30748 15904
rect 30800 15852 30806 15904
rect 32030 15852 32036 15904
rect 32088 15892 32094 15904
rect 32125 15895 32183 15901
rect 32125 15892 32137 15895
rect 32088 15864 32137 15892
rect 32088 15852 32094 15864
rect 32125 15861 32137 15864
rect 32171 15861 32183 15895
rect 32125 15855 32183 15861
rect 32490 15852 32496 15904
rect 32548 15852 32554 15904
rect 33318 15852 33324 15904
rect 33376 15852 33382 15904
rect 34606 15852 34612 15904
rect 34664 15892 34670 15904
rect 34977 15895 35035 15901
rect 34977 15892 34989 15895
rect 34664 15864 34989 15892
rect 34664 15852 34670 15864
rect 34977 15861 34989 15864
rect 35023 15861 35035 15895
rect 34977 15855 35035 15861
rect 37366 15852 37372 15904
rect 37424 15852 37430 15904
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 11054 15648 11060 15700
rect 11112 15648 11118 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 11256 15660 11621 15688
rect 9490 15580 9496 15632
rect 9548 15620 9554 15632
rect 11072 15620 11100 15648
rect 9548 15592 11100 15620
rect 9548 15580 9554 15592
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15552 8815 15555
rect 9582 15552 9588 15564
rect 8803 15524 9588 15552
rect 8803 15521 8815 15524
rect 8757 15515 8815 15521
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 7006 15444 7012 15496
rect 7064 15444 7070 15496
rect 9968 15493 9996 15592
rect 11146 15580 11152 15632
rect 11204 15580 11210 15632
rect 11256 15496 11284 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 11977 15691 12035 15697
rect 11977 15657 11989 15691
rect 12023 15688 12035 15691
rect 12158 15688 12164 15700
rect 12023 15660 12164 15688
rect 12023 15657 12035 15660
rect 11977 15651 12035 15657
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 16022 15648 16028 15700
rect 16080 15648 16086 15700
rect 17696 15660 19288 15688
rect 14182 15552 14188 15564
rect 11716 15524 14188 15552
rect 9953 15487 10011 15493
rect 9953 15453 9965 15487
rect 9999 15453 10011 15487
rect 9953 15447 10011 15453
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 7282 15376 7288 15428
rect 7340 15376 7346 15428
rect 8570 15416 8576 15428
rect 8510 15388 8576 15416
rect 8570 15376 8576 15388
rect 8628 15376 8634 15428
rect 9401 15419 9459 15425
rect 9401 15385 9413 15419
rect 9447 15416 9459 15419
rect 10045 15419 10103 15425
rect 10045 15416 10057 15419
rect 9447 15388 10057 15416
rect 9447 15385 9459 15388
rect 9401 15379 9459 15385
rect 10045 15385 10057 15388
rect 10091 15385 10103 15419
rect 10045 15379 10103 15385
rect 10980 15416 11008 15447
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 11238 15444 11244 15496
rect 11296 15444 11302 15496
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15484 11391 15487
rect 11514 15484 11520 15496
rect 11379 15456 11520 15484
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 11716 15494 11744 15524
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 11624 15493 11744 15494
rect 11609 15487 11744 15493
rect 11609 15453 11621 15487
rect 11655 15466 11744 15487
rect 11793 15487 11851 15493
rect 11655 15453 11667 15466
rect 11609 15447 11667 15453
rect 11793 15453 11805 15487
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 11808 15416 11836 15447
rect 15194 15444 15200 15496
rect 15252 15493 15258 15496
rect 15252 15484 15264 15493
rect 15252 15456 15297 15484
rect 15252 15447 15264 15456
rect 15252 15444 15258 15447
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 15436 15456 15485 15484
rect 15436 15444 15442 15456
rect 15473 15453 15485 15456
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 15841 15487 15899 15493
rect 15841 15453 15853 15487
rect 15887 15484 15899 15487
rect 16040 15484 16068 15648
rect 17696 15564 17724 15660
rect 17586 15512 17592 15564
rect 17644 15512 17650 15564
rect 17678 15512 17684 15564
rect 17736 15512 17742 15564
rect 19260 15561 19288 15660
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 21726 15688 21732 15700
rect 20312 15660 21732 15688
rect 20312 15648 20318 15660
rect 21726 15648 21732 15660
rect 21784 15648 21790 15700
rect 22554 15648 22560 15700
rect 22612 15648 22618 15700
rect 23198 15648 23204 15700
rect 23256 15648 23262 15700
rect 23382 15648 23388 15700
rect 23440 15648 23446 15700
rect 26602 15648 26608 15700
rect 26660 15688 26666 15700
rect 26881 15691 26939 15697
rect 26881 15688 26893 15691
rect 26660 15660 26893 15688
rect 26660 15648 26666 15660
rect 26881 15657 26893 15660
rect 26927 15657 26939 15691
rect 26881 15651 26939 15657
rect 27798 15648 27804 15700
rect 27856 15648 27862 15700
rect 29914 15648 29920 15700
rect 29972 15688 29978 15700
rect 31481 15691 31539 15697
rect 31481 15688 31493 15691
rect 29972 15660 31493 15688
rect 29972 15648 29978 15660
rect 31481 15657 31493 15660
rect 31527 15688 31539 15691
rect 32490 15688 32496 15700
rect 31527 15660 32496 15688
rect 31527 15657 31539 15660
rect 31481 15651 31539 15657
rect 32490 15648 32496 15660
rect 32548 15648 32554 15700
rect 34054 15648 34060 15700
rect 34112 15688 34118 15700
rect 34149 15691 34207 15697
rect 34149 15688 34161 15691
rect 34112 15660 34161 15688
rect 34112 15648 34118 15660
rect 34149 15657 34161 15660
rect 34195 15657 34207 15691
rect 34149 15651 34207 15657
rect 34698 15648 34704 15700
rect 34756 15648 34762 15700
rect 35342 15648 35348 15700
rect 35400 15688 35406 15700
rect 36357 15691 36415 15697
rect 36357 15688 36369 15691
rect 35400 15660 36369 15688
rect 35400 15648 35406 15660
rect 36357 15657 36369 15660
rect 36403 15657 36415 15691
rect 36357 15651 36415 15657
rect 19245 15555 19303 15561
rect 19245 15521 19257 15555
rect 19291 15552 19303 15555
rect 19518 15552 19524 15564
rect 19291 15524 19524 15552
rect 19291 15521 19303 15524
rect 19245 15515 19303 15521
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 19794 15512 19800 15564
rect 19852 15512 19858 15564
rect 19889 15555 19947 15561
rect 19889 15521 19901 15555
rect 19935 15552 19947 15555
rect 20349 15555 20407 15561
rect 20349 15552 20361 15555
rect 19935 15524 20361 15552
rect 19935 15521 19947 15524
rect 19889 15515 19947 15521
rect 20349 15521 20361 15524
rect 20395 15521 20407 15555
rect 20349 15515 20407 15521
rect 21174 15512 21180 15564
rect 21232 15512 21238 15564
rect 22005 15555 22063 15561
rect 22005 15521 22017 15555
rect 22051 15552 22063 15555
rect 22572 15552 22600 15648
rect 23400 15552 23428 15648
rect 27816 15552 27844 15648
rect 30834 15620 30840 15632
rect 29840 15592 30840 15620
rect 29840 15552 29868 15592
rect 30834 15580 30840 15592
rect 30892 15620 30898 15632
rect 34716 15620 34744 15648
rect 30892 15592 31340 15620
rect 30892 15580 30898 15592
rect 22051 15524 22600 15552
rect 23216 15524 23428 15552
rect 26712 15524 27844 15552
rect 29748 15524 29868 15552
rect 29917 15555 29975 15561
rect 22051 15521 22063 15524
rect 22005 15515 22063 15521
rect 15887 15456 16068 15484
rect 17604 15484 17632 15512
rect 18966 15484 18972 15496
rect 17604 15456 18972 15484
rect 15887 15453 15899 15456
rect 15841 15447 15899 15453
rect 18966 15444 18972 15456
rect 19024 15484 19030 15496
rect 19061 15487 19119 15493
rect 19061 15484 19073 15487
rect 19024 15456 19073 15484
rect 19024 15444 19030 15456
rect 19061 15453 19073 15456
rect 19107 15484 19119 15487
rect 19702 15484 19708 15496
rect 19107 15456 19708 15484
rect 19107 15453 19119 15456
rect 19061 15447 19119 15453
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 19812 15484 19840 15512
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 19812 15456 20177 15484
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20254 15444 20260 15496
rect 20312 15444 20318 15496
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15453 20499 15487
rect 20441 15447 20499 15453
rect 14182 15416 14188 15428
rect 10980 15388 11836 15416
rect 11900 15388 14188 15416
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 9490 15308 9496 15360
rect 9548 15308 9554 15360
rect 9582 15308 9588 15360
rect 9640 15348 9646 15360
rect 10980 15348 11008 15388
rect 9640 15320 11008 15348
rect 9640 15308 9646 15320
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 11900 15348 11928 15388
rect 14182 15376 14188 15388
rect 14240 15376 14246 15428
rect 14550 15376 14556 15428
rect 14608 15416 14614 15428
rect 16574 15416 16580 15428
rect 14608 15388 16580 15416
rect 14608 15376 14614 15388
rect 11572 15320 11928 15348
rect 11572 15308 11578 15320
rect 14090 15308 14096 15360
rect 14148 15308 14154 15360
rect 15746 15308 15752 15360
rect 15804 15308 15810 15360
rect 16224 15357 16252 15388
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 17344 15419 17402 15425
rect 17344 15385 17356 15419
rect 17390 15416 17402 15419
rect 17494 15416 17500 15428
rect 17390 15388 17500 15416
rect 17390 15385 17402 15388
rect 17344 15379 17402 15385
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 18816 15419 18874 15425
rect 18816 15385 18828 15419
rect 18862 15416 18874 15419
rect 18862 15388 19012 15416
rect 18862 15385 18874 15388
rect 18816 15379 18874 15385
rect 16209 15351 16267 15357
rect 16209 15317 16221 15351
rect 16255 15317 16267 15351
rect 16209 15311 16267 15317
rect 17678 15308 17684 15360
rect 17736 15308 17742 15360
rect 18984 15348 19012 15388
rect 19444 15388 20024 15416
rect 19444 15348 19472 15388
rect 19996 15357 20024 15388
rect 18984 15320 19472 15348
rect 19981 15351 20039 15357
rect 19981 15317 19993 15351
rect 20027 15317 20039 15351
rect 19981 15311 20039 15317
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 20456 15348 20484 15447
rect 21450 15444 21456 15496
rect 21508 15486 21514 15496
rect 21546 15487 21604 15493
rect 21546 15486 21558 15487
rect 21508 15458 21558 15486
rect 21508 15444 21514 15458
rect 21546 15453 21558 15458
rect 21592 15453 21604 15487
rect 21546 15447 21604 15453
rect 21726 15444 21732 15496
rect 21784 15444 21790 15496
rect 22097 15487 22155 15493
rect 22097 15453 22109 15487
rect 22143 15484 22155 15487
rect 22143 15456 22324 15484
rect 22143 15453 22155 15456
rect 22097 15447 22155 15453
rect 21634 15376 21640 15428
rect 21692 15376 21698 15428
rect 21867 15419 21925 15425
rect 21867 15385 21879 15419
rect 21913 15416 21925 15419
rect 22186 15416 22192 15428
rect 21913 15388 22192 15416
rect 21913 15385 21925 15388
rect 21867 15379 21925 15385
rect 22186 15376 22192 15388
rect 22244 15376 22250 15428
rect 20128 15320 20484 15348
rect 20128 15308 20134 15320
rect 20622 15308 20628 15360
rect 20680 15308 20686 15360
rect 21361 15351 21419 15357
rect 21361 15317 21373 15351
rect 21407 15348 21419 15351
rect 22296 15348 22324 15456
rect 22646 15444 22652 15496
rect 22704 15444 22710 15496
rect 23014 15444 23020 15496
rect 23072 15444 23078 15496
rect 23216 15493 23244 15524
rect 23201 15487 23259 15493
rect 23201 15453 23213 15487
rect 23247 15453 23259 15487
rect 23201 15447 23259 15453
rect 23290 15444 23296 15496
rect 23348 15444 23354 15496
rect 23474 15444 23480 15496
rect 23532 15484 23538 15496
rect 23934 15484 23940 15496
rect 23532 15456 23940 15484
rect 23532 15444 23538 15456
rect 23934 15444 23940 15456
rect 23992 15484 23998 15496
rect 24121 15487 24179 15493
rect 24121 15484 24133 15487
rect 23992 15456 24133 15484
rect 23992 15444 23998 15456
rect 24121 15453 24133 15456
rect 24167 15453 24179 15487
rect 24121 15447 24179 15453
rect 24397 15487 24455 15493
rect 24397 15453 24409 15487
rect 24443 15484 24455 15487
rect 25130 15484 25136 15496
rect 24443 15456 25136 15484
rect 24443 15453 24455 15456
rect 24397 15447 24455 15453
rect 22664 15416 22692 15444
rect 24872 15428 24900 15456
rect 25130 15444 25136 15456
rect 25188 15444 25194 15496
rect 25682 15444 25688 15496
rect 25740 15484 25746 15496
rect 26712 15493 26740 15524
rect 26329 15487 26387 15493
rect 26329 15484 26341 15487
rect 25740 15456 26341 15484
rect 25740 15444 25746 15456
rect 26329 15453 26341 15456
rect 26375 15453 26387 15487
rect 26329 15447 26387 15453
rect 26697 15487 26755 15493
rect 26697 15453 26709 15487
rect 26743 15453 26755 15487
rect 26697 15447 26755 15453
rect 26970 15444 26976 15496
rect 27028 15444 27034 15496
rect 27798 15444 27804 15496
rect 27856 15444 27862 15496
rect 29748 15493 29776 15524
rect 29917 15521 29929 15555
rect 29963 15552 29975 15555
rect 30098 15552 30104 15564
rect 29963 15524 30104 15552
rect 29963 15521 29975 15524
rect 29917 15515 29975 15521
rect 30098 15512 30104 15524
rect 30156 15512 30162 15564
rect 30742 15512 30748 15564
rect 30800 15552 30806 15564
rect 30800 15524 31064 15552
rect 30800 15512 30806 15524
rect 29733 15487 29791 15493
rect 29733 15453 29745 15487
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 29822 15444 29828 15496
rect 29880 15444 29886 15496
rect 30006 15444 30012 15496
rect 30064 15484 30070 15496
rect 31036 15493 31064 15524
rect 31312 15496 31340 15592
rect 34164 15592 34744 15620
rect 30285 15487 30343 15493
rect 30285 15484 30297 15487
rect 30064 15456 30297 15484
rect 30064 15444 30070 15456
rect 30285 15453 30297 15456
rect 30331 15453 30343 15487
rect 30285 15447 30343 15453
rect 31021 15487 31079 15493
rect 31021 15453 31033 15487
rect 31067 15453 31079 15487
rect 31021 15447 31079 15453
rect 23385 15419 23443 15425
rect 23385 15416 23397 15419
rect 22664 15388 23397 15416
rect 23385 15385 23397 15388
rect 23431 15385 23443 15419
rect 23385 15379 23443 15385
rect 24486 15376 24492 15428
rect 24544 15416 24550 15428
rect 24642 15419 24700 15425
rect 24642 15416 24654 15419
rect 24544 15388 24654 15416
rect 24544 15376 24550 15388
rect 24642 15385 24654 15388
rect 24688 15385 24700 15419
rect 24642 15379 24700 15385
rect 24854 15376 24860 15428
rect 24912 15376 24918 15428
rect 25314 15376 25320 15428
rect 25372 15416 25378 15428
rect 25700 15416 25728 15444
rect 25372 15388 25728 15416
rect 25372 15376 25378 15388
rect 26510 15376 26516 15428
rect 26568 15376 26574 15428
rect 26605 15419 26663 15425
rect 26605 15385 26617 15419
rect 26651 15416 26663 15419
rect 29840 15416 29868 15444
rect 30300 15416 30328 15447
rect 31294 15444 31300 15496
rect 31352 15444 31358 15496
rect 31478 15444 31484 15496
rect 31536 15484 31542 15496
rect 32030 15493 32036 15496
rect 31757 15487 31815 15493
rect 31757 15484 31769 15487
rect 31536 15456 31769 15484
rect 31536 15444 31542 15456
rect 31757 15453 31769 15456
rect 31803 15453 31815 15487
rect 32024 15484 32036 15493
rect 31991 15456 32036 15484
rect 31757 15447 31815 15453
rect 32024 15447 32036 15456
rect 32030 15444 32036 15447
rect 32088 15444 32094 15496
rect 33778 15444 33784 15496
rect 33836 15444 33842 15496
rect 33870 15444 33876 15496
rect 33928 15484 33934 15496
rect 34164 15493 34192 15592
rect 34977 15555 35035 15561
rect 34977 15552 34989 15555
rect 34348 15524 34989 15552
rect 34348 15496 34376 15524
rect 34977 15521 34989 15524
rect 35023 15521 35035 15555
rect 36372 15552 36400 15651
rect 37001 15555 37059 15561
rect 37001 15552 37013 15555
rect 36372 15524 37013 15552
rect 34977 15515 35035 15521
rect 37001 15521 37013 15524
rect 37047 15521 37059 15555
rect 37001 15515 37059 15521
rect 33965 15487 34023 15493
rect 33965 15484 33977 15487
rect 33928 15456 33977 15484
rect 33928 15444 33934 15456
rect 33965 15453 33977 15456
rect 34011 15453 34023 15487
rect 33965 15447 34023 15453
rect 34149 15487 34207 15493
rect 34149 15453 34161 15487
rect 34195 15453 34207 15487
rect 34149 15447 34207 15453
rect 34241 15487 34299 15493
rect 34241 15453 34253 15487
rect 34287 15453 34299 15487
rect 34241 15447 34299 15453
rect 31113 15419 31171 15425
rect 31113 15416 31125 15419
rect 26651 15388 26685 15416
rect 29840 15388 29960 15416
rect 30300 15388 31125 15416
rect 26651 15385 26663 15388
rect 26605 15379 26663 15385
rect 21407 15320 22324 15348
rect 21407 15317 21419 15320
rect 21361 15311 21419 15317
rect 22738 15308 22744 15360
rect 22796 15308 22802 15360
rect 23566 15308 23572 15360
rect 23624 15308 23630 15360
rect 25777 15351 25835 15357
rect 25777 15317 25789 15351
rect 25823 15348 25835 15351
rect 26620 15348 26648 15379
rect 29932 15360 29960 15388
rect 31113 15385 31125 15388
rect 31159 15385 31171 15419
rect 33318 15416 33324 15428
rect 31113 15379 31171 15385
rect 33152 15388 33324 15416
rect 26786 15348 26792 15360
rect 25823 15320 26792 15348
rect 25823 15317 25835 15320
rect 25777 15311 25835 15317
rect 26786 15308 26792 15320
rect 26844 15308 26850 15360
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 27617 15351 27675 15357
rect 27617 15348 27629 15351
rect 27580 15320 27629 15348
rect 27580 15308 27586 15320
rect 27617 15317 27629 15320
rect 27663 15317 27675 15351
rect 27617 15311 27675 15317
rect 28442 15308 28448 15360
rect 28500 15308 28506 15360
rect 29546 15308 29552 15360
rect 29604 15308 29610 15360
rect 29914 15308 29920 15360
rect 29972 15308 29978 15360
rect 30926 15308 30932 15360
rect 30984 15308 30990 15360
rect 33152 15357 33180 15388
rect 33318 15376 33324 15388
rect 33376 15416 33382 15428
rect 34256 15416 34284 15447
rect 34330 15444 34336 15496
rect 34388 15444 34394 15496
rect 34606 15444 34612 15496
rect 34664 15444 34670 15496
rect 34701 15487 34759 15493
rect 34701 15453 34713 15487
rect 34747 15484 34759 15487
rect 34790 15484 34796 15496
rect 34747 15456 34796 15484
rect 34747 15453 34759 15456
rect 34701 15447 34759 15453
rect 34790 15444 34796 15456
rect 34848 15444 34854 15496
rect 37366 15444 37372 15496
rect 37424 15484 37430 15496
rect 68278 15484 68284 15496
rect 37424 15456 68284 15484
rect 37424 15444 37430 15456
rect 68278 15444 68284 15456
rect 68336 15444 68342 15496
rect 33376 15388 34284 15416
rect 33376 15376 33382 15388
rect 33137 15351 33195 15357
rect 33137 15317 33149 15351
rect 33183 15317 33195 15351
rect 33137 15311 33195 15317
rect 33226 15308 33232 15360
rect 33284 15308 33290 15360
rect 33686 15308 33692 15360
rect 33744 15348 33750 15360
rect 34333 15351 34391 15357
rect 34333 15348 34345 15351
rect 33744 15320 34345 15348
rect 33744 15308 33750 15320
rect 34333 15317 34345 15320
rect 34379 15317 34391 15351
rect 34624 15348 34652 15444
rect 35244 15419 35302 15425
rect 35244 15385 35256 15419
rect 35290 15416 35302 15419
rect 35342 15416 35348 15428
rect 35290 15388 35348 15416
rect 35290 15385 35302 15388
rect 35244 15379 35302 15385
rect 35342 15376 35348 15388
rect 35400 15376 35406 15428
rect 34793 15351 34851 15357
rect 34793 15348 34805 15351
rect 34624 15320 34805 15348
rect 34333 15311 34391 15317
rect 34793 15317 34805 15320
rect 34839 15317 34851 15351
rect 34793 15311 34851 15317
rect 36446 15308 36452 15360
rect 36504 15308 36510 15360
rect 37274 15308 37280 15360
rect 37332 15308 37338 15360
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 7929 15147 7987 15153
rect 7929 15144 7941 15147
rect 7340 15116 7941 15144
rect 7340 15104 7346 15116
rect 7929 15113 7941 15116
rect 7975 15113 7987 15147
rect 7929 15107 7987 15113
rect 8570 15104 8576 15156
rect 8628 15104 8634 15156
rect 9030 15104 9036 15156
rect 9088 15104 9094 15156
rect 9674 15104 9680 15156
rect 9732 15104 9738 15156
rect 12618 15144 12624 15156
rect 11808 15116 12624 15144
rect 9048 15076 9076 15104
rect 8128 15048 9076 15076
rect 8128 15017 8156 15048
rect 9582 15036 9588 15088
rect 9640 15036 9646 15088
rect 9845 15079 9903 15085
rect 9845 15045 9857 15079
rect 9891 15076 9903 15079
rect 9950 15076 9956 15088
rect 9891 15048 9956 15076
rect 9891 15045 9903 15048
rect 9845 15039 9903 15045
rect 9950 15036 9956 15048
rect 10008 15036 10014 15088
rect 10045 15079 10103 15085
rect 10045 15045 10057 15079
rect 10091 15045 10103 15079
rect 10045 15039 10103 15045
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 8662 14968 8668 15020
rect 8720 14968 8726 15020
rect 9600 15008 9628 15036
rect 10060 15008 10088 15039
rect 11330 15036 11336 15088
rect 11388 15076 11394 15088
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 11388 15048 11529 15076
rect 11388 15036 11394 15048
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 11517 15039 11575 15045
rect 9600 14980 10088 15008
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 11808 15017 11836 15116
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 13265 15147 13323 15153
rect 13265 15144 13277 15147
rect 12768 15116 13277 15144
rect 12768 15104 12774 15116
rect 13265 15113 13277 15116
rect 13311 15113 13323 15147
rect 13265 15107 13323 15113
rect 14182 15104 14188 15156
rect 14240 15104 14246 15156
rect 14752 15116 15884 15144
rect 11882 15036 11888 15088
rect 11940 15076 11946 15088
rect 11940 15048 12204 15076
rect 11940 15036 11946 15048
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11204 14980 11713 15008
rect 11204 14968 11210 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 14977 11851 15011
rect 12069 15011 12127 15017
rect 12069 15008 12081 15011
rect 11793 14971 11851 14977
rect 11992 14980 12081 15008
rect 11992 14881 12020 14980
rect 12069 14977 12081 14980
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 11977 14875 12035 14881
rect 11977 14841 11989 14875
rect 12023 14841 12035 14875
rect 12176 14872 12204 15048
rect 12250 15036 12256 15088
rect 12308 15076 12314 15088
rect 12308 15048 13768 15076
rect 12308 15036 12314 15048
rect 12529 15014 12587 15017
rect 12529 15011 12756 15014
rect 12529 14977 12541 15011
rect 12575 15008 12756 15011
rect 12894 15008 12900 15020
rect 12575 14986 12900 15008
rect 12575 14980 12596 14986
rect 12728 14980 12900 14986
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 12986 14968 12992 15020
rect 13044 15008 13050 15020
rect 13740 15017 13768 15048
rect 14090 15036 14096 15088
rect 14148 15076 14154 15088
rect 14148 15048 14688 15076
rect 14148 15036 14154 15048
rect 14292 15017 14320 15048
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 13044 14980 13093 15008
rect 13044 14968 13050 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 13081 14971 13139 14977
rect 13188 14980 13553 15008
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 12768 14912 12817 14940
rect 12768 14900 12774 14912
rect 12805 14909 12817 14912
rect 12851 14940 12863 14943
rect 13188 14940 13216 14980
rect 13541 14977 13553 14980
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14550 14968 14556 15020
rect 14608 14968 14614 15020
rect 14660 15017 14688 15048
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 12851 14912 13216 14940
rect 13449 14943 13507 14949
rect 12851 14909 12863 14912
rect 12805 14903 12863 14909
rect 13449 14909 13461 14943
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14909 13691 14943
rect 14752 14940 14780 15116
rect 14844 15048 15792 15076
rect 14844 15017 14872 15048
rect 15764 15020 15792 15048
rect 15856 15020 15884 15116
rect 15930 15104 15936 15156
rect 15988 15144 15994 15156
rect 15988 15116 16988 15144
rect 15988 15104 15994 15116
rect 16485 15079 16543 15085
rect 16485 15045 16497 15079
rect 16531 15076 16543 15079
rect 16853 15079 16911 15085
rect 16853 15076 16865 15079
rect 16531 15048 16865 15076
rect 16531 15045 16543 15048
rect 16485 15039 16543 15045
rect 16853 15045 16865 15048
rect 16899 15045 16911 15079
rect 16853 15039 16911 15045
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 14977 14887 15011
rect 14829 14971 14887 14977
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 14977 15071 15011
rect 15013 14971 15071 14977
rect 13633 14903 13691 14909
rect 14660 14912 14780 14940
rect 15028 14940 15056 14971
rect 15746 14968 15752 15020
rect 15804 14968 15810 15020
rect 15838 14968 15844 15020
rect 15896 14968 15902 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16960 15017 16988 15116
rect 17494 15104 17500 15156
rect 17552 15144 17558 15156
rect 17681 15147 17739 15153
rect 17681 15144 17693 15147
rect 17552 15116 17693 15144
rect 17552 15104 17558 15116
rect 17681 15113 17693 15116
rect 17727 15113 17739 15147
rect 17681 15107 17739 15113
rect 18693 15147 18751 15153
rect 18693 15113 18705 15147
rect 18739 15144 18751 15147
rect 19242 15144 19248 15156
rect 18739 15116 19248 15144
rect 18739 15113 18751 15116
rect 18693 15107 18751 15113
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 19426 15104 19432 15156
rect 19484 15104 19490 15156
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 19576 15116 20024 15144
rect 19576 15104 19582 15116
rect 19444 15076 19472 15104
rect 19996 15085 20024 15116
rect 20070 15104 20076 15156
rect 20128 15104 20134 15156
rect 22005 15147 22063 15153
rect 22005 15113 22017 15147
rect 22051 15113 22063 15147
rect 22005 15107 22063 15113
rect 18524 15048 19472 15076
rect 19981 15079 20039 15085
rect 18524 15017 18552 15048
rect 19981 15045 19993 15079
rect 20027 15045 20039 15079
rect 19981 15039 20039 15045
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16632 14980 16681 15008
rect 16632 14968 16638 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 18509 15011 18567 15017
rect 18509 14977 18521 15011
rect 18555 14977 18567 15011
rect 18509 14971 18567 14977
rect 18966 14968 18972 15020
rect 19024 14968 19030 15020
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 15006 19211 15011
rect 20088 15008 20116 15104
rect 20622 15076 20628 15088
rect 20272 15048 20628 15076
rect 20272 15017 20300 15048
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 22020 15076 22048 15107
rect 23474 15104 23480 15156
rect 23532 15104 23538 15156
rect 23750 15104 23756 15156
rect 23808 15104 23814 15156
rect 24397 15147 24455 15153
rect 24397 15113 24409 15147
rect 24443 15144 24455 15147
rect 24486 15144 24492 15156
rect 24443 15116 24492 15144
rect 24443 15113 24455 15116
rect 24397 15107 24455 15113
rect 24486 15104 24492 15116
rect 24544 15104 24550 15156
rect 27617 15147 27675 15153
rect 27617 15144 27629 15147
rect 24596 15116 26188 15144
rect 22342 15079 22400 15085
rect 22342 15076 22354 15079
rect 22020 15048 22354 15076
rect 22342 15045 22354 15048
rect 22388 15045 22400 15079
rect 24596 15076 24624 15116
rect 26160 15088 26188 15116
rect 26804 15116 27629 15144
rect 26804 15088 26832 15116
rect 27617 15113 27629 15116
rect 27663 15113 27675 15147
rect 27617 15107 27675 15113
rect 29457 15147 29515 15153
rect 29457 15113 29469 15147
rect 29503 15144 29515 15147
rect 30006 15144 30012 15156
rect 29503 15116 30012 15144
rect 29503 15113 29515 15116
rect 29457 15107 29515 15113
rect 30006 15104 30012 15116
rect 30064 15104 30070 15156
rect 30926 15104 30932 15156
rect 30984 15104 30990 15156
rect 31849 15147 31907 15153
rect 31849 15113 31861 15147
rect 31895 15144 31907 15147
rect 33778 15144 33784 15156
rect 31895 15116 33784 15144
rect 31895 15113 31907 15116
rect 31849 15107 31907 15113
rect 33778 15104 33784 15116
rect 33836 15104 33842 15156
rect 35342 15104 35348 15156
rect 35400 15104 35406 15156
rect 36446 15104 36452 15156
rect 36504 15104 36510 15156
rect 37090 15104 37096 15156
rect 37148 15104 37154 15156
rect 22342 15039 22400 15045
rect 24228 15048 24624 15076
rect 19336 15006 20116 15008
rect 19199 14980 20116 15006
rect 20257 15011 20315 15017
rect 19199 14978 19364 14980
rect 19199 14977 19211 14978
rect 19153 14971 19211 14977
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20438 14968 20444 15020
rect 20496 14968 20502 15020
rect 20530 14968 20536 15020
rect 20588 14968 20594 15020
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 15008 20775 15011
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 20763 14980 21833 15008
rect 20763 14977 20775 14980
rect 20717 14971 20775 14977
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 22094 14968 22100 15020
rect 22152 14968 22158 15020
rect 23566 14968 23572 15020
rect 23624 15008 23630 15020
rect 23694 15011 23752 15017
rect 23694 15008 23706 15011
rect 23624 14980 23706 15008
rect 23624 14968 23630 14980
rect 23694 14977 23706 14980
rect 23740 14977 23752 15011
rect 23694 14971 23752 14977
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 24228 15017 24256 15048
rect 25038 15036 25044 15088
rect 25096 15076 25102 15088
rect 25133 15079 25191 15085
rect 25133 15076 25145 15079
rect 25096 15048 25145 15076
rect 25096 15036 25102 15048
rect 25133 15045 25145 15048
rect 25179 15045 25191 15079
rect 25133 15039 25191 15045
rect 26142 15036 26148 15088
rect 26200 15036 26206 15088
rect 26786 15036 26792 15088
rect 26844 15036 26850 15088
rect 27801 15079 27859 15085
rect 27801 15045 27813 15079
rect 27847 15076 27859 15079
rect 29546 15076 29552 15088
rect 27847 15048 29552 15076
rect 27847 15045 27859 15048
rect 27801 15039 27859 15045
rect 29546 15036 29552 15048
rect 29604 15036 29610 15088
rect 30024 15076 30052 15104
rect 30469 15079 30527 15085
rect 30469 15076 30481 15079
rect 30024 15048 30481 15076
rect 30469 15045 30481 15048
rect 30515 15045 30527 15079
rect 30469 15039 30527 15045
rect 30674 15079 30732 15085
rect 30674 15045 30686 15079
rect 30720 15076 30732 15079
rect 30720 15048 30788 15076
rect 30720 15045 30732 15048
rect 30674 15039 30732 15045
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 24305 15011 24363 15017
rect 24305 14977 24317 15011
rect 24351 14977 24363 15011
rect 24305 14971 24363 14977
rect 15657 14943 15715 14949
rect 15028 14912 15608 14940
rect 12176 14844 12296 14872
rect 11977 14835 12035 14841
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 11054 14804 11060 14816
rect 9907 14776 11060 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 11793 14807 11851 14813
rect 11793 14773 11805 14807
rect 11839 14804 11851 14807
rect 12158 14804 12164 14816
rect 11839 14776 12164 14804
rect 11839 14773 11851 14776
rect 11793 14767 11851 14773
rect 12158 14764 12164 14776
rect 12216 14764 12222 14816
rect 12268 14813 12296 14844
rect 12434 14832 12440 14884
rect 12492 14832 12498 14884
rect 12621 14875 12679 14881
rect 12621 14841 12633 14875
rect 12667 14872 12679 14875
rect 12989 14875 13047 14881
rect 12989 14872 13001 14875
rect 12667 14844 13001 14872
rect 12667 14841 12679 14844
rect 12621 14835 12679 14841
rect 12989 14841 13001 14844
rect 13035 14841 13047 14875
rect 12989 14835 13047 14841
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14773 12311 14807
rect 12452 14804 12480 14832
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12452 14776 12909 14804
rect 12253 14767 12311 14773
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 13464 14804 13492 14903
rect 13648 14872 13676 14903
rect 14660 14872 14688 14912
rect 13648 14844 14688 14872
rect 14734 14832 14740 14884
rect 14792 14832 14798 14884
rect 15286 14872 15292 14884
rect 15028 14844 15292 14872
rect 13136 14776 13492 14804
rect 14369 14807 14427 14813
rect 13136 14764 13142 14776
rect 14369 14773 14381 14807
rect 14415 14804 14427 14807
rect 15028 14804 15056 14844
rect 15286 14832 15292 14844
rect 15344 14832 15350 14884
rect 14415 14776 15056 14804
rect 15105 14807 15163 14813
rect 14415 14773 14427 14776
rect 14369 14767 14427 14773
rect 15105 14773 15117 14807
rect 15151 14804 15163 14807
rect 15194 14804 15200 14816
rect 15151 14776 15200 14804
rect 15151 14773 15163 14776
rect 15105 14767 15163 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 15580 14804 15608 14912
rect 15657 14909 15669 14943
rect 15703 14909 15715 14943
rect 15657 14903 15715 14909
rect 15672 14872 15700 14903
rect 17034 14900 17040 14952
rect 17092 14900 17098 14952
rect 18782 14900 18788 14952
rect 18840 14900 18846 14952
rect 19245 14943 19303 14949
rect 19245 14909 19257 14943
rect 19291 14909 19303 14943
rect 20548 14940 20576 14968
rect 19245 14903 19303 14909
rect 20088 14912 20576 14940
rect 21453 14943 21511 14949
rect 16669 14875 16727 14881
rect 16669 14872 16681 14875
rect 15672 14844 16681 14872
rect 16669 14841 16681 14844
rect 16715 14841 16727 14875
rect 16669 14835 16727 14841
rect 18966 14832 18972 14884
rect 19024 14832 19030 14884
rect 19150 14832 19156 14884
rect 19208 14872 19214 14884
rect 19260 14872 19288 14903
rect 20088 14872 20116 14912
rect 21453 14909 21465 14943
rect 21499 14940 21511 14943
rect 21634 14940 21640 14952
rect 21499 14912 21640 14940
rect 21499 14909 21511 14912
rect 21453 14903 21511 14909
rect 21634 14900 21640 14912
rect 21692 14900 21698 14952
rect 24320 14940 24348 14971
rect 24486 14968 24492 15020
rect 24544 14968 24550 15020
rect 24762 14968 24768 15020
rect 24820 15008 24826 15020
rect 25498 15008 25504 15020
rect 24820 14980 25504 15008
rect 24820 14968 24826 14980
rect 25498 14968 25504 14980
rect 25556 15008 25562 15020
rect 27062 15008 27068 15020
rect 25556 14980 27068 15008
rect 25556 14968 25562 14980
rect 27062 14968 27068 14980
rect 27120 15008 27126 15020
rect 27249 15011 27307 15017
rect 27249 15008 27261 15011
rect 27120 14980 27261 15008
rect 27120 14968 27126 14980
rect 27249 14977 27261 14980
rect 27295 14977 27307 15011
rect 27249 14971 27307 14977
rect 27522 14968 27528 15020
rect 27580 14968 27586 15020
rect 27614 14968 27620 15020
rect 27672 14968 27678 15020
rect 27982 14968 27988 15020
rect 28040 15008 28046 15020
rect 28077 15011 28135 15017
rect 28077 15008 28089 15011
rect 28040 14980 28089 15008
rect 28040 14968 28046 14980
rect 28077 14977 28089 14980
rect 28123 14977 28135 15011
rect 28077 14971 28135 14977
rect 28166 14968 28172 15020
rect 28224 15008 28230 15020
rect 28333 15011 28391 15017
rect 28333 15008 28345 15011
rect 28224 14980 28345 15008
rect 28224 14968 28230 14980
rect 28333 14977 28345 14980
rect 28379 14977 28391 15011
rect 28333 14971 28391 14977
rect 23584 14912 24348 14940
rect 25041 14943 25099 14949
rect 23584 14881 23612 14912
rect 25041 14909 25053 14943
rect 25087 14940 25099 14943
rect 25406 14940 25412 14952
rect 25087 14912 25412 14940
rect 25087 14909 25099 14912
rect 25041 14903 25099 14909
rect 25406 14900 25412 14912
rect 25464 14900 25470 14952
rect 25685 14943 25743 14949
rect 25685 14909 25697 14943
rect 25731 14909 25743 14943
rect 25685 14903 25743 14909
rect 19208 14844 19288 14872
rect 19812 14844 20116 14872
rect 20165 14875 20223 14881
rect 19208 14832 19214 14844
rect 18874 14804 18880 14816
rect 15580 14776 18880 14804
rect 18874 14764 18880 14776
rect 18932 14764 18938 14816
rect 18984 14804 19012 14832
rect 19812 14804 19840 14844
rect 20165 14841 20177 14875
rect 20211 14872 20223 14875
rect 20809 14875 20867 14881
rect 20809 14872 20821 14875
rect 20211 14844 20821 14872
rect 20211 14841 20223 14844
rect 20165 14835 20223 14841
rect 20809 14841 20821 14844
rect 20855 14841 20867 14875
rect 20809 14835 20867 14841
rect 23569 14875 23627 14881
rect 23569 14841 23581 14875
rect 23615 14841 23627 14875
rect 23569 14835 23627 14841
rect 24578 14832 24584 14884
rect 24636 14832 24642 14884
rect 24949 14875 25007 14881
rect 24949 14841 24961 14875
rect 24995 14872 25007 14875
rect 25590 14872 25596 14884
rect 24995 14844 25596 14872
rect 24995 14841 25007 14844
rect 24949 14835 25007 14841
rect 25590 14832 25596 14844
rect 25648 14832 25654 14884
rect 18984 14776 19840 14804
rect 19889 14807 19947 14813
rect 19889 14773 19901 14807
rect 19935 14804 19947 14807
rect 19978 14804 19984 14816
rect 19935 14776 19984 14804
rect 19935 14773 19947 14776
rect 19889 14767 19947 14773
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 20070 14764 20076 14816
rect 20128 14764 20134 14816
rect 25406 14764 25412 14816
rect 25464 14804 25470 14816
rect 25700 14804 25728 14903
rect 26326 14900 26332 14952
rect 26384 14940 26390 14952
rect 26697 14943 26755 14949
rect 26697 14940 26709 14943
rect 26384 14912 26709 14940
rect 26384 14900 26390 14912
rect 26697 14909 26709 14912
rect 26743 14909 26755 14943
rect 26697 14903 26755 14909
rect 26973 14943 27031 14949
rect 26973 14909 26985 14943
rect 27019 14940 27031 14943
rect 27632 14940 27660 14968
rect 30760 14952 30788 15048
rect 30944 15017 30972 15104
rect 31021 15079 31079 15085
rect 31021 15045 31033 15079
rect 31067 15076 31079 15079
rect 31754 15076 31760 15088
rect 31067 15048 31248 15076
rect 31067 15045 31079 15048
rect 31021 15039 31079 15045
rect 31220 15017 31248 15048
rect 31404 15048 31760 15076
rect 31404 15017 31432 15048
rect 31754 15036 31760 15048
rect 31812 15036 31818 15088
rect 33226 15036 33232 15088
rect 33284 15085 33290 15088
rect 33284 15076 33296 15085
rect 34330 15076 34336 15088
rect 33284 15048 33329 15076
rect 33520 15048 34336 15076
rect 33284 15039 33296 15048
rect 33284 15036 33290 15039
rect 30929 15011 30987 15017
rect 30929 14977 30941 15011
rect 30975 14977 30987 15011
rect 30929 14971 30987 14977
rect 31113 15011 31171 15017
rect 31113 14977 31125 15011
rect 31159 14977 31171 15011
rect 31113 14971 31171 14977
rect 31205 15011 31263 15017
rect 31205 14977 31217 15011
rect 31251 14977 31263 15011
rect 31205 14971 31263 14977
rect 31389 15011 31447 15017
rect 31389 14977 31401 15011
rect 31435 14977 31447 15011
rect 31389 14971 31447 14977
rect 31481 15011 31539 15017
rect 31481 14977 31493 15011
rect 31527 14977 31539 15011
rect 31481 14971 31539 14977
rect 31573 15011 31631 15017
rect 31573 14977 31585 15011
rect 31619 15008 31631 15011
rect 31619 14980 31754 15008
rect 31619 14977 31631 14980
rect 31573 14971 31631 14977
rect 27019 14912 27660 14940
rect 27019 14909 27031 14912
rect 26973 14903 27031 14909
rect 30742 14900 30748 14952
rect 30800 14940 30806 14952
rect 31128 14940 31156 14971
rect 30800 14912 31156 14940
rect 30800 14900 30806 14912
rect 31294 14900 31300 14952
rect 31352 14940 31358 14952
rect 31496 14940 31524 14971
rect 31352 14912 31524 14940
rect 31352 14900 31358 14912
rect 25774 14832 25780 14884
rect 25832 14872 25838 14884
rect 26145 14875 26203 14881
rect 26145 14872 26157 14875
rect 25832 14844 26157 14872
rect 25832 14832 25838 14844
rect 26145 14841 26157 14844
rect 26191 14841 26203 14875
rect 26145 14835 26203 14841
rect 25464 14776 25728 14804
rect 25464 14764 25470 14776
rect 25866 14764 25872 14816
rect 25924 14804 25930 14816
rect 26510 14804 26516 14816
rect 25924 14776 26516 14804
rect 25924 14764 25930 14776
rect 26510 14764 26516 14776
rect 26568 14804 26574 14816
rect 27065 14807 27123 14813
rect 27065 14804 27077 14807
rect 26568 14776 27077 14804
rect 26568 14764 26574 14776
rect 27065 14773 27077 14776
rect 27111 14773 27123 14807
rect 27065 14767 27123 14773
rect 27430 14764 27436 14816
rect 27488 14764 27494 14816
rect 27798 14764 27804 14816
rect 27856 14764 27862 14816
rect 30650 14764 30656 14816
rect 30708 14764 30714 14816
rect 30834 14764 30840 14816
rect 30892 14764 30898 14816
rect 31726 14804 31754 14980
rect 33410 14968 33416 15020
rect 33468 15008 33474 15020
rect 33520 15017 33548 15048
rect 34330 15036 34336 15048
rect 34388 15036 34394 15088
rect 36464 15076 36492 15104
rect 35544 15048 36492 15076
rect 33505 15011 33563 15017
rect 33505 15008 33517 15011
rect 33468 14980 33517 15008
rect 33468 14968 33474 14980
rect 33505 14977 33517 14980
rect 33551 14977 33563 15011
rect 33505 14971 33563 14977
rect 33594 14968 33600 15020
rect 33652 14968 33658 15020
rect 35544 15017 35572 15048
rect 35529 15011 35587 15017
rect 35529 14977 35541 15011
rect 35575 14977 35587 15011
rect 35529 14971 35587 14977
rect 35621 15011 35679 15017
rect 35621 14977 35633 15011
rect 35667 14977 35679 15011
rect 35621 14971 35679 14977
rect 32125 14807 32183 14813
rect 32125 14804 32137 14807
rect 31726 14776 32137 14804
rect 32125 14773 32137 14776
rect 32171 14804 32183 14807
rect 32582 14804 32588 14816
rect 32171 14776 32588 14804
rect 32171 14773 32183 14776
rect 32125 14767 32183 14773
rect 32582 14764 32588 14776
rect 32640 14764 32646 14816
rect 35636 14804 35664 14971
rect 35710 14968 35716 15020
rect 35768 15008 35774 15020
rect 35805 15011 35863 15017
rect 35805 15008 35817 15011
rect 35768 14980 35817 15008
rect 35768 14968 35774 14980
rect 35805 14977 35817 14980
rect 35851 14977 35863 15011
rect 35805 14971 35863 14977
rect 35897 15011 35955 15017
rect 35897 14977 35909 15011
rect 35943 15008 35955 15011
rect 37108 15008 37136 15104
rect 35943 14980 37136 15008
rect 35943 14977 35955 14980
rect 35897 14971 35955 14977
rect 35820 14940 35848 14971
rect 67634 14940 67640 14952
rect 35820 14912 41414 14940
rect 41386 14872 41414 14912
rect 45526 14912 67640 14940
rect 45526 14872 45554 14912
rect 67634 14900 67640 14912
rect 67692 14900 67698 14952
rect 41386 14844 45554 14872
rect 37274 14804 37280 14816
rect 35636 14776 37280 14804
rect 37274 14764 37280 14776
rect 37332 14764 37338 14816
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 11422 14600 11428 14612
rect 10928 14572 11428 14600
rect 10928 14560 10934 14572
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 12124 14572 13277 14600
rect 12124 14560 12130 14572
rect 13265 14569 13277 14572
rect 13311 14569 13323 14603
rect 13265 14563 13323 14569
rect 14734 14560 14740 14612
rect 14792 14600 14798 14612
rect 15654 14600 15660 14612
rect 14792 14572 15660 14600
rect 14792 14560 14798 14572
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 15838 14560 15844 14612
rect 15896 14600 15902 14612
rect 15933 14603 15991 14609
rect 15933 14600 15945 14603
rect 15896 14572 15945 14600
rect 15896 14560 15902 14572
rect 15933 14569 15945 14572
rect 15979 14569 15991 14603
rect 15933 14563 15991 14569
rect 16669 14603 16727 14609
rect 16669 14569 16681 14603
rect 16715 14600 16727 14603
rect 17034 14600 17040 14612
rect 16715 14572 17040 14600
rect 16715 14569 16727 14572
rect 16669 14563 16727 14569
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 19208 14572 19257 14600
rect 19208 14560 19214 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 20070 14600 20076 14612
rect 19245 14563 19303 14569
rect 19352 14572 20076 14600
rect 11054 14532 11060 14544
rect 10060 14504 11060 14532
rect 10060 14473 10088 14504
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14433 10103 14467
rect 11440 14464 11468 14560
rect 12158 14492 12164 14544
rect 12216 14532 12222 14544
rect 12805 14535 12863 14541
rect 12805 14532 12817 14535
rect 12216 14504 12817 14532
rect 12216 14492 12222 14504
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 10045 14427 10103 14433
rect 10152 14436 10732 14464
rect 11440 14436 11529 14464
rect 10152 14408 10180 14436
rect 9122 14356 9128 14408
rect 9180 14356 9186 14408
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14396 9459 14399
rect 9490 14396 9496 14408
rect 9447 14368 9496 14396
rect 9447 14365 9459 14368
rect 9401 14359 9459 14365
rect 9490 14356 9496 14368
rect 9548 14356 9554 14408
rect 10134 14356 10140 14408
rect 10192 14356 10198 14408
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 10704 14405 10732 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 12066 14424 12072 14476
rect 12124 14424 12130 14476
rect 11348 14405 11468 14406
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 11333 14399 11468 14405
rect 11333 14365 11345 14399
rect 11379 14396 11468 14399
rect 11882 14396 11888 14408
rect 11379 14378 11888 14396
rect 11379 14365 11391 14378
rect 11440 14368 11888 14378
rect 11333 14359 11391 14365
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12452 14405 12480 14504
rect 12805 14501 12817 14504
rect 12851 14501 12863 14535
rect 12805 14495 12863 14501
rect 18506 14492 18512 14544
rect 18564 14532 18570 14544
rect 19352 14532 19380 14572
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 21177 14603 21235 14609
rect 21177 14569 21189 14603
rect 21223 14600 21235 14603
rect 21634 14600 21640 14612
rect 21223 14572 21640 14600
rect 21223 14569 21235 14572
rect 21177 14563 21235 14569
rect 18564 14504 19380 14532
rect 18564 14492 18570 14504
rect 19426 14492 19432 14544
rect 19484 14532 19490 14544
rect 19521 14535 19579 14541
rect 19521 14532 19533 14535
rect 19484 14504 19533 14532
rect 19484 14492 19490 14504
rect 19521 14501 19533 14504
rect 19567 14501 19579 14535
rect 19521 14495 19579 14501
rect 19613 14535 19671 14541
rect 19613 14501 19625 14535
rect 19659 14532 19671 14535
rect 21192 14532 21220 14563
rect 21634 14560 21640 14572
rect 21692 14560 21698 14612
rect 24486 14560 24492 14612
rect 24544 14600 24550 14612
rect 25130 14600 25136 14612
rect 24544 14572 25136 14600
rect 24544 14560 24550 14572
rect 25130 14560 25136 14572
rect 25188 14600 25194 14612
rect 25682 14600 25688 14612
rect 25188 14572 25688 14600
rect 25188 14560 25194 14572
rect 25682 14560 25688 14572
rect 25740 14560 25746 14612
rect 26050 14560 26056 14612
rect 26108 14600 26114 14612
rect 26108 14572 27108 14600
rect 26108 14560 26114 14572
rect 19659 14504 21220 14532
rect 19659 14501 19671 14504
rect 19613 14495 19671 14501
rect 14185 14467 14243 14473
rect 14185 14464 14197 14467
rect 12544 14436 14197 14464
rect 12544 14405 12572 14436
rect 14185 14433 14197 14436
rect 14231 14433 14243 14467
rect 14185 14427 14243 14433
rect 16850 14424 16856 14476
rect 16908 14424 16914 14476
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17402 14464 17408 14476
rect 17175 14436 17408 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 18782 14424 18788 14476
rect 18840 14424 18846 14476
rect 19628 14464 19656 14495
rect 19306 14436 19656 14464
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14365 12403 14399
rect 12345 14359 12403 14365
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14365 12495 14399
rect 12437 14359 12495 14365
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14365 12587 14399
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 12529 14359 12587 14365
rect 13004 14368 13829 14396
rect 9508 14328 9536 14356
rect 10229 14331 10287 14337
rect 10229 14328 10241 14331
rect 9508 14300 10241 14328
rect 10229 14297 10241 14300
rect 10275 14297 10287 14331
rect 10428 14328 10456 14356
rect 11974 14328 11980 14340
rect 10428 14300 11980 14328
rect 10229 14291 10287 14297
rect 11974 14288 11980 14300
rect 12032 14328 12038 14340
rect 12227 14331 12285 14337
rect 12227 14328 12239 14331
rect 12032 14300 12239 14328
rect 12032 14288 12038 14300
rect 12227 14297 12239 14300
rect 12273 14297 12285 14331
rect 12227 14291 12285 14297
rect 8938 14220 8944 14272
rect 8996 14220 9002 14272
rect 9309 14263 9367 14269
rect 9309 14229 9321 14263
rect 9355 14260 9367 14263
rect 9493 14263 9551 14269
rect 9493 14260 9505 14263
rect 9355 14232 9505 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 9493 14229 9505 14232
rect 9539 14229 9551 14263
rect 9493 14223 9551 14229
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10643 14232 11161 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 11149 14229 11161 14232
rect 11195 14260 11207 14263
rect 11330 14260 11336 14272
rect 11195 14232 11336 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 11422 14220 11428 14272
rect 11480 14260 11486 14272
rect 12360 14260 12388 14359
rect 13004 14340 13032 14368
rect 13817 14365 13829 14368
rect 13863 14365 13875 14399
rect 13817 14359 13875 14365
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14365 14151 14399
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 14093 14359 14151 14365
rect 14200 14368 14289 14396
rect 12713 14331 12771 14337
rect 12713 14297 12725 14331
rect 12759 14328 12771 14331
rect 12894 14328 12900 14340
rect 12759 14300 12900 14328
rect 12759 14297 12771 14300
rect 12713 14291 12771 14297
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 12986 14288 12992 14340
rect 13044 14288 13050 14340
rect 13078 14288 13084 14340
rect 13136 14328 13142 14340
rect 13173 14331 13231 14337
rect 13173 14328 13185 14331
rect 13136 14300 13185 14328
rect 13136 14288 13142 14300
rect 13173 14297 13185 14300
rect 13219 14328 13231 14331
rect 14114 14328 14142 14359
rect 13219 14300 14142 14328
rect 13219 14297 13231 14300
rect 13173 14291 13231 14297
rect 11480 14232 12388 14260
rect 11480 14220 11486 14232
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 13004 14260 13032 14288
rect 14200 14272 14228 14368
rect 14277 14365 14289 14368
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14396 14611 14399
rect 15102 14396 15108 14408
rect 14599 14368 15108 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 15102 14356 15108 14368
rect 15160 14396 15166 14408
rect 15378 14396 15384 14408
rect 15160 14368 15384 14396
rect 15160 14356 15166 14368
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14396 17095 14399
rect 17310 14396 17316 14408
rect 17083 14368 17316 14396
rect 17083 14365 17095 14368
rect 17037 14359 17095 14365
rect 14820 14331 14878 14337
rect 14820 14297 14832 14331
rect 14866 14328 14878 14331
rect 14918 14328 14924 14340
rect 14866 14300 14924 14328
rect 14866 14297 14878 14300
rect 14820 14291 14878 14297
rect 14918 14288 14924 14300
rect 14976 14288 14982 14340
rect 16960 14328 16988 14359
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 18138 14356 18144 14408
rect 18196 14356 18202 14408
rect 18800 14396 18828 14424
rect 19306 14396 19334 14436
rect 20254 14424 20260 14476
rect 20312 14464 20318 14476
rect 20809 14467 20867 14473
rect 20809 14464 20821 14467
rect 20312 14436 20821 14464
rect 20312 14424 20318 14436
rect 20809 14433 20821 14436
rect 20855 14464 20867 14467
rect 23753 14467 23811 14473
rect 20855 14436 21404 14464
rect 20855 14433 20867 14436
rect 20809 14427 20867 14433
rect 18800 14368 19334 14396
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 19518 14396 19524 14408
rect 19475 14368 19524 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14396 19763 14399
rect 19751 14368 19840 14396
rect 19751 14365 19763 14368
rect 19705 14359 19763 14365
rect 16960 14300 19334 14328
rect 14182 14260 14188 14272
rect 12860 14232 14188 14260
rect 12860 14220 12866 14232
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 17586 14220 17592 14272
rect 17644 14220 17650 14272
rect 19306 14260 19334 14300
rect 19702 14260 19708 14272
rect 19306 14232 19708 14260
rect 19702 14220 19708 14232
rect 19760 14220 19766 14272
rect 19812 14260 19840 14368
rect 19886 14356 19892 14408
rect 19944 14356 19950 14408
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14396 20039 14399
rect 20070 14396 20076 14408
rect 20027 14368 20076 14396
rect 20027 14365 20039 14368
rect 19981 14359 20039 14365
rect 20070 14356 20076 14368
rect 20128 14396 20134 14408
rect 21376 14396 21404 14436
rect 23753 14433 23765 14467
rect 23799 14464 23811 14467
rect 24504 14464 24532 14560
rect 24578 14492 24584 14544
rect 24636 14492 24642 14544
rect 24946 14532 24952 14544
rect 24688 14504 24952 14532
rect 23799 14436 24532 14464
rect 23799 14433 23811 14436
rect 23753 14427 23811 14433
rect 22557 14399 22615 14405
rect 22557 14396 22569 14399
rect 20128 14368 21312 14396
rect 21376 14368 22569 14396
rect 20128 14356 20134 14368
rect 20438 14260 20444 14272
rect 19812 14232 20444 14260
rect 20438 14220 20444 14232
rect 20496 14220 20502 14272
rect 21284 14260 21312 14368
rect 22112 14340 22140 14368
rect 22557 14365 22569 14368
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 22738 14356 22744 14408
rect 22796 14356 22802 14408
rect 23014 14356 23020 14408
rect 23072 14396 23078 14408
rect 23477 14399 23535 14405
rect 23477 14396 23489 14399
rect 23072 14368 23489 14396
rect 23072 14356 23078 14368
rect 23477 14365 23489 14368
rect 23523 14365 23535 14399
rect 24596 14396 24624 14492
rect 24688 14473 24716 14504
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 24673 14467 24731 14473
rect 24673 14433 24685 14467
rect 24719 14433 24731 14467
rect 24673 14427 24731 14433
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 25317 14467 25375 14473
rect 25317 14464 25329 14467
rect 24912 14436 25329 14464
rect 24912 14424 24918 14436
rect 25317 14433 25329 14436
rect 25363 14433 25375 14467
rect 25317 14427 25375 14433
rect 26786 14424 26792 14476
rect 26844 14464 26850 14476
rect 26844 14436 27016 14464
rect 26844 14424 26850 14436
rect 24596 14368 24716 14396
rect 23477 14359 23535 14365
rect 22094 14288 22100 14340
rect 22152 14288 22158 14340
rect 22312 14331 22370 14337
rect 22312 14297 22324 14331
rect 22358 14328 22370 14331
rect 22756 14328 22784 14356
rect 22358 14300 22784 14328
rect 24688 14328 24716 14368
rect 24762 14356 24768 14408
rect 24820 14396 24826 14408
rect 26988 14405 27016 14436
rect 27080 14405 27108 14572
rect 27430 14560 27436 14612
rect 27488 14560 27494 14612
rect 27632 14572 30604 14600
rect 27249 14467 27307 14473
rect 27249 14433 27261 14467
rect 27295 14464 27307 14467
rect 27338 14464 27344 14476
rect 27295 14436 27344 14464
rect 27295 14433 27307 14436
rect 27249 14427 27307 14433
rect 27338 14424 27344 14436
rect 27396 14424 27402 14476
rect 27448 14464 27476 14560
rect 27632 14544 27660 14572
rect 27614 14492 27620 14544
rect 27672 14492 27678 14544
rect 28166 14492 28172 14544
rect 28224 14492 28230 14544
rect 27801 14467 27859 14473
rect 27801 14464 27813 14467
rect 27448 14436 27813 14464
rect 27801 14433 27813 14436
rect 27847 14433 27859 14467
rect 27801 14427 27859 14433
rect 27908 14436 29960 14464
rect 26973 14399 27031 14405
rect 24820 14368 26924 14396
rect 24820 14356 24826 14368
rect 25562 14331 25620 14337
rect 25562 14328 25574 14331
rect 24688 14300 25574 14328
rect 22358 14297 22370 14300
rect 22312 14291 22370 14297
rect 25562 14297 25574 14300
rect 25608 14297 25620 14331
rect 25562 14291 25620 14297
rect 25682 14288 25688 14340
rect 25740 14328 25746 14340
rect 26896 14328 26924 14368
rect 26973 14365 26985 14399
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 27065 14399 27123 14405
rect 27065 14365 27077 14399
rect 27111 14396 27123 14399
rect 27908 14396 27936 14436
rect 27111 14368 27936 14396
rect 27985 14399 28043 14405
rect 27111 14365 27123 14368
rect 27065 14359 27123 14365
rect 27985 14365 27997 14399
rect 28031 14398 28043 14399
rect 28169 14399 28227 14405
rect 28031 14370 28120 14398
rect 28031 14365 28043 14370
rect 27985 14359 28043 14365
rect 27614 14328 27620 14340
rect 25740 14300 26832 14328
rect 26896 14300 27620 14328
rect 25740 14288 25746 14300
rect 24670 14260 24676 14272
rect 21284 14232 24676 14260
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 25222 14220 25228 14272
rect 25280 14220 25286 14272
rect 26694 14220 26700 14272
rect 26752 14220 26758 14272
rect 26804 14260 26832 14300
rect 27614 14288 27620 14300
rect 27672 14288 27678 14340
rect 28092 14328 28120 14370
rect 28169 14365 28181 14399
rect 28215 14396 28227 14399
rect 28442 14396 28448 14408
rect 28215 14368 28448 14396
rect 28215 14365 28227 14368
rect 28169 14359 28227 14365
rect 28442 14356 28448 14368
rect 28500 14356 28506 14408
rect 28092 14300 29592 14328
rect 28092 14260 28120 14300
rect 29564 14272 29592 14300
rect 26804 14232 28120 14260
rect 29546 14220 29552 14272
rect 29604 14220 29610 14272
rect 29638 14220 29644 14272
rect 29696 14260 29702 14272
rect 29825 14263 29883 14269
rect 29825 14260 29837 14263
rect 29696 14232 29837 14260
rect 29696 14220 29702 14232
rect 29825 14229 29837 14232
rect 29871 14229 29883 14263
rect 29932 14260 29960 14436
rect 30009 14399 30067 14405
rect 30009 14365 30021 14399
rect 30055 14398 30067 14399
rect 30055 14396 30144 14398
rect 30374 14396 30380 14408
rect 30055 14370 30380 14396
rect 30055 14365 30067 14370
rect 30116 14368 30380 14370
rect 30009 14359 30067 14365
rect 30374 14356 30380 14368
rect 30432 14356 30438 14408
rect 30576 14328 30604 14572
rect 30834 14560 30840 14612
rect 30892 14560 30898 14612
rect 31757 14603 31815 14609
rect 31757 14569 31769 14603
rect 31803 14600 31815 14603
rect 35710 14600 35716 14612
rect 31803 14572 35716 14600
rect 31803 14569 31815 14572
rect 31757 14563 31815 14569
rect 35710 14560 35716 14572
rect 35768 14560 35774 14612
rect 30852 14396 30880 14560
rect 33594 14492 33600 14544
rect 33652 14492 33658 14544
rect 31573 14399 31631 14405
rect 31573 14396 31585 14399
rect 30852 14368 31585 14396
rect 31573 14365 31585 14368
rect 31619 14365 31631 14399
rect 32861 14399 32919 14405
rect 32861 14396 32873 14399
rect 31573 14359 31631 14365
rect 31726 14368 32873 14396
rect 31726 14328 31754 14368
rect 32861 14365 32873 14368
rect 32907 14396 32919 14399
rect 33612 14396 33640 14492
rect 32907 14368 33640 14396
rect 32907 14365 32919 14368
rect 32861 14359 32919 14365
rect 33778 14356 33784 14408
rect 33836 14396 33842 14408
rect 34517 14399 34575 14405
rect 34517 14396 34529 14399
rect 33836 14368 34529 14396
rect 33836 14356 33842 14368
rect 34517 14365 34529 14368
rect 34563 14396 34575 14399
rect 34563 14368 36124 14396
rect 34563 14365 34575 14368
rect 34517 14359 34575 14365
rect 30576 14300 31754 14328
rect 33502 14288 33508 14340
rect 33560 14328 33566 14340
rect 33689 14331 33747 14337
rect 33689 14328 33701 14331
rect 33560 14300 33701 14328
rect 33560 14288 33566 14300
rect 33689 14297 33701 14300
rect 33735 14328 33747 14331
rect 35342 14328 35348 14340
rect 33735 14300 35348 14328
rect 33735 14297 33747 14300
rect 33689 14291 33747 14297
rect 35342 14288 35348 14300
rect 35400 14288 35406 14340
rect 36096 14272 36124 14368
rect 31938 14260 31944 14272
rect 29932 14232 31944 14260
rect 29825 14223 29883 14229
rect 31938 14220 31944 14232
rect 31996 14220 32002 14272
rect 34330 14220 34336 14272
rect 34388 14260 34394 14272
rect 34425 14263 34483 14269
rect 34425 14260 34437 14263
rect 34388 14232 34437 14260
rect 34388 14220 34394 14232
rect 34425 14229 34437 14232
rect 34471 14229 34483 14263
rect 34425 14223 34483 14229
rect 36078 14220 36084 14272
rect 36136 14220 36142 14272
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 9122 14016 9128 14068
rect 9180 14016 9186 14068
rect 9309 14059 9367 14065
rect 9309 14025 9321 14059
rect 9355 14025 9367 14059
rect 9309 14019 9367 14025
rect 8110 13988 8116 14000
rect 7576 13960 8116 13988
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7576 13929 7604 13960
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 7561 13923 7619 13929
rect 7561 13920 7573 13923
rect 7064 13892 7573 13920
rect 7064 13880 7070 13892
rect 7561 13889 7573 13892
rect 7607 13889 7619 13923
rect 7561 13883 7619 13889
rect 9140 13852 9168 14016
rect 9324 13988 9352 14019
rect 10134 14016 10140 14068
rect 10192 14016 10198 14068
rect 10962 14016 10968 14068
rect 11020 14016 11026 14068
rect 11057 14059 11115 14065
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 12250 14056 12256 14068
rect 11103 14028 12256 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 10686 13997 10692 14000
rect 10668 13991 10692 13997
rect 9324 13960 10272 13988
rect 9950 13880 9956 13932
rect 10008 13918 10014 13932
rect 10244 13929 10272 13960
rect 10668 13957 10680 13991
rect 10668 13951 10692 13957
rect 10686 13948 10692 13951
rect 10744 13948 10750 14000
rect 10870 13948 10876 14000
rect 10928 13948 10934 14000
rect 10980 13929 11008 14016
rect 10045 13923 10103 13929
rect 10045 13918 10057 13923
rect 10008 13890 10057 13918
rect 10008 13880 10014 13890
rect 10045 13889 10057 13890
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10275 13892 10977 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 9140 13824 10548 13852
rect 8938 13744 8944 13796
rect 8996 13744 9002 13796
rect 10520 13793 10548 13824
rect 10505 13787 10563 13793
rect 10505 13753 10517 13787
rect 10551 13753 10563 13787
rect 10505 13747 10563 13753
rect 7824 13719 7882 13725
rect 7824 13685 7836 13719
rect 7870 13716 7882 13719
rect 8956 13716 8984 13744
rect 7870 13688 8984 13716
rect 10689 13719 10747 13725
rect 7870 13685 7882 13688
rect 7824 13679 7882 13685
rect 10689 13685 10701 13719
rect 10735 13716 10747 13719
rect 11072 13716 11100 14019
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12636 14028 15148 14056
rect 12636 13929 12664 14028
rect 15120 14000 15148 14028
rect 17586 14016 17592 14068
rect 17644 14016 17650 14068
rect 17687 14059 17745 14065
rect 17687 14025 17699 14059
rect 17733 14056 17745 14059
rect 18138 14056 18144 14068
rect 17733 14028 18144 14056
rect 17733 14025 17745 14028
rect 17687 14019 17745 14025
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 18877 14059 18935 14065
rect 18877 14025 18889 14059
rect 18923 14056 18935 14059
rect 18923 14028 19472 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 12894 13948 12900 14000
rect 12952 13948 12958 14000
rect 13906 13948 13912 14000
rect 13964 13948 13970 14000
rect 14918 13948 14924 14000
rect 14976 13948 14982 14000
rect 15102 13948 15108 14000
rect 15160 13948 15166 14000
rect 17604 13988 17632 14016
rect 17236 13960 17632 13988
rect 17773 13991 17831 13997
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 11882 13744 11888 13796
rect 11940 13784 11946 13796
rect 12636 13784 12664 13883
rect 14936 13852 14964 13948
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13920 15071 13923
rect 15059 13892 15148 13920
rect 15059 13889 15071 13892
rect 15013 13883 15071 13889
rect 15120 13852 15148 13892
rect 15194 13880 15200 13932
rect 15252 13880 15258 13932
rect 17236 13929 17264 13960
rect 17773 13957 17785 13991
rect 17819 13988 17831 13991
rect 17957 13991 18015 13997
rect 17957 13988 17969 13991
rect 17819 13960 17969 13988
rect 17819 13957 17831 13960
rect 17773 13951 17831 13957
rect 17957 13957 17969 13960
rect 18003 13957 18015 13991
rect 17957 13951 18015 13957
rect 18506 13948 18512 14000
rect 18564 13948 18570 14000
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13889 17095 13923
rect 17037 13883 17095 13889
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 17589 13923 17647 13929
rect 17589 13889 17601 13923
rect 17635 13920 17647 13923
rect 17678 13920 17684 13932
rect 17635 13892 17684 13920
rect 17635 13889 17647 13892
rect 17589 13883 17647 13889
rect 17052 13852 17080 13883
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 18230 13920 18236 13932
rect 17911 13892 18236 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 18230 13880 18236 13892
rect 18288 13920 18294 13932
rect 18524 13920 18552 13948
rect 19444 13932 19472 14028
rect 20622 14016 20628 14068
rect 20680 14016 20686 14068
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 21140 14028 21833 14056
rect 21140 14016 21146 14028
rect 21821 14025 21833 14028
rect 21867 14025 21879 14059
rect 23658 14056 23664 14068
rect 21821 14019 21879 14025
rect 22066 14028 23664 14056
rect 19978 13948 19984 14000
rect 20036 13997 20042 14000
rect 20036 13988 20048 13997
rect 20036 13960 20081 13988
rect 20036 13951 20048 13960
rect 20036 13948 20042 13951
rect 18288 13892 18552 13920
rect 18288 13880 18294 13892
rect 19426 13880 19432 13932
rect 19484 13880 19490 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 20640 13920 20668 14016
rect 20579 13892 20668 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 14936 13824 15056 13852
rect 15120 13824 17908 13852
rect 11940 13756 12664 13784
rect 11940 13744 11946 13756
rect 14182 13744 14188 13796
rect 14240 13784 14246 13796
rect 14369 13787 14427 13793
rect 14369 13784 14381 13787
rect 14240 13756 14381 13784
rect 14240 13744 14246 13756
rect 14369 13753 14381 13756
rect 14415 13753 14427 13787
rect 15028 13784 15056 13824
rect 15197 13787 15255 13793
rect 15197 13784 15209 13787
rect 15028 13756 15209 13784
rect 14369 13747 14427 13753
rect 15197 13753 15209 13756
rect 15243 13753 15255 13787
rect 15197 13747 15255 13753
rect 17880 13728 17908 13824
rect 18506 13812 18512 13864
rect 18564 13812 18570 13864
rect 20254 13812 20260 13864
rect 20312 13812 20318 13864
rect 20438 13812 20444 13864
rect 20496 13852 20502 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20496 13824 20637 13852
rect 20496 13812 20502 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 22066 13852 22094 14028
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 23753 14059 23811 14065
rect 23753 14025 23765 14059
rect 23799 14025 23811 14059
rect 23753 14019 23811 14025
rect 22189 13991 22247 13997
rect 22189 13957 22201 13991
rect 22235 13988 22247 13991
rect 23768 13988 23796 14019
rect 24854 14016 24860 14068
rect 24912 14016 24918 14068
rect 25225 14059 25283 14065
rect 25225 14025 25237 14059
rect 25271 14056 25283 14059
rect 25406 14056 25412 14068
rect 25271 14028 25412 14056
rect 25271 14025 25283 14028
rect 25225 14019 25283 14025
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 26237 14059 26295 14065
rect 26237 14025 26249 14059
rect 26283 14056 26295 14059
rect 26326 14056 26332 14068
rect 26283 14028 26332 14056
rect 26283 14025 26295 14028
rect 26237 14019 26295 14025
rect 26326 14016 26332 14028
rect 26384 14016 26390 14068
rect 29638 14056 29644 14068
rect 29472 14028 29644 14056
rect 24762 13988 24768 14000
rect 22235 13960 23704 13988
rect 23768 13960 24768 13988
rect 22235 13957 22247 13960
rect 22189 13951 22247 13957
rect 22281 13923 22339 13929
rect 22281 13889 22293 13923
rect 22327 13920 22339 13923
rect 23106 13920 23112 13932
rect 22327 13892 23112 13920
rect 22327 13889 22339 13892
rect 22281 13883 22339 13889
rect 23106 13880 23112 13892
rect 23164 13880 23170 13932
rect 23201 13923 23259 13929
rect 23201 13889 23213 13923
rect 23247 13889 23259 13923
rect 23676 13920 23704 13960
rect 24762 13948 24768 13960
rect 24820 13948 24826 14000
rect 24872 13988 24900 14016
rect 29472 13997 29500 14028
rect 29638 14016 29644 14028
rect 29696 14016 29702 14068
rect 33778 14056 33784 14068
rect 29840 14028 31984 14056
rect 29457 13991 29515 13997
rect 24872 13960 29224 13988
rect 24877 13923 24935 13929
rect 23676 13892 24164 13920
rect 23201 13883 23259 13889
rect 20625 13815 20683 13821
rect 20732 13824 22094 13852
rect 22373 13855 22431 13861
rect 10735 13688 11100 13716
rect 10735 13685 10747 13688
rect 10689 13679 10747 13685
rect 17218 13676 17224 13728
rect 17276 13676 17282 13728
rect 17862 13676 17868 13728
rect 17920 13716 17926 13728
rect 20732 13716 20760 13824
rect 22373 13821 22385 13855
rect 22419 13821 22431 13855
rect 22373 13815 22431 13821
rect 22388 13784 22416 13815
rect 23014 13812 23020 13864
rect 23072 13852 23078 13864
rect 23216 13852 23244 13883
rect 23072 13824 23244 13852
rect 23072 13812 23078 13824
rect 23474 13812 23480 13864
rect 23532 13812 23538 13864
rect 22462 13784 22468 13796
rect 22388 13756 22468 13784
rect 22462 13744 22468 13756
rect 22520 13744 22526 13796
rect 17920 13688 20760 13716
rect 24136 13716 24164 13892
rect 24877 13889 24889 13923
rect 24923 13920 24935 13923
rect 25038 13920 25044 13932
rect 24923 13892 25044 13920
rect 24923 13889 24935 13892
rect 24877 13883 24935 13889
rect 25038 13880 25044 13892
rect 25096 13880 25102 13932
rect 25148 13929 25176 13960
rect 26988 13932 27016 13960
rect 25133 13923 25191 13929
rect 25133 13889 25145 13923
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 25222 13880 25228 13932
rect 25280 13920 25286 13932
rect 25409 13923 25467 13929
rect 25409 13920 25421 13923
rect 25280 13892 25421 13920
rect 25280 13880 25286 13892
rect 25409 13889 25421 13892
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25498 13880 25504 13932
rect 25556 13920 25562 13932
rect 25685 13923 25743 13929
rect 25685 13920 25697 13923
rect 25556 13892 25697 13920
rect 25556 13880 25562 13892
rect 25685 13889 25697 13892
rect 25731 13889 25743 13923
rect 25685 13883 25743 13889
rect 25866 13880 25872 13932
rect 25924 13920 25930 13932
rect 26145 13923 26203 13929
rect 26145 13920 26157 13923
rect 25924 13892 26157 13920
rect 25924 13880 25930 13892
rect 26145 13889 26157 13892
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 26329 13923 26387 13929
rect 26329 13889 26341 13923
rect 26375 13920 26387 13923
rect 26418 13920 26424 13932
rect 26375 13892 26424 13920
rect 26375 13889 26387 13892
rect 26329 13883 26387 13889
rect 25593 13855 25651 13861
rect 25593 13821 25605 13855
rect 25639 13852 25651 13855
rect 25774 13852 25780 13864
rect 25639 13824 25780 13852
rect 25639 13821 25651 13824
rect 25593 13815 25651 13821
rect 25774 13812 25780 13824
rect 25832 13812 25838 13864
rect 26160 13852 26188 13883
rect 26418 13880 26424 13892
rect 26476 13880 26482 13932
rect 26694 13880 26700 13932
rect 26752 13880 26758 13932
rect 26970 13880 26976 13932
rect 27028 13880 27034 13932
rect 27246 13929 27252 13932
rect 27240 13920 27252 13929
rect 27207 13892 27252 13920
rect 27240 13883 27252 13892
rect 27246 13880 27252 13883
rect 27304 13880 27310 13932
rect 29196 13929 29224 13960
rect 29457 13957 29469 13991
rect 29503 13957 29515 13991
rect 29457 13951 29515 13957
rect 29546 13948 29552 14000
rect 29604 13988 29610 14000
rect 29840 13988 29868 14028
rect 31849 13991 31907 13997
rect 31849 13988 31861 13991
rect 29604 13960 29868 13988
rect 30682 13960 31861 13988
rect 29604 13948 29610 13960
rect 31849 13957 31861 13960
rect 31895 13957 31907 13991
rect 31849 13951 31907 13957
rect 31956 13988 31984 14028
rect 33060 14028 33784 14056
rect 33060 13988 33088 14028
rect 33778 14016 33784 14028
rect 33836 14016 33842 14068
rect 31956 13960 33088 13988
rect 31956 13929 31984 13960
rect 29181 13923 29239 13929
rect 29181 13889 29193 13923
rect 29227 13889 29239 13923
rect 29181 13883 29239 13889
rect 31941 13923 31999 13929
rect 31941 13889 31953 13923
rect 31987 13889 31999 13923
rect 31941 13883 31999 13889
rect 32582 13880 32588 13932
rect 32640 13880 32646 13932
rect 33060 13929 33088 13960
rect 34330 13948 34336 14000
rect 34388 13948 34394 14000
rect 33045 13923 33103 13929
rect 33045 13889 33057 13923
rect 33091 13889 33103 13923
rect 33045 13883 33103 13889
rect 35069 13923 35127 13929
rect 35069 13889 35081 13923
rect 35115 13920 35127 13923
rect 35115 13892 35388 13920
rect 35115 13889 35127 13892
rect 35069 13883 35127 13889
rect 35360 13864 35388 13892
rect 35434 13880 35440 13932
rect 35492 13920 35498 13932
rect 35989 13923 36047 13929
rect 35989 13920 36001 13923
rect 35492 13892 36001 13920
rect 35492 13880 35498 13892
rect 35989 13889 36001 13892
rect 36035 13889 36047 13923
rect 35989 13883 36047 13889
rect 36170 13880 36176 13932
rect 36228 13880 36234 13932
rect 26605 13855 26663 13861
rect 26605 13852 26617 13855
rect 26160 13824 26617 13852
rect 26605 13821 26617 13824
rect 26651 13821 26663 13855
rect 26605 13815 26663 13821
rect 30929 13855 30987 13861
rect 30929 13821 30941 13855
rect 30975 13852 30987 13855
rect 31202 13852 31208 13864
rect 30975 13824 31208 13852
rect 30975 13821 30987 13824
rect 30929 13815 30987 13821
rect 25501 13787 25559 13793
rect 25501 13753 25513 13787
rect 25547 13784 25559 13787
rect 25958 13784 25964 13796
rect 25547 13756 25964 13784
rect 25547 13753 25559 13756
rect 25501 13747 25559 13753
rect 25958 13744 25964 13756
rect 26016 13744 26022 13796
rect 30558 13744 30564 13796
rect 30616 13784 30622 13796
rect 30944 13784 30972 13815
rect 31202 13812 31208 13824
rect 31260 13852 31266 13864
rect 31573 13855 31631 13861
rect 31573 13852 31585 13855
rect 31260 13824 31585 13852
rect 31260 13812 31266 13824
rect 31573 13821 31585 13824
rect 31619 13821 31631 13855
rect 31573 13815 31631 13821
rect 32674 13812 32680 13864
rect 32732 13812 32738 13864
rect 34790 13812 34796 13864
rect 34848 13812 34854 13864
rect 35253 13855 35311 13861
rect 35253 13821 35265 13855
rect 35299 13821 35311 13855
rect 35253 13815 35311 13821
rect 30616 13756 30972 13784
rect 30616 13744 30622 13756
rect 26050 13716 26056 13728
rect 24136 13688 26056 13716
rect 17920 13676 17926 13688
rect 26050 13676 26056 13688
rect 26108 13676 26114 13728
rect 28350 13676 28356 13728
rect 28408 13676 28414 13728
rect 31018 13676 31024 13728
rect 31076 13676 31082 13728
rect 33134 13676 33140 13728
rect 33192 13676 33198 13728
rect 33321 13719 33379 13725
rect 33321 13685 33333 13719
rect 33367 13716 33379 13719
rect 34146 13716 34152 13728
rect 33367 13688 34152 13716
rect 33367 13685 33379 13688
rect 33321 13679 33379 13685
rect 34146 13676 34152 13688
rect 34204 13716 34210 13728
rect 35268 13716 35296 13815
rect 35342 13812 35348 13864
rect 35400 13812 35406 13864
rect 35897 13855 35955 13861
rect 35897 13821 35909 13855
rect 35943 13852 35955 13855
rect 36354 13852 36360 13864
rect 35943 13824 36360 13852
rect 35943 13821 35955 13824
rect 35897 13815 35955 13821
rect 36354 13812 36360 13824
rect 36412 13812 36418 13864
rect 34204 13688 35296 13716
rect 35989 13719 36047 13725
rect 34204 13676 34210 13688
rect 35989 13685 36001 13719
rect 36035 13716 36047 13719
rect 36262 13716 36268 13728
rect 36035 13688 36268 13716
rect 36035 13685 36047 13688
rect 35989 13679 36047 13685
rect 36262 13676 36268 13688
rect 36320 13676 36326 13728
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 8570 13472 8576 13524
rect 8628 13472 8634 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10686 13512 10692 13524
rect 10008 13484 10692 13512
rect 10008 13472 10014 13484
rect 10686 13472 10692 13484
rect 10744 13512 10750 13524
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 10744 13484 10885 13512
rect 10744 13472 10750 13484
rect 10873 13481 10885 13484
rect 10919 13481 10931 13515
rect 10873 13475 10931 13481
rect 12069 13515 12127 13521
rect 12069 13481 12081 13515
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 9968 13444 9996 13472
rect 9600 13416 9996 13444
rect 9600 13385 9628 13416
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11517 13447 11575 13453
rect 11517 13444 11529 13447
rect 11112 13416 11529 13444
rect 11112 13404 11118 13416
rect 11517 13413 11529 13416
rect 11563 13444 11575 13447
rect 11885 13447 11943 13453
rect 11885 13444 11897 13447
rect 11563 13416 11897 13444
rect 11563 13413 11575 13416
rect 11517 13407 11575 13413
rect 11885 13413 11897 13416
rect 11931 13413 11943 13447
rect 11885 13407 11943 13413
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13345 9643 13379
rect 9585 13339 9643 13345
rect 9692 13348 10548 13376
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 8662 13308 8668 13320
rect 8527 13280 8668 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 8662 13268 8668 13280
rect 8720 13308 8726 13320
rect 9692 13317 9720 13348
rect 9677 13311 9735 13317
rect 8720 13280 9628 13308
rect 8720 13268 8726 13280
rect 9600 13252 9628 13280
rect 9677 13277 9689 13311
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13308 10011 13311
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 9999 13280 10149 13308
rect 9999 13277 10011 13280
rect 9953 13271 10011 13277
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10410 13268 10416 13320
rect 10468 13268 10474 13320
rect 9582 13200 9588 13252
rect 9640 13200 9646 13252
rect 10045 13243 10103 13249
rect 10045 13209 10057 13243
rect 10091 13240 10103 13243
rect 10428 13240 10456 13268
rect 10091 13212 10456 13240
rect 10520 13240 10548 13348
rect 11330 13336 11336 13388
rect 11388 13376 11394 13388
rect 12084 13376 12112 13475
rect 12526 13472 12532 13524
rect 12584 13472 12590 13524
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13512 13875 13515
rect 13906 13512 13912 13524
rect 13863 13484 13912 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18506 13512 18512 13524
rect 18012 13484 18512 13512
rect 18012 13472 18018 13484
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 22465 13515 22523 13521
rect 22465 13481 22477 13515
rect 22511 13512 22523 13515
rect 22830 13512 22836 13524
rect 22511 13484 22836 13512
rect 22511 13481 22523 13484
rect 22465 13475 22523 13481
rect 22830 13472 22836 13484
rect 22888 13472 22894 13524
rect 30374 13472 30380 13524
rect 30432 13472 30438 13524
rect 30650 13472 30656 13524
rect 30708 13512 30714 13524
rect 30837 13515 30895 13521
rect 30837 13512 30849 13515
rect 30708 13484 30849 13512
rect 30708 13472 30714 13484
rect 30837 13481 30849 13484
rect 30883 13481 30895 13515
rect 30837 13475 30895 13481
rect 31018 13472 31024 13524
rect 31076 13472 31082 13524
rect 33965 13515 34023 13521
rect 33965 13481 33977 13515
rect 34011 13512 34023 13515
rect 34333 13515 34391 13521
rect 34333 13512 34345 13515
rect 34011 13484 34345 13512
rect 34011 13481 34023 13484
rect 33965 13475 34023 13481
rect 34333 13481 34345 13484
rect 34379 13512 34391 13515
rect 34422 13512 34428 13524
rect 34379 13484 34428 13512
rect 34379 13481 34391 13484
rect 34333 13475 34391 13481
rect 34422 13472 34428 13484
rect 34480 13472 34486 13524
rect 34701 13515 34759 13521
rect 34701 13481 34713 13515
rect 34747 13512 34759 13515
rect 34790 13512 34796 13524
rect 34747 13484 34796 13512
rect 34747 13481 34759 13484
rect 34701 13475 34759 13481
rect 34790 13472 34796 13484
rect 34848 13472 34854 13524
rect 35434 13472 35440 13524
rect 35492 13472 35498 13524
rect 12158 13404 12164 13456
rect 12216 13444 12222 13456
rect 13078 13444 13084 13456
rect 12216 13416 13084 13444
rect 12216 13404 12222 13416
rect 12802 13376 12808 13388
rect 11388 13348 11744 13376
rect 12084 13348 12808 13376
rect 11388 13336 11394 13348
rect 11716 13320 11744 13348
rect 12802 13336 12808 13348
rect 12860 13376 12866 13388
rect 12860 13348 12940 13376
rect 12860 13336 12866 13348
rect 10686 13268 10692 13320
rect 10744 13268 10750 13320
rect 11054 13268 11060 13320
rect 11112 13268 11118 13320
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11609 13311 11667 13317
rect 11609 13308 11621 13311
rect 11296 13307 11376 13308
rect 11532 13307 11621 13308
rect 11296 13280 11621 13307
rect 11296 13268 11302 13280
rect 11348 13279 11560 13280
rect 11333 13243 11391 13249
rect 11333 13240 11345 13243
rect 10520 13212 11345 13240
rect 10091 13209 10103 13212
rect 10045 13203 10103 13209
rect 11333 13209 11345 13212
rect 11379 13209 11391 13243
rect 11333 13203 11391 13209
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9401 13175 9459 13181
rect 9401 13172 9413 13175
rect 8996 13144 9413 13172
rect 8996 13132 9002 13144
rect 9401 13141 9413 13144
rect 9447 13141 9459 13175
rect 9401 13135 9459 13141
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 11440 13172 11468 13279
rect 11609 13277 11621 13280
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 11698 13268 11704 13320
rect 11756 13268 11762 13320
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 12912 13317 12940 13348
rect 13004 13317 13032 13416
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 29086 13404 29092 13456
rect 29144 13444 29150 13456
rect 30561 13447 30619 13453
rect 30561 13444 30573 13447
rect 29144 13416 30573 13444
rect 29144 13404 29150 13416
rect 30561 13413 30573 13416
rect 30607 13413 30619 13447
rect 31036 13444 31064 13472
rect 30561 13407 30619 13413
rect 30668 13416 31064 13444
rect 34517 13447 34575 13453
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 13872 13348 13952 13376
rect 13872 13336 13878 13348
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13277 12955 13311
rect 12897 13271 12955 13277
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 13630 13268 13636 13320
rect 13688 13268 13694 13320
rect 13924 13317 13952 13348
rect 15102 13336 15108 13388
rect 15160 13336 15166 13388
rect 20073 13379 20131 13385
rect 20073 13345 20085 13379
rect 20119 13376 20131 13379
rect 20254 13376 20260 13388
rect 20119 13348 20260 13376
rect 20119 13345 20131 13348
rect 20073 13339 20131 13345
rect 20254 13336 20260 13348
rect 20312 13336 20318 13388
rect 22462 13336 22468 13388
rect 22520 13376 22526 13388
rect 23017 13379 23075 13385
rect 23017 13376 23029 13379
rect 22520 13348 23029 13376
rect 22520 13336 22526 13348
rect 23017 13345 23029 13348
rect 23063 13376 23075 13379
rect 23750 13376 23756 13388
rect 23063 13348 23756 13376
rect 23063 13345 23075 13348
rect 23017 13339 23075 13345
rect 23750 13336 23756 13348
rect 23808 13336 23814 13388
rect 26970 13336 26976 13388
rect 27028 13336 27034 13388
rect 28350 13336 28356 13388
rect 28408 13376 28414 13388
rect 28721 13379 28779 13385
rect 28721 13376 28733 13379
rect 28408 13348 28733 13376
rect 28408 13336 28414 13348
rect 28721 13345 28733 13348
rect 28767 13345 28779 13379
rect 28721 13339 28779 13345
rect 29825 13379 29883 13385
rect 29825 13345 29837 13379
rect 29871 13376 29883 13379
rect 29871 13348 30604 13376
rect 29871 13345 29883 13348
rect 29825 13339 29883 13345
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13277 13967 13311
rect 15120 13308 15148 13336
rect 30576 13320 30604 13348
rect 30668 13327 30696 13416
rect 34517 13413 34529 13447
rect 34563 13444 34575 13447
rect 35452 13444 35480 13472
rect 36170 13444 36176 13456
rect 34563 13416 35480 13444
rect 35544 13416 36176 13444
rect 34563 13413 34575 13416
rect 34517 13407 34575 13413
rect 32217 13379 32275 13385
rect 32217 13345 32229 13379
rect 32263 13376 32275 13379
rect 33502 13376 33508 13388
rect 32263 13348 33508 13376
rect 32263 13345 32275 13348
rect 32217 13339 32275 13345
rect 33502 13336 33508 13348
rect 33560 13336 33566 13388
rect 30653 13321 30711 13327
rect 16577 13311 16635 13317
rect 16577 13308 16589 13311
rect 15120 13280 16589 13308
rect 13909 13271 13967 13277
rect 16577 13277 16589 13280
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 16844 13311 16902 13317
rect 16844 13277 16856 13311
rect 16890 13308 16902 13311
rect 17218 13308 17224 13320
rect 16890 13280 17224 13308
rect 16890 13277 16902 13280
rect 16844 13271 16902 13277
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 17862 13268 17868 13320
rect 17920 13308 17926 13320
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 17920 13280 18061 13308
rect 17920 13268 17926 13280
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 18230 13268 18236 13320
rect 18288 13268 18294 13320
rect 20438 13268 20444 13320
rect 20496 13268 20502 13320
rect 27614 13268 27620 13320
rect 27672 13308 27678 13320
rect 27801 13311 27859 13317
rect 27801 13308 27813 13311
rect 27672 13280 27813 13308
rect 27672 13268 27678 13280
rect 27801 13277 27813 13280
rect 27847 13277 27859 13311
rect 27801 13271 27859 13277
rect 29914 13268 29920 13320
rect 29972 13308 29978 13320
rect 30009 13311 30067 13317
rect 30009 13308 30021 13311
rect 29972 13280 30021 13308
rect 29972 13268 29978 13280
rect 30009 13277 30021 13280
rect 30055 13277 30067 13311
rect 30009 13271 30067 13277
rect 30469 13311 30527 13317
rect 30469 13277 30481 13311
rect 30515 13277 30527 13311
rect 30469 13271 30527 13277
rect 12253 13243 12311 13249
rect 12253 13209 12265 13243
rect 12299 13240 12311 13243
rect 12728 13240 12756 13268
rect 13648 13240 13676 13268
rect 15378 13249 15384 13252
rect 12299 13212 13676 13240
rect 12299 13209 12311 13212
rect 12253 13203 12311 13209
rect 15372 13203 15384 13249
rect 15378 13200 15384 13203
rect 15436 13200 15442 13252
rect 21450 13200 21456 13252
rect 21508 13200 21514 13252
rect 22925 13243 22983 13249
rect 22925 13240 22937 13243
rect 21882 13212 22937 13240
rect 21882 13184 21910 13212
rect 22925 13209 22937 13212
rect 22971 13209 22983 13243
rect 22925 13203 22983 13209
rect 30484 13240 30512 13271
rect 30558 13268 30564 13320
rect 30616 13268 30622 13320
rect 30653 13287 30665 13321
rect 30699 13287 30711 13321
rect 35544 13320 35572 13416
rect 36170 13404 36176 13416
rect 36228 13444 36234 13456
rect 36228 13416 36676 13444
rect 36228 13404 36234 13416
rect 36081 13379 36139 13385
rect 35636 13348 36032 13376
rect 30926 13308 30932 13320
rect 30653 13281 30711 13287
rect 30760 13280 30932 13308
rect 30760 13240 30788 13280
rect 30926 13268 30932 13280
rect 30984 13268 30990 13320
rect 35345 13311 35403 13317
rect 35345 13277 35357 13311
rect 35391 13308 35403 13311
rect 35437 13311 35495 13317
rect 35437 13308 35449 13311
rect 35391 13280 35449 13308
rect 35391 13277 35403 13280
rect 35345 13271 35403 13277
rect 35437 13277 35449 13280
rect 35483 13277 35495 13311
rect 35437 13271 35495 13277
rect 35526 13268 35532 13320
rect 35584 13268 35590 13320
rect 35636 13317 35664 13348
rect 35621 13311 35679 13317
rect 35621 13277 35633 13311
rect 35667 13277 35679 13311
rect 36004 13310 36032 13348
rect 36081 13345 36093 13379
rect 36127 13376 36139 13379
rect 36354 13376 36360 13388
rect 36127 13348 36360 13376
rect 36127 13345 36139 13348
rect 36081 13339 36139 13345
rect 36354 13336 36360 13348
rect 36412 13336 36418 13388
rect 36004 13308 36124 13310
rect 36262 13308 36268 13320
rect 36004 13282 36268 13308
rect 36096 13280 36268 13282
rect 35621 13271 35679 13277
rect 36262 13268 36268 13280
rect 36320 13308 36326 13320
rect 36648 13317 36676 13416
rect 36633 13311 36691 13317
rect 36320 13280 36400 13308
rect 36320 13268 36326 13280
rect 30484 13212 30788 13240
rect 10744 13144 11468 13172
rect 12053 13175 12111 13181
rect 10744 13132 10750 13144
rect 12053 13141 12065 13175
rect 12099 13172 12111 13175
rect 12158 13172 12164 13184
rect 12099 13144 12164 13172
rect 12099 13141 12111 13144
rect 12053 13135 12111 13141
rect 12158 13132 12164 13144
rect 12216 13132 12222 13184
rect 16485 13175 16543 13181
rect 16485 13141 16497 13175
rect 16531 13172 16543 13175
rect 16942 13172 16948 13184
rect 16531 13144 16948 13172
rect 16531 13141 16543 13144
rect 16485 13135 16543 13141
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 18141 13175 18199 13181
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 18230 13172 18236 13184
rect 18187 13144 18236 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 18230 13132 18236 13144
rect 18288 13132 18294 13184
rect 21818 13132 21824 13184
rect 21876 13181 21910 13184
rect 21876 13175 21925 13181
rect 21876 13141 21879 13175
rect 21913 13141 21925 13175
rect 21876 13135 21925 13141
rect 21876 13132 21882 13135
rect 22830 13132 22836 13184
rect 22888 13132 22894 13184
rect 28166 13132 28172 13184
rect 28224 13132 28230 13184
rect 29917 13175 29975 13181
rect 29917 13141 29929 13175
rect 29963 13172 29975 13175
rect 30098 13172 30104 13184
rect 29963 13144 30104 13172
rect 29963 13141 29975 13144
rect 29917 13135 29975 13141
rect 30098 13132 30104 13144
rect 30156 13172 30162 13184
rect 30484 13172 30512 13212
rect 32490 13200 32496 13252
rect 32548 13200 32554 13252
rect 33134 13200 33140 13252
rect 33192 13200 33198 13252
rect 34146 13200 34152 13252
rect 34204 13200 34210 13252
rect 34365 13243 34423 13249
rect 34365 13209 34377 13243
rect 34411 13240 34423 13243
rect 34606 13240 34612 13252
rect 34411 13212 34612 13240
rect 34411 13209 34423 13212
rect 34365 13203 34423 13209
rect 34606 13200 34612 13212
rect 34664 13240 34670 13252
rect 35713 13243 35771 13249
rect 34664 13212 34928 13240
rect 34664 13200 34670 13212
rect 30156 13144 30512 13172
rect 34900 13172 34928 13212
rect 35713 13209 35725 13243
rect 35759 13209 35771 13243
rect 35713 13203 35771 13209
rect 35728 13172 35756 13203
rect 35802 13200 35808 13252
rect 35860 13200 35866 13252
rect 35986 13249 35992 13252
rect 35943 13243 35992 13249
rect 35943 13209 35955 13243
rect 35989 13209 35992 13243
rect 35943 13203 35992 13209
rect 35986 13200 35992 13203
rect 36044 13240 36050 13252
rect 36044 13212 36124 13240
rect 36044 13200 36050 13212
rect 34900 13144 35756 13172
rect 36096 13172 36124 13212
rect 36170 13200 36176 13252
rect 36228 13200 36234 13252
rect 36372 13249 36400 13280
rect 36633 13277 36645 13311
rect 36679 13277 36691 13311
rect 36633 13271 36691 13277
rect 36817 13311 36875 13317
rect 36817 13277 36829 13311
rect 36863 13277 36875 13311
rect 36817 13271 36875 13277
rect 36357 13243 36415 13249
rect 36357 13209 36369 13243
rect 36403 13209 36415 13243
rect 36357 13203 36415 13209
rect 36832 13184 36860 13271
rect 36541 13175 36599 13181
rect 36541 13172 36553 13175
rect 36096 13144 36553 13172
rect 30156 13132 30162 13144
rect 36541 13141 36553 13144
rect 36587 13141 36599 13175
rect 36541 13135 36599 13141
rect 36722 13132 36728 13184
rect 36780 13132 36786 13184
rect 36814 13132 36820 13184
rect 36872 13132 36878 13184
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 11882 12968 11888 12980
rect 8404 12940 11888 12968
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8404 12841 8432 12940
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 12032 12940 12874 12968
rect 12032 12928 12038 12940
rect 8665 12903 8723 12909
rect 8665 12869 8677 12903
rect 8711 12900 8723 12903
rect 8938 12900 8944 12912
rect 8711 12872 8944 12900
rect 8711 12869 8723 12872
rect 8665 12863 8723 12869
rect 8938 12860 8944 12872
rect 8996 12860 9002 12912
rect 9674 12860 9680 12912
rect 9732 12860 9738 12912
rect 11054 12860 11060 12912
rect 11112 12860 11118 12912
rect 12846 12909 12874 12940
rect 17862 12928 17868 12980
rect 17920 12928 17926 12980
rect 18138 12968 18144 12980
rect 17972 12940 18144 12968
rect 11241 12903 11299 12909
rect 11241 12869 11253 12903
rect 11287 12900 11299 12903
rect 12621 12903 12679 12909
rect 12621 12900 12633 12903
rect 11287 12872 12633 12900
rect 11287 12869 11299 12872
rect 11241 12863 11299 12869
rect 12621 12869 12633 12872
rect 12667 12869 12679 12903
rect 12621 12863 12679 12869
rect 12831 12903 12889 12909
rect 12831 12869 12843 12903
rect 12877 12869 12889 12903
rect 12831 12863 12889 12869
rect 14829 12903 14887 12909
rect 14829 12869 14841 12903
rect 14875 12900 14887 12903
rect 15102 12900 15108 12912
rect 14875 12872 15108 12900
rect 14875 12869 14887 12872
rect 14829 12863 14887 12869
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 17681 12903 17739 12909
rect 17681 12869 17693 12903
rect 17727 12900 17739 12903
rect 17880 12900 17908 12928
rect 17727 12872 17908 12900
rect 17727 12869 17739 12872
rect 17681 12863 17739 12869
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8352 12804 8401 12832
rect 8352 12792 8358 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 11072 12832 11100 12860
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 11072 12804 11161 12832
rect 8389 12795 8447 12801
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 11756 12804 11897 12832
rect 11756 12792 11762 12804
rect 11885 12801 11897 12804
rect 11931 12832 11943 12835
rect 11931 12804 12296 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 10686 12764 10692 12776
rect 10183 12736 10692 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 12158 12724 12164 12776
rect 12216 12724 12222 12776
rect 12268 12764 12296 12804
rect 12526 12792 12532 12844
rect 12584 12792 12590 12844
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12801 12771 12835
rect 12713 12795 12771 12801
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12832 14059 12835
rect 15470 12832 15476 12844
rect 14047 12804 15476 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 12728 12764 12756 12795
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 16942 12792 16948 12844
rect 17000 12792 17006 12844
rect 17862 12792 17868 12844
rect 17920 12792 17926 12844
rect 17972 12841 18000 12940
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 20438 12928 20444 12980
rect 20496 12928 20502 12980
rect 20622 12928 20628 12980
rect 20680 12928 20686 12980
rect 20898 12928 20904 12980
rect 20956 12928 20962 12980
rect 21450 12928 21456 12980
rect 21508 12928 21514 12980
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 24581 12971 24639 12977
rect 24581 12968 24593 12971
rect 22888 12940 24593 12968
rect 22888 12928 22894 12940
rect 24581 12937 24593 12940
rect 24627 12937 24639 12971
rect 24581 12931 24639 12937
rect 24949 12971 25007 12977
rect 24949 12937 24961 12971
rect 24995 12968 25007 12971
rect 27295 12971 27353 12977
rect 27295 12968 27307 12971
rect 24995 12940 27307 12968
rect 24995 12937 25007 12940
rect 24949 12931 25007 12937
rect 27295 12937 27307 12940
rect 27341 12968 27353 12971
rect 27341 12940 29224 12968
rect 27341 12937 27353 12940
rect 27295 12931 27353 12937
rect 20254 12900 20260 12912
rect 18156 12872 20260 12900
rect 18156 12841 18184 12872
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 20640 12900 20668 12928
rect 20364 12872 20668 12900
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12801 18015 12835
rect 17957 12795 18015 12801
rect 18141 12835 18199 12841
rect 18141 12801 18153 12835
rect 18187 12801 18199 12835
rect 18141 12795 18199 12801
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 20364 12841 20392 12872
rect 18397 12835 18455 12841
rect 18397 12832 18409 12835
rect 18288 12804 18409 12832
rect 18288 12792 18294 12804
rect 18397 12801 18409 12804
rect 18443 12801 18455 12835
rect 18397 12795 18455 12801
rect 20349 12835 20407 12841
rect 20349 12801 20361 12835
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12832 20591 12835
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20579 12804 20637 12832
rect 20579 12801 20591 12804
rect 20533 12795 20591 12801
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20916 12832 20944 12928
rect 23753 12903 23811 12909
rect 23753 12900 23765 12903
rect 23322 12872 23765 12900
rect 23753 12869 23765 12872
rect 23799 12869 23811 12903
rect 25958 12900 25964 12912
rect 23753 12863 23811 12869
rect 25608 12872 25964 12900
rect 21361 12835 21419 12841
rect 21361 12832 21373 12835
rect 20916 12804 21373 12832
rect 20625 12795 20683 12801
rect 21361 12801 21373 12804
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 23106 12792 23112 12844
rect 23164 12792 23170 12844
rect 23474 12792 23480 12844
rect 23532 12832 23538 12844
rect 25608 12841 25636 12872
rect 25958 12860 25964 12872
rect 26016 12900 26022 12912
rect 26513 12903 26571 12909
rect 26513 12900 26525 12903
rect 26016 12872 26525 12900
rect 26016 12860 26022 12872
rect 26513 12869 26525 12872
rect 26559 12869 26571 12903
rect 26513 12863 26571 12869
rect 28350 12860 28356 12912
rect 28408 12860 28414 12912
rect 29086 12860 29092 12912
rect 29144 12860 29150 12912
rect 23845 12835 23903 12841
rect 23845 12832 23857 12835
rect 23532 12804 23857 12832
rect 23532 12792 23538 12804
rect 23845 12801 23857 12804
rect 23891 12832 23903 12835
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 23891 12804 24900 12832
rect 23891 12801 23903 12804
rect 23845 12795 23903 12801
rect 12268 12736 12756 12764
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12764 13047 12767
rect 13265 12767 13323 12773
rect 13265 12764 13277 12767
rect 13035 12736 13277 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 13265 12733 13277 12736
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 13688 12736 13829 12764
rect 13688 12724 13694 12736
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 15378 12724 15384 12776
rect 15436 12724 15442 12776
rect 16960 12764 16988 12792
rect 17770 12764 17776 12776
rect 16960 12736 17776 12764
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 20165 12767 20223 12773
rect 20165 12733 20177 12767
rect 20211 12733 20223 12767
rect 20165 12727 20223 12733
rect 15396 12696 15424 12724
rect 17681 12699 17739 12705
rect 17681 12696 17693 12699
rect 15396 12668 17693 12696
rect 17681 12665 17693 12668
rect 17727 12665 17739 12699
rect 17681 12659 17739 12665
rect 19521 12699 19579 12705
rect 19521 12665 19533 12699
rect 19567 12696 19579 12699
rect 20180 12696 20208 12727
rect 20898 12724 20904 12776
rect 20956 12764 20962 12776
rect 21177 12767 21235 12773
rect 21177 12764 21189 12767
rect 20956 12736 21189 12764
rect 20956 12724 20962 12736
rect 21177 12733 21189 12736
rect 21223 12733 21235 12767
rect 21177 12727 21235 12733
rect 21542 12724 21548 12776
rect 21600 12764 21606 12776
rect 21821 12767 21879 12773
rect 21821 12764 21833 12767
rect 21600 12736 21833 12764
rect 21600 12724 21606 12736
rect 21821 12733 21833 12736
rect 21867 12733 21879 12767
rect 21821 12727 21879 12733
rect 22094 12724 22100 12776
rect 22152 12724 22158 12776
rect 23124 12764 23152 12792
rect 23569 12767 23627 12773
rect 23569 12764 23581 12767
rect 23124 12736 23581 12764
rect 23569 12733 23581 12736
rect 23615 12733 23627 12767
rect 23569 12727 23627 12733
rect 19567 12668 20208 12696
rect 19567 12665 19579 12668
rect 19521 12659 19579 12665
rect 11514 12588 11520 12640
rect 11572 12588 11578 12640
rect 12342 12588 12348 12640
rect 12400 12588 12406 12640
rect 17586 12588 17592 12640
rect 17644 12588 17650 12640
rect 19610 12588 19616 12640
rect 19668 12588 19674 12640
rect 24872 12628 24900 12804
rect 25056 12804 25421 12832
rect 25056 12773 25084 12804
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 25593 12835 25651 12841
rect 25593 12801 25605 12835
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12832 26479 12835
rect 28721 12835 28779 12841
rect 26467 12804 28028 12832
rect 26467 12801 26479 12804
rect 26421 12795 26479 12801
rect 25041 12767 25099 12773
rect 25041 12764 25053 12767
rect 24964 12736 25053 12764
rect 24964 12708 24992 12736
rect 25041 12733 25053 12736
rect 25087 12733 25099 12767
rect 25041 12727 25099 12733
rect 25225 12767 25283 12773
rect 25225 12733 25237 12767
rect 25271 12764 25283 12767
rect 26142 12764 26148 12776
rect 25271 12736 26148 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 26142 12724 26148 12736
rect 26200 12764 26206 12776
rect 26605 12767 26663 12773
rect 26605 12764 26617 12767
rect 26200 12736 26617 12764
rect 26200 12724 26206 12736
rect 26605 12733 26617 12736
rect 26651 12764 26663 12767
rect 26786 12764 26792 12776
rect 26651 12736 26792 12764
rect 26651 12733 26663 12736
rect 26605 12727 26663 12733
rect 26786 12724 26792 12736
rect 26844 12724 26850 12776
rect 28000 12764 28028 12804
rect 28721 12801 28733 12835
rect 28767 12832 28779 12835
rect 29104 12832 29132 12860
rect 28767 12804 29132 12832
rect 28767 12801 28779 12804
rect 28721 12795 28779 12801
rect 28534 12764 28540 12776
rect 28000 12736 28540 12764
rect 28534 12724 28540 12736
rect 28592 12724 28598 12776
rect 29086 12724 29092 12776
rect 29144 12724 29150 12776
rect 29196 12764 29224 12940
rect 32490 12928 32496 12980
rect 32548 12968 32554 12980
rect 32769 12971 32827 12977
rect 32769 12968 32781 12971
rect 32548 12940 32781 12968
rect 32548 12928 32554 12940
rect 32769 12937 32781 12940
rect 32815 12937 32827 12971
rect 32769 12931 32827 12937
rect 34422 12928 34428 12980
rect 34480 12968 34486 12980
rect 35802 12968 35808 12980
rect 34480 12940 35808 12968
rect 34480 12928 34486 12940
rect 30285 12903 30343 12909
rect 30285 12869 30297 12903
rect 30331 12900 30343 12903
rect 30469 12903 30527 12909
rect 30469 12900 30481 12903
rect 30331 12872 30481 12900
rect 30331 12869 30343 12872
rect 30285 12863 30343 12869
rect 30469 12869 30481 12872
rect 30515 12869 30527 12903
rect 30469 12863 30527 12869
rect 30650 12860 30656 12912
rect 30708 12860 30714 12912
rect 31021 12903 31079 12909
rect 31021 12869 31033 12903
rect 31067 12900 31079 12903
rect 31067 12872 31432 12900
rect 31067 12869 31079 12872
rect 31021 12863 31079 12869
rect 29917 12835 29975 12841
rect 29917 12832 29929 12835
rect 29748 12804 29929 12832
rect 29748 12773 29776 12804
rect 29917 12801 29929 12804
rect 29963 12801 29975 12835
rect 29917 12795 29975 12801
rect 30101 12835 30159 12841
rect 30101 12801 30113 12835
rect 30147 12801 30159 12835
rect 30101 12795 30159 12801
rect 29733 12767 29791 12773
rect 29733 12764 29745 12767
rect 29196 12736 29745 12764
rect 29733 12733 29745 12736
rect 29779 12733 29791 12767
rect 29733 12727 29791 12733
rect 30116 12764 30144 12795
rect 30374 12792 30380 12844
rect 30432 12792 30438 12844
rect 30926 12792 30932 12844
rect 30984 12792 30990 12844
rect 31113 12835 31171 12841
rect 31113 12801 31125 12835
rect 31159 12801 31171 12835
rect 31113 12795 31171 12801
rect 31128 12764 31156 12795
rect 31202 12792 31208 12844
rect 31260 12792 31266 12844
rect 31404 12841 31432 12872
rect 34146 12860 34152 12912
rect 34204 12900 34210 12912
rect 34204 12872 34652 12900
rect 34204 12860 34210 12872
rect 31389 12835 31447 12841
rect 31389 12801 31401 12835
rect 31435 12832 31447 12835
rect 32953 12835 33011 12841
rect 31435 12804 31754 12832
rect 31435 12801 31447 12804
rect 31389 12795 31447 12801
rect 30116 12736 31156 12764
rect 24946 12656 24952 12708
rect 25004 12656 25010 12708
rect 25056 12668 25544 12696
rect 25056 12628 25084 12668
rect 24872 12600 25084 12628
rect 25406 12588 25412 12640
rect 25464 12588 25470 12640
rect 25516 12628 25544 12668
rect 26050 12656 26056 12708
rect 26108 12656 26114 12708
rect 30116 12696 30144 12736
rect 29104 12668 30144 12696
rect 28258 12628 28264 12640
rect 25516 12600 28264 12628
rect 28258 12588 28264 12600
rect 28316 12588 28322 12640
rect 28534 12588 28540 12640
rect 28592 12628 28598 12640
rect 29104 12628 29132 12668
rect 28592 12600 29132 12628
rect 28592 12588 28598 12600
rect 29178 12588 29184 12640
rect 29236 12588 29242 12640
rect 30650 12588 30656 12640
rect 30708 12588 30714 12640
rect 31386 12588 31392 12640
rect 31444 12628 31450 12640
rect 31573 12631 31631 12637
rect 31573 12628 31585 12631
rect 31444 12600 31585 12628
rect 31444 12588 31450 12600
rect 31573 12597 31585 12600
rect 31619 12597 31631 12631
rect 31726 12628 31754 12804
rect 32953 12801 32965 12835
rect 32999 12832 33011 12835
rect 32999 12804 34100 12832
rect 32999 12801 33011 12804
rect 32953 12795 33011 12801
rect 34072 12705 34100 12804
rect 34238 12792 34244 12844
rect 34296 12832 34302 12844
rect 34425 12835 34483 12841
rect 34425 12832 34437 12835
rect 34296 12804 34437 12832
rect 34296 12792 34302 12804
rect 34425 12801 34437 12804
rect 34471 12801 34483 12835
rect 34425 12795 34483 12801
rect 34517 12767 34575 12773
rect 34517 12764 34529 12767
rect 34440 12736 34529 12764
rect 34440 12708 34468 12736
rect 34517 12733 34529 12736
rect 34563 12733 34575 12767
rect 34517 12727 34575 12733
rect 34057 12699 34115 12705
rect 34057 12665 34069 12699
rect 34103 12665 34115 12699
rect 34057 12659 34115 12665
rect 34422 12656 34428 12708
rect 34480 12656 34486 12708
rect 34624 12696 34652 12872
rect 35268 12841 35296 12940
rect 35802 12928 35808 12940
rect 35860 12928 35866 12980
rect 35621 12903 35679 12909
rect 35621 12869 35633 12903
rect 35667 12900 35679 12903
rect 35894 12900 35900 12912
rect 35667 12872 35900 12900
rect 35667 12869 35679 12872
rect 35621 12863 35679 12869
rect 35894 12860 35900 12872
rect 35952 12860 35958 12912
rect 36354 12860 36360 12912
rect 36412 12860 36418 12912
rect 35253 12835 35311 12841
rect 35253 12832 35265 12835
rect 34716 12804 35265 12832
rect 34716 12773 34744 12804
rect 35253 12801 35265 12804
rect 35299 12801 35311 12835
rect 35253 12795 35311 12801
rect 34701 12767 34759 12773
rect 34701 12733 34713 12767
rect 34747 12733 34759 12767
rect 34701 12727 34759 12733
rect 34790 12724 34796 12776
rect 34848 12764 34854 12776
rect 35161 12767 35219 12773
rect 35161 12764 35173 12767
rect 34848 12736 35173 12764
rect 34848 12724 34854 12736
rect 35161 12733 35173 12736
rect 35207 12733 35219 12767
rect 35161 12727 35219 12733
rect 34624 12668 35112 12696
rect 33962 12628 33968 12640
rect 31726 12600 33968 12628
rect 31573 12591 31631 12597
rect 33962 12588 33968 12600
rect 34020 12588 34026 12640
rect 34514 12588 34520 12640
rect 34572 12628 34578 12640
rect 35084 12637 35112 12668
rect 34885 12631 34943 12637
rect 34885 12628 34897 12631
rect 34572 12600 34897 12628
rect 34572 12588 34578 12600
rect 34885 12597 34897 12600
rect 34931 12597 34943 12631
rect 34885 12591 34943 12597
rect 35069 12631 35127 12637
rect 35069 12597 35081 12631
rect 35115 12597 35127 12631
rect 35176 12628 35204 12727
rect 35342 12724 35348 12776
rect 35400 12724 35406 12776
rect 37829 12767 37887 12773
rect 37829 12764 37841 12767
rect 37108 12736 37841 12764
rect 36814 12628 36820 12640
rect 35176 12600 36820 12628
rect 35069 12591 35127 12597
rect 36814 12588 36820 12600
rect 36872 12628 36878 12640
rect 37108 12637 37136 12736
rect 37829 12733 37841 12736
rect 37875 12733 37887 12767
rect 37829 12727 37887 12733
rect 37093 12631 37151 12637
rect 37093 12628 37105 12631
rect 36872 12600 37105 12628
rect 36872 12588 36878 12600
rect 37093 12597 37105 12600
rect 37139 12597 37151 12631
rect 37093 12591 37151 12597
rect 37274 12588 37280 12640
rect 37332 12588 37338 12640
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9674 12424 9680 12436
rect 9447 12396 9680 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13688 12396 13737 12424
rect 13688 12384 13694 12396
rect 13725 12393 13737 12396
rect 13771 12393 13783 12427
rect 13725 12387 13783 12393
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 20070 12424 20076 12436
rect 15528 12396 20076 12424
rect 15528 12384 15534 12396
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 20714 12424 20720 12436
rect 20180 12396 20720 12424
rect 17313 12359 17371 12365
rect 17313 12325 17325 12359
rect 17359 12356 17371 12359
rect 17862 12356 17868 12368
rect 17359 12328 17868 12356
rect 17359 12325 17371 12328
rect 17313 12319 17371 12325
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 20180 12356 20208 12396
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22281 12427 22339 12433
rect 22281 12424 22293 12427
rect 22152 12396 22293 12424
rect 22152 12384 22158 12396
rect 22281 12393 22293 12396
rect 22327 12393 22339 12427
rect 25958 12424 25964 12436
rect 22281 12387 22339 12393
rect 24688 12396 25964 12424
rect 17972 12328 20208 12356
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 11977 12291 12035 12297
rect 11977 12288 11989 12291
rect 11940 12260 11989 12288
rect 11940 12248 11946 12260
rect 11977 12257 11989 12260
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 12342 12288 12348 12300
rect 12299 12260 12348 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 17144 12260 17724 12288
rect 17144 12232 17172 12260
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 10873 12223 10931 12229
rect 9355 12192 9628 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 9600 12164 9628 12192
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 11514 12220 11520 12232
rect 10919 12192 11520 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 17402 12180 17408 12232
rect 17460 12180 17466 12232
rect 17494 12180 17500 12232
rect 17552 12180 17558 12232
rect 17696 12229 17724 12260
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 9582 12112 9588 12164
rect 9640 12112 9646 12164
rect 12986 12112 12992 12164
rect 13044 12112 13050 12164
rect 16482 12112 16488 12164
rect 16540 12152 16546 12164
rect 17972 12152 18000 12328
rect 20622 12316 20628 12368
rect 20680 12316 20686 12368
rect 19429 12291 19487 12297
rect 19429 12257 19441 12291
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 19521 12291 19579 12297
rect 19521 12257 19533 12291
rect 19567 12288 19579 12291
rect 20640 12288 20668 12316
rect 19567 12260 20668 12288
rect 22005 12291 22063 12297
rect 19567 12257 19579 12260
rect 19521 12251 19579 12257
rect 22005 12257 22017 12291
rect 22051 12288 22063 12291
rect 22649 12291 22707 12297
rect 22649 12288 22661 12291
rect 22051 12260 22661 12288
rect 22051 12257 22063 12260
rect 22005 12251 22063 12257
rect 22649 12257 22661 12260
rect 22695 12257 22707 12291
rect 22649 12251 22707 12257
rect 22741 12291 22799 12297
rect 22741 12257 22753 12291
rect 22787 12288 22799 12291
rect 22925 12291 22983 12297
rect 22925 12288 22937 12291
rect 22787 12260 22937 12288
rect 22787 12257 22799 12260
rect 22741 12251 22799 12257
rect 22925 12257 22937 12260
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 16540 12124 18000 12152
rect 19444 12152 19472 12251
rect 19610 12180 19616 12232
rect 19668 12180 19674 12232
rect 20070 12180 20076 12232
rect 20128 12220 20134 12232
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 20128 12192 20637 12220
rect 20128 12180 20134 12192
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 21637 12223 21695 12229
rect 21637 12189 21649 12223
rect 21683 12189 21695 12223
rect 21637 12183 21695 12189
rect 20898 12152 20904 12164
rect 19444 12124 20904 12152
rect 16540 12112 16546 12124
rect 20898 12112 20904 12124
rect 20956 12112 20962 12164
rect 21358 12112 21364 12164
rect 21416 12112 21422 12164
rect 10686 12044 10692 12096
rect 10744 12044 10750 12096
rect 17681 12087 17739 12093
rect 17681 12053 17693 12087
rect 17727 12084 17739 12087
rect 18322 12084 18328 12096
rect 17727 12056 18328 12084
rect 17727 12053 17739 12056
rect 17681 12047 17739 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 18414 12044 18420 12096
rect 18472 12084 18478 12096
rect 19334 12084 19340 12096
rect 18472 12056 19340 12084
rect 18472 12044 18478 12056
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 19978 12044 19984 12096
rect 20036 12044 20042 12096
rect 21652 12084 21680 12183
rect 21818 12180 21824 12232
rect 21876 12180 21882 12232
rect 21910 12180 21916 12232
rect 21968 12220 21974 12232
rect 22465 12223 22523 12229
rect 22465 12220 22477 12223
rect 21968 12192 22477 12220
rect 21968 12180 21974 12192
rect 22465 12189 22477 12192
rect 22511 12189 22523 12223
rect 22465 12183 22523 12189
rect 22833 12223 22891 12229
rect 22833 12189 22845 12223
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 23017 12223 23075 12229
rect 23017 12189 23029 12223
rect 23063 12220 23075 12223
rect 23106 12220 23112 12232
rect 23063 12192 23112 12220
rect 23063 12189 23075 12192
rect 23017 12183 23075 12189
rect 21836 12152 21864 12180
rect 22848 12152 22876 12183
rect 21836 12124 22876 12152
rect 22186 12084 22192 12096
rect 21652 12056 22192 12084
rect 22186 12044 22192 12056
rect 22244 12084 22250 12096
rect 23032 12084 23060 12183
rect 23106 12180 23112 12192
rect 23164 12180 23170 12232
rect 24688 12229 24716 12396
rect 25958 12384 25964 12396
rect 26016 12424 26022 12436
rect 26694 12424 26700 12436
rect 26016 12396 26700 12424
rect 26016 12384 26022 12396
rect 26694 12384 26700 12396
rect 26752 12424 26758 12436
rect 26789 12427 26847 12433
rect 26789 12424 26801 12427
rect 26752 12396 26801 12424
rect 26752 12384 26758 12396
rect 26789 12393 26801 12396
rect 26835 12393 26847 12427
rect 26789 12387 26847 12393
rect 28997 12427 29055 12433
rect 28997 12393 29009 12427
rect 29043 12424 29055 12427
rect 30374 12424 30380 12436
rect 29043 12396 30380 12424
rect 29043 12393 29055 12396
rect 28997 12387 29055 12393
rect 30374 12384 30380 12396
rect 30432 12384 30438 12436
rect 31389 12427 31447 12433
rect 31389 12393 31401 12427
rect 31435 12424 31447 12427
rect 33686 12424 33692 12436
rect 31435 12396 33692 12424
rect 31435 12393 31447 12396
rect 31389 12387 31447 12393
rect 33686 12384 33692 12396
rect 33744 12384 33750 12436
rect 34146 12384 34152 12436
rect 34204 12384 34210 12436
rect 34238 12384 34244 12436
rect 34296 12424 34302 12436
rect 34701 12427 34759 12433
rect 34701 12424 34713 12427
rect 34296 12396 34713 12424
rect 34296 12384 34302 12396
rect 34701 12393 34713 12396
rect 34747 12393 34759 12427
rect 34701 12387 34759 12393
rect 35894 12384 35900 12436
rect 35952 12384 35958 12436
rect 36354 12384 36360 12436
rect 36412 12384 36418 12436
rect 32674 12356 32680 12368
rect 31588 12328 32680 12356
rect 25038 12248 25044 12300
rect 25096 12288 25102 12300
rect 27246 12288 27252 12300
rect 25096 12260 27252 12288
rect 25096 12248 25102 12260
rect 27246 12248 27252 12260
rect 27304 12288 27310 12300
rect 28445 12291 28503 12297
rect 28445 12288 28457 12291
rect 27304 12260 28457 12288
rect 27304 12248 27310 12260
rect 28445 12257 28457 12260
rect 28491 12288 28503 12291
rect 28994 12288 29000 12300
rect 28491 12260 29000 12288
rect 28491 12257 28503 12260
rect 28445 12251 28503 12257
rect 28994 12248 29000 12260
rect 29052 12248 29058 12300
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12220 24823 12223
rect 24946 12220 24952 12232
rect 24811 12192 24952 12220
rect 24811 12189 24823 12192
rect 24765 12183 24823 12189
rect 24688 12152 24716 12183
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 27706 12180 27712 12232
rect 27764 12180 27770 12232
rect 28534 12180 28540 12232
rect 28592 12220 28598 12232
rect 28905 12223 28963 12229
rect 28905 12220 28917 12223
rect 28592 12192 28917 12220
rect 28592 12180 28598 12192
rect 28905 12189 28917 12192
rect 28951 12189 28963 12223
rect 28905 12183 28963 12189
rect 24688 12124 24808 12152
rect 24780 12096 24808 12124
rect 25314 12112 25320 12164
rect 25372 12112 25378 12164
rect 25590 12112 25596 12164
rect 25648 12152 25654 12164
rect 28920 12152 28948 12183
rect 29086 12180 29092 12232
rect 29144 12180 29150 12232
rect 30837 12223 30895 12229
rect 30837 12189 30849 12223
rect 30883 12189 30895 12223
rect 30837 12183 30895 12189
rect 30742 12152 30748 12164
rect 25648 12124 25806 12152
rect 28920 12124 30748 12152
rect 25648 12112 25654 12124
rect 30742 12112 30748 12124
rect 30800 12152 30806 12164
rect 30852 12152 30880 12183
rect 30926 12180 30932 12232
rect 30984 12220 30990 12232
rect 31021 12223 31079 12229
rect 31021 12220 31033 12223
rect 30984 12192 31033 12220
rect 30984 12180 30990 12192
rect 31021 12189 31033 12192
rect 31067 12189 31079 12223
rect 31021 12183 31079 12189
rect 30800 12124 30880 12152
rect 31036 12152 31064 12183
rect 31202 12180 31208 12232
rect 31260 12220 31266 12232
rect 31588 12229 31616 12328
rect 32674 12316 32680 12328
rect 32732 12316 32738 12368
rect 33318 12356 33324 12368
rect 32784 12328 33324 12356
rect 32784 12288 32812 12328
rect 33318 12316 33324 12328
rect 33376 12356 33382 12368
rect 33870 12356 33876 12368
rect 33376 12328 33876 12356
rect 33376 12316 33382 12328
rect 33870 12316 33876 12328
rect 33928 12316 33934 12368
rect 33962 12316 33968 12368
rect 34020 12356 34026 12368
rect 35526 12356 35532 12368
rect 34020 12328 35532 12356
rect 34020 12316 34026 12328
rect 32508 12260 32812 12288
rect 32508 12229 32536 12260
rect 32858 12248 32864 12300
rect 32916 12288 32922 12300
rect 34514 12288 34520 12300
rect 32916 12260 34520 12288
rect 32916 12248 32922 12260
rect 34514 12248 34520 12260
rect 34572 12248 34578 12300
rect 31297 12223 31355 12229
rect 31297 12220 31309 12223
rect 31260 12192 31309 12220
rect 31260 12180 31266 12192
rect 31297 12189 31309 12192
rect 31343 12189 31355 12223
rect 31297 12183 31355 12189
rect 31573 12223 31631 12229
rect 31573 12189 31585 12223
rect 31619 12189 31631 12223
rect 31573 12183 31631 12189
rect 31665 12223 31723 12229
rect 31665 12189 31677 12223
rect 31711 12189 31723 12223
rect 31665 12183 31723 12189
rect 32493 12223 32551 12229
rect 32493 12189 32505 12223
rect 32539 12189 32551 12223
rect 32493 12183 32551 12189
rect 32677 12223 32735 12229
rect 32677 12189 32689 12223
rect 32723 12220 32735 12223
rect 32950 12220 32956 12232
rect 32723 12192 32956 12220
rect 32723 12189 32735 12192
rect 32677 12183 32735 12189
rect 31036 12124 31340 12152
rect 30800 12112 30806 12124
rect 31312 12096 31340 12124
rect 22244 12056 23060 12084
rect 22244 12044 22250 12056
rect 24762 12044 24768 12096
rect 24820 12044 24826 12096
rect 24949 12087 25007 12093
rect 24949 12053 24961 12087
rect 24995 12084 25007 12087
rect 25682 12084 25688 12096
rect 24995 12056 25688 12084
rect 24995 12053 25007 12056
rect 24949 12047 25007 12053
rect 25682 12044 25688 12056
rect 25740 12044 25746 12096
rect 31110 12044 31116 12096
rect 31168 12084 31174 12096
rect 31205 12087 31263 12093
rect 31205 12084 31217 12087
rect 31168 12056 31217 12084
rect 31168 12044 31174 12056
rect 31205 12053 31217 12056
rect 31251 12053 31263 12087
rect 31205 12047 31263 12053
rect 31294 12044 31300 12096
rect 31352 12044 31358 12096
rect 31680 12084 31708 12183
rect 32950 12180 32956 12192
rect 33008 12220 33014 12232
rect 33410 12220 33416 12232
rect 33008 12192 33416 12220
rect 33008 12180 33014 12192
rect 33410 12180 33416 12192
rect 33468 12180 33474 12232
rect 33781 12223 33839 12229
rect 33781 12189 33793 12223
rect 33827 12189 33839 12223
rect 33781 12183 33839 12189
rect 31754 12084 31760 12096
rect 31680 12056 31760 12084
rect 31754 12044 31760 12056
rect 31812 12044 31818 12096
rect 31846 12044 31852 12096
rect 31904 12044 31910 12096
rect 32582 12044 32588 12096
rect 32640 12044 32646 12096
rect 33594 12044 33600 12096
rect 33652 12044 33658 12096
rect 33796 12084 33824 12183
rect 33870 12180 33876 12232
rect 33928 12180 33934 12232
rect 34238 12180 34244 12232
rect 34296 12180 34302 12232
rect 34900 12229 34928 12328
rect 35526 12316 35532 12328
rect 35584 12316 35590 12368
rect 37274 12288 37280 12300
rect 35636 12260 37280 12288
rect 34701 12223 34759 12229
rect 34701 12189 34713 12223
rect 34747 12189 34759 12223
rect 34701 12183 34759 12189
rect 34885 12223 34943 12229
rect 34885 12189 34897 12223
rect 34931 12189 34943 12223
rect 34885 12183 34943 12189
rect 35345 12223 35403 12229
rect 35345 12189 35357 12223
rect 35391 12220 35403 12223
rect 35434 12220 35440 12232
rect 35391 12192 35440 12220
rect 35391 12189 35403 12192
rect 35345 12183 35403 12189
rect 34716 12152 34744 12183
rect 35434 12180 35440 12192
rect 35492 12180 35498 12232
rect 35636 12229 35664 12260
rect 37274 12248 37280 12260
rect 37332 12248 37338 12300
rect 35621 12223 35679 12229
rect 35621 12189 35633 12223
rect 35667 12189 35679 12223
rect 35621 12183 35679 12189
rect 35713 12223 35771 12229
rect 35713 12189 35725 12223
rect 35759 12220 35771 12223
rect 35986 12220 35992 12232
rect 35759 12192 35992 12220
rect 35759 12189 35771 12192
rect 35713 12183 35771 12189
rect 35986 12180 35992 12192
rect 36044 12180 36050 12232
rect 36078 12180 36084 12232
rect 36136 12220 36142 12232
rect 36262 12220 36268 12232
rect 36136 12192 36268 12220
rect 36136 12180 36142 12192
rect 36262 12180 36268 12192
rect 36320 12180 36326 12232
rect 36630 12180 36636 12232
rect 36688 12180 36694 12232
rect 35250 12152 35256 12164
rect 34716 12124 35256 12152
rect 35250 12112 35256 12124
rect 35308 12112 35314 12164
rect 35529 12155 35587 12161
rect 35529 12121 35541 12155
rect 35575 12152 35587 12155
rect 36648 12152 36676 12180
rect 35575 12124 36676 12152
rect 35575 12121 35587 12124
rect 35529 12115 35587 12121
rect 34790 12084 34796 12096
rect 33796 12056 34796 12084
rect 34790 12044 34796 12056
rect 34848 12044 34854 12096
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 13044 11852 13093 11880
rect 13044 11840 13050 11852
rect 13081 11849 13093 11852
rect 13127 11849 13139 11883
rect 13081 11843 13139 11849
rect 17770 11840 17776 11892
rect 17828 11840 17834 11892
rect 17954 11840 17960 11892
rect 18012 11840 18018 11892
rect 21358 11880 21364 11892
rect 19168 11852 21364 11880
rect 15470 11772 15476 11824
rect 15528 11812 15534 11824
rect 15749 11815 15807 11821
rect 15749 11812 15761 11815
rect 15528 11784 15761 11812
rect 15528 11772 15534 11784
rect 15749 11781 15761 11784
rect 15795 11781 15807 11815
rect 15749 11775 15807 11781
rect 16482 11772 16488 11824
rect 16540 11772 16546 11824
rect 17681 11815 17739 11821
rect 17681 11781 17693 11815
rect 17727 11812 17739 11815
rect 17972 11812 18000 11840
rect 17727 11784 18000 11812
rect 17727 11781 17739 11784
rect 17681 11775 17739 11781
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 9640 11716 11713 11744
rect 9640 11704 9646 11716
rect 11701 11713 11713 11716
rect 11747 11744 11759 11747
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 11747 11716 13001 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 12989 11713 13001 11716
rect 13035 11744 13047 11747
rect 16301 11747 16359 11753
rect 13035 11716 13860 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 13832 11620 13860 11716
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16500 11744 16528 11772
rect 16347 11716 16528 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 17126 11704 17132 11756
rect 17184 11704 17190 11756
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11744 17371 11747
rect 17494 11744 17500 11756
rect 17359 11716 17500 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 17494 11704 17500 11716
rect 17552 11744 17558 11756
rect 19168 11753 19196 11852
rect 21358 11840 21364 11852
rect 21416 11880 21422 11892
rect 22554 11880 22560 11892
rect 21416 11852 22560 11880
rect 21416 11840 21422 11852
rect 22554 11840 22560 11852
rect 22612 11840 22618 11892
rect 23247 11883 23305 11889
rect 23247 11849 23259 11883
rect 23293 11880 23305 11883
rect 24946 11880 24952 11892
rect 23293 11852 24952 11880
rect 23293 11849 23305 11852
rect 23247 11843 23305 11849
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 25038 11840 25044 11892
rect 25096 11840 25102 11892
rect 25314 11840 25320 11892
rect 25372 11840 25378 11892
rect 25516 11852 26740 11880
rect 19429 11815 19487 11821
rect 19429 11781 19441 11815
rect 19475 11812 19487 11815
rect 19702 11812 19708 11824
rect 19475 11784 19708 11812
rect 19475 11781 19487 11784
rect 19429 11775 19487 11781
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 21085 11815 21143 11821
rect 21085 11812 21097 11815
rect 20654 11784 21097 11812
rect 21085 11781 21097 11784
rect 21131 11781 21143 11815
rect 21085 11775 21143 11781
rect 21818 11772 21824 11824
rect 21876 11772 21882 11824
rect 22462 11772 22468 11824
rect 22520 11772 22526 11824
rect 23934 11772 23940 11824
rect 23992 11772 23998 11824
rect 19153 11747 19211 11753
rect 17552 11716 17632 11744
rect 17552 11704 17558 11716
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 17604 11685 17632 11716
rect 19153 11713 19165 11747
rect 19199 11713 19211 11747
rect 19153 11707 19211 11713
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11713 21235 11747
rect 21177 11707 21235 11713
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14700 11648 14933 11676
rect 14700 11636 14706 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 17589 11679 17647 11685
rect 17589 11645 17601 11679
rect 17635 11676 17647 11679
rect 17862 11676 17868 11688
rect 17635 11648 17868 11676
rect 17635 11645 17647 11648
rect 17589 11639 17647 11645
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 21192 11676 21220 11707
rect 21726 11704 21732 11756
rect 21784 11744 21790 11756
rect 21910 11744 21916 11756
rect 21784 11716 21916 11744
rect 21784 11704 21790 11716
rect 21910 11704 21916 11716
rect 21968 11744 21974 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21968 11716 22017 11744
rect 21968 11704 21974 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 22005 11707 22063 11713
rect 22112 11716 22385 11744
rect 21818 11676 21824 11688
rect 21192 11648 21824 11676
rect 21818 11636 21824 11648
rect 21876 11636 21882 11688
rect 13814 11568 13820 11620
rect 13872 11608 13878 11620
rect 18782 11608 18788 11620
rect 13872 11580 18788 11608
rect 13872 11568 13878 11580
rect 18782 11568 18788 11580
rect 18840 11568 18846 11620
rect 22112 11608 22140 11716
rect 22373 11713 22385 11716
rect 22419 11713 22431 11747
rect 22480 11744 22508 11772
rect 25056 11753 25084 11840
rect 22833 11747 22891 11753
rect 22833 11744 22845 11747
rect 22480 11716 22845 11744
rect 22373 11707 22431 11713
rect 22833 11713 22845 11716
rect 22879 11713 22891 11747
rect 25052 11747 25110 11753
rect 22833 11707 22891 11713
rect 24596 11728 24992 11744
rect 24596 11716 25018 11728
rect 22186 11636 22192 11688
rect 22244 11636 22250 11688
rect 22278 11636 22284 11688
rect 22336 11676 22342 11688
rect 22557 11679 22615 11685
rect 22557 11676 22569 11679
rect 22336 11648 22569 11676
rect 22336 11636 22342 11648
rect 22557 11645 22569 11648
rect 22603 11645 22615 11679
rect 22557 11639 22615 11645
rect 22649 11679 22707 11685
rect 22649 11645 22661 11679
rect 22695 11676 22707 11679
rect 24596 11676 24624 11716
rect 24964 11700 25018 11716
rect 25052 11713 25064 11747
rect 25098 11713 25110 11747
rect 25052 11707 25110 11713
rect 25222 11704 25228 11756
rect 25280 11744 25286 11756
rect 25516 11753 25544 11852
rect 25590 11772 25596 11824
rect 25648 11812 25654 11824
rect 25648 11784 25820 11812
rect 25648 11772 25654 11784
rect 25501 11747 25559 11753
rect 25501 11744 25513 11747
rect 25280 11716 25513 11744
rect 25280 11704 25286 11716
rect 25501 11713 25513 11716
rect 25547 11713 25559 11747
rect 25501 11707 25559 11713
rect 25682 11704 25688 11756
rect 25740 11704 25746 11756
rect 25792 11753 25820 11784
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11713 25835 11747
rect 25777 11707 25835 11713
rect 26605 11747 26663 11753
rect 26605 11713 26617 11747
rect 26651 11713 26663 11747
rect 26712 11744 26740 11852
rect 26786 11840 26792 11892
rect 26844 11840 26850 11892
rect 27801 11883 27859 11889
rect 27801 11849 27813 11883
rect 27847 11880 27859 11883
rect 28166 11880 28172 11892
rect 27847 11852 28172 11880
rect 27847 11849 27859 11852
rect 27801 11843 27859 11849
rect 28166 11840 28172 11852
rect 28224 11840 28230 11892
rect 30742 11840 30748 11892
rect 30800 11840 30806 11892
rect 31294 11840 31300 11892
rect 31352 11880 31358 11892
rect 32217 11883 32275 11889
rect 32217 11880 32229 11883
rect 31352 11852 32229 11880
rect 31352 11840 31358 11852
rect 32217 11849 32229 11852
rect 32263 11849 32275 11883
rect 32217 11843 32275 11849
rect 33134 11840 33140 11892
rect 33192 11840 33198 11892
rect 33321 11883 33379 11889
rect 33321 11849 33333 11883
rect 33367 11849 33379 11883
rect 33321 11843 33379 11849
rect 27893 11815 27951 11821
rect 27893 11812 27905 11815
rect 27172 11784 27905 11812
rect 27172 11756 27200 11784
rect 27893 11781 27905 11784
rect 27939 11781 27951 11815
rect 27893 11775 27951 11781
rect 30006 11772 30012 11824
rect 30064 11772 30070 11824
rect 30760 11812 30788 11840
rect 31389 11815 31447 11821
rect 31389 11812 31401 11815
rect 30760 11784 31401 11812
rect 31389 11781 31401 11784
rect 31435 11781 31447 11815
rect 33336 11812 33364 11843
rect 34606 11840 34612 11892
rect 34664 11880 34670 11892
rect 34701 11883 34759 11889
rect 34701 11880 34713 11883
rect 34664 11852 34713 11880
rect 34664 11840 34670 11852
rect 34701 11849 34713 11852
rect 34747 11849 34759 11883
rect 34701 11843 34759 11849
rect 31389 11775 31447 11781
rect 32416 11784 33364 11812
rect 27154 11744 27160 11756
rect 26712 11716 27160 11744
rect 26605 11707 26663 11713
rect 22695 11648 24624 11676
rect 24673 11679 24731 11685
rect 22695 11645 22707 11648
rect 22649 11639 22707 11645
rect 24673 11645 24685 11679
rect 24719 11676 24731 11679
rect 24854 11676 24860 11688
rect 24719 11648 24860 11676
rect 24719 11645 24731 11648
rect 24673 11639 24731 11645
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 24990 11676 25018 11700
rect 26620 11676 26648 11707
rect 27154 11704 27160 11716
rect 27212 11704 27218 11756
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11744 27399 11747
rect 28261 11747 28319 11753
rect 28261 11744 28273 11747
rect 27387 11716 28273 11744
rect 27387 11713 27399 11716
rect 27341 11707 27399 11713
rect 28261 11713 28273 11716
rect 28307 11713 28319 11747
rect 28261 11707 28319 11713
rect 28994 11704 29000 11756
rect 29052 11704 29058 11756
rect 31205 11747 31263 11753
rect 31205 11713 31217 11747
rect 31251 11713 31263 11747
rect 31205 11707 31263 11713
rect 24990 11648 25077 11676
rect 26620 11648 27476 11676
rect 20824 11580 22140 11608
rect 11606 11500 11612 11552
rect 11664 11500 11670 11552
rect 16390 11500 16396 11552
rect 16448 11500 16454 11552
rect 16945 11543 17003 11549
rect 16945 11509 16957 11543
rect 16991 11540 17003 11543
rect 18046 11540 18052 11552
rect 16991 11512 18052 11540
rect 16991 11509 17003 11512
rect 16945 11503 17003 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18138 11500 18144 11552
rect 18196 11500 18202 11552
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 20824 11540 20852 11580
rect 22370 11568 22376 11620
rect 22428 11568 22434 11620
rect 22741 11611 22799 11617
rect 22741 11577 22753 11611
rect 22787 11608 22799 11611
rect 25049 11608 25077 11648
rect 22787 11580 23980 11608
rect 25049 11580 25820 11608
rect 22787 11577 22799 11580
rect 22741 11571 22799 11577
rect 18748 11512 20852 11540
rect 18748 11500 18754 11512
rect 20898 11500 20904 11552
rect 20956 11500 20962 11552
rect 22388 11540 22416 11568
rect 23017 11543 23075 11549
rect 23017 11540 23029 11543
rect 22388 11512 23029 11540
rect 23017 11509 23029 11512
rect 23063 11509 23075 11543
rect 23952 11540 23980 11580
rect 25222 11540 25228 11552
rect 23952 11512 25228 11540
rect 23017 11503 23075 11509
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 25792 11540 25820 11580
rect 25958 11568 25964 11620
rect 26016 11608 26022 11620
rect 27448 11617 27476 11648
rect 28074 11636 28080 11688
rect 28132 11676 28138 11688
rect 28810 11676 28816 11688
rect 28132 11648 28816 11676
rect 28132 11636 28138 11648
rect 28810 11636 28816 11648
rect 28868 11636 28874 11688
rect 29273 11679 29331 11685
rect 29273 11645 29285 11679
rect 29319 11676 29331 11679
rect 30650 11676 30656 11688
rect 29319 11648 30656 11676
rect 29319 11645 29331 11648
rect 29273 11639 29331 11645
rect 30650 11636 30656 11648
rect 30708 11636 30714 11688
rect 27249 11611 27307 11617
rect 27249 11608 27261 11611
rect 26016 11580 27261 11608
rect 26016 11568 26022 11580
rect 27249 11577 27261 11580
rect 27295 11577 27307 11611
rect 27249 11571 27307 11577
rect 27433 11611 27491 11617
rect 27433 11577 27445 11611
rect 27479 11577 27491 11611
rect 27433 11571 27491 11577
rect 30282 11540 30288 11552
rect 25792 11512 30288 11540
rect 30282 11500 30288 11512
rect 30340 11500 30346 11552
rect 31018 11500 31024 11552
rect 31076 11500 31082 11552
rect 31220 11540 31248 11707
rect 31294 11704 31300 11756
rect 31352 11704 31358 11756
rect 32416 11753 32444 11784
rect 33410 11772 33416 11824
rect 33468 11812 33474 11824
rect 33965 11815 34023 11821
rect 33965 11812 33977 11815
rect 33468 11784 33977 11812
rect 33468 11772 33474 11784
rect 33965 11781 33977 11784
rect 34011 11781 34023 11815
rect 34716 11812 34744 11843
rect 35250 11840 35256 11892
rect 35308 11880 35314 11892
rect 35434 11880 35440 11892
rect 35308 11852 35440 11880
rect 35308 11840 35314 11852
rect 35434 11840 35440 11852
rect 35492 11840 35498 11892
rect 34716 11784 35388 11812
rect 33965 11775 34023 11781
rect 31507 11747 31565 11753
rect 31507 11744 31519 11747
rect 31404 11716 31519 11744
rect 31404 11688 31432 11716
rect 31507 11713 31519 11716
rect 31553 11713 31565 11747
rect 31507 11707 31565 11713
rect 32401 11747 32459 11753
rect 32401 11713 32413 11747
rect 32447 11713 32459 11747
rect 32401 11707 32459 11713
rect 32766 11704 32772 11756
rect 32824 11704 32830 11756
rect 32858 11704 32864 11756
rect 32916 11742 32922 11756
rect 32953 11747 33011 11753
rect 32953 11742 32965 11747
rect 32916 11714 32965 11742
rect 32916 11704 32922 11714
rect 32953 11713 32965 11714
rect 32999 11713 33011 11747
rect 32953 11707 33011 11713
rect 33134 11704 33140 11756
rect 33192 11753 33198 11756
rect 33192 11747 33224 11753
rect 33212 11744 33224 11747
rect 33505 11747 33563 11753
rect 33212 11714 33241 11744
rect 33212 11713 33224 11714
rect 33192 11707 33224 11713
rect 33505 11713 33517 11747
rect 33551 11744 33563 11747
rect 33686 11744 33692 11756
rect 33551 11716 33692 11744
rect 33551 11713 33563 11716
rect 33505 11707 33563 11713
rect 33192 11704 33198 11707
rect 33686 11704 33692 11716
rect 33744 11704 33750 11756
rect 34790 11704 34796 11756
rect 34848 11744 34854 11756
rect 35360 11753 35388 11784
rect 34885 11747 34943 11753
rect 34885 11744 34897 11747
rect 34848 11716 34897 11744
rect 34848 11704 34854 11716
rect 34885 11713 34897 11716
rect 34931 11713 34943 11747
rect 34885 11707 34943 11713
rect 35345 11747 35403 11753
rect 35345 11713 35357 11747
rect 35391 11713 35403 11747
rect 35345 11707 35403 11713
rect 31386 11636 31392 11688
rect 31444 11636 31450 11688
rect 31662 11636 31668 11688
rect 31720 11636 31726 11688
rect 32876 11608 32904 11704
rect 33597 11679 33655 11685
rect 33597 11676 33609 11679
rect 33428 11648 33609 11676
rect 32784 11580 32904 11608
rect 32784 11552 32812 11580
rect 33226 11568 33232 11620
rect 33284 11568 33290 11620
rect 31754 11540 31760 11552
rect 31220 11512 31760 11540
rect 31754 11500 31760 11512
rect 31812 11500 31818 11552
rect 32490 11500 32496 11552
rect 32548 11500 32554 11552
rect 32766 11500 32772 11552
rect 32824 11500 32830 11552
rect 32858 11500 32864 11552
rect 32916 11500 32922 11552
rect 33244 11540 33272 11568
rect 33428 11540 33456 11648
rect 33597 11645 33609 11648
rect 33643 11645 33655 11679
rect 33597 11639 33655 11645
rect 34422 11636 34428 11688
rect 34480 11676 34486 11688
rect 35069 11679 35127 11685
rect 35069 11676 35081 11679
rect 34480 11648 35081 11676
rect 34480 11636 34486 11648
rect 35069 11645 35081 11648
rect 35115 11645 35127 11679
rect 35069 11639 35127 11645
rect 33244 11512 33456 11540
rect 33594 11500 33600 11552
rect 33652 11500 33658 11552
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 10584 11339 10642 11345
rect 10584 11305 10596 11339
rect 10630 11336 10642 11339
rect 10686 11336 10692 11348
rect 10630 11308 10692 11336
rect 10630 11305 10642 11308
rect 10584 11299 10642 11305
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 18138 11296 18144 11348
rect 18196 11296 18202 11348
rect 18690 11296 18696 11348
rect 18748 11296 18754 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 19429 11339 19487 11345
rect 19429 11336 19441 11339
rect 19392 11308 19441 11336
rect 19392 11296 19398 11308
rect 19429 11305 19441 11308
rect 19475 11305 19487 11339
rect 19429 11299 19487 11305
rect 19702 11296 19708 11348
rect 19760 11296 19766 11348
rect 20622 11296 20628 11348
rect 20680 11336 20686 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20680 11308 21005 11336
rect 20680 11296 20686 11308
rect 20993 11305 21005 11308
rect 21039 11336 21051 11339
rect 21726 11336 21732 11348
rect 21039 11308 21732 11336
rect 21039 11305 21051 11308
rect 20993 11299 21051 11305
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 23934 11296 23940 11348
rect 23992 11296 23998 11348
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 25958 11336 25964 11348
rect 24912 11308 25964 11336
rect 24912 11296 24918 11308
rect 25958 11296 25964 11308
rect 26016 11296 26022 11348
rect 26712 11308 28764 11336
rect 18046 11268 18052 11280
rect 17972 11240 18052 11268
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 15657 11203 15715 11209
rect 10367 11172 14688 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 14660 11144 14688 11172
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 17972 11200 18000 11240
rect 18046 11228 18052 11240
rect 18104 11228 18110 11280
rect 15703 11172 18000 11200
rect 18156 11200 18184 11296
rect 19245 11271 19303 11277
rect 19245 11268 19257 11271
rect 18616 11240 19257 11268
rect 18156 11172 18368 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 11664 11104 11730 11132
rect 11664 11092 11670 11104
rect 12158 11092 12164 11144
rect 12216 11132 12222 11144
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 12216 11104 12357 11132
rect 12216 11092 12222 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 14642 11092 14648 11144
rect 14700 11132 14706 11144
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 14700 11104 15393 11132
rect 14700 11092 14706 11104
rect 15381 11101 15393 11104
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 17126 11092 17132 11144
rect 17184 11132 17190 11144
rect 17405 11135 17463 11141
rect 17405 11132 17417 11135
rect 17184 11104 17417 11132
rect 17184 11092 17190 11104
rect 17405 11101 17417 11104
rect 17451 11101 17463 11135
rect 17405 11095 17463 11101
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 16390 11024 16396 11076
rect 16448 11024 16454 11076
rect 18064 11064 18092 11095
rect 18138 11092 18144 11144
rect 18196 11092 18202 11144
rect 18340 11064 18368 11172
rect 18616 11141 18644 11240
rect 19245 11237 19257 11240
rect 19291 11237 19303 11271
rect 26712 11268 26740 11308
rect 19245 11231 19303 11237
rect 19812 11240 26740 11268
rect 18690 11160 18696 11212
rect 18748 11200 18754 11212
rect 19702 11200 19708 11212
rect 18748 11172 19708 11200
rect 18748 11160 18754 11172
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 18568 11135 18644 11141
rect 18568 11101 18580 11135
rect 18614 11104 18644 11135
rect 18614 11101 18626 11104
rect 18568 11095 18626 11101
rect 18782 11092 18788 11144
rect 18840 11132 18846 11144
rect 19812 11132 19840 11240
rect 26786 11228 26792 11280
rect 26844 11268 26850 11280
rect 26844 11240 27384 11268
rect 26844 11228 26850 11240
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11200 20499 11203
rect 20898 11200 20904 11212
rect 20487 11172 20904 11200
rect 20487 11169 20499 11172
rect 20441 11163 20499 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 22186 11200 22192 11212
rect 21652 11172 22192 11200
rect 18840 11104 19840 11132
rect 19889 11135 19947 11141
rect 18840 11092 18846 11104
rect 19889 11101 19901 11135
rect 19935 11132 19947 11135
rect 19996 11132 20024 11160
rect 19935 11104 20024 11132
rect 20257 11135 20315 11141
rect 19935 11101 19947 11104
rect 19889 11095 19947 11101
rect 20257 11101 20269 11135
rect 20303 11132 20315 11135
rect 20303 11104 20392 11132
rect 20303 11101 20315 11104
rect 20257 11095 20315 11101
rect 18443 11067 18501 11073
rect 18443 11064 18455 11067
rect 18064 11036 18276 11064
rect 18340 11036 18455 11064
rect 18248 10996 18276 11036
rect 18443 11033 18455 11036
rect 18489 11033 18501 11067
rect 19242 11064 19248 11076
rect 18443 11027 18501 11033
rect 18616 11036 19248 11064
rect 18616 10996 18644 11036
rect 19242 11024 19248 11036
rect 19300 11064 19306 11076
rect 19613 11067 19671 11073
rect 19613 11064 19625 11067
rect 19300 11036 19625 11064
rect 19300 11024 19306 11036
rect 19613 11033 19625 11036
rect 19659 11033 19671 11067
rect 19613 11027 19671 11033
rect 19702 11024 19708 11076
rect 19760 11064 19766 11076
rect 20073 11067 20131 11073
rect 20073 11064 20085 11067
rect 19760 11036 20085 11064
rect 19760 11024 19766 11036
rect 20073 11033 20085 11036
rect 20119 11064 20131 11067
rect 20364 11064 20392 11104
rect 20806 11092 20812 11144
rect 20864 11092 20870 11144
rect 21652 11141 21680 11172
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 27246 11160 27252 11212
rect 27304 11160 27310 11212
rect 27356 11200 27384 11240
rect 27525 11203 27583 11209
rect 27525 11200 27537 11203
rect 27356 11172 27537 11200
rect 27525 11169 27537 11172
rect 27571 11169 27583 11203
rect 28736 11200 28764 11308
rect 28810 11296 28816 11348
rect 28868 11336 28874 11348
rect 28997 11339 29055 11345
rect 28997 11336 29009 11339
rect 28868 11308 29009 11336
rect 28868 11296 28874 11308
rect 28997 11305 29009 11308
rect 29043 11305 29055 11339
rect 28997 11299 29055 11305
rect 30006 11296 30012 11348
rect 30064 11336 30070 11348
rect 30101 11339 30159 11345
rect 30101 11336 30113 11339
rect 30064 11308 30113 11336
rect 30064 11296 30070 11308
rect 30101 11305 30113 11308
rect 30147 11305 30159 11339
rect 30101 11299 30159 11305
rect 31205 11339 31263 11345
rect 31205 11305 31217 11339
rect 31251 11336 31263 11339
rect 31294 11336 31300 11348
rect 31251 11308 31300 11336
rect 31251 11305 31263 11308
rect 31205 11299 31263 11305
rect 31294 11296 31300 11308
rect 31352 11296 31358 11348
rect 31754 11296 31760 11348
rect 31812 11296 31818 11348
rect 31846 11296 31852 11348
rect 31904 11336 31910 11348
rect 34057 11339 34115 11345
rect 31904 11308 32444 11336
rect 31904 11296 31910 11308
rect 31938 11268 31944 11280
rect 30024 11240 31944 11268
rect 30024 11200 30052 11240
rect 31938 11228 31944 11240
rect 31996 11228 32002 11280
rect 28736 11172 30052 11200
rect 27525 11163 27583 11169
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 21726 11092 21732 11144
rect 21784 11092 21790 11144
rect 21818 11092 21824 11144
rect 21876 11132 21882 11144
rect 23842 11132 23848 11144
rect 21876 11104 23848 11132
rect 21876 11092 21882 11104
rect 23842 11092 23848 11104
rect 23900 11092 23906 11144
rect 25498 11092 25504 11144
rect 25556 11092 25562 11144
rect 25685 11135 25743 11141
rect 25685 11101 25697 11135
rect 25731 11132 25743 11135
rect 25774 11132 25780 11144
rect 25731 11104 25780 11132
rect 25731 11101 25743 11104
rect 25685 11095 25743 11101
rect 25774 11092 25780 11104
rect 25832 11092 25838 11144
rect 30024 11141 30052 11172
rect 30282 11160 30288 11212
rect 30340 11200 30346 11212
rect 30340 11172 31800 11200
rect 30340 11160 30346 11172
rect 25869 11135 25927 11141
rect 25869 11101 25881 11135
rect 25915 11101 25927 11135
rect 25869 11095 25927 11101
rect 29273 11135 29331 11141
rect 29273 11101 29285 11135
rect 29319 11101 29331 11135
rect 29273 11095 29331 11101
rect 30009 11135 30067 11141
rect 30009 11101 30021 11135
rect 30055 11101 30067 11135
rect 30009 11095 30067 11101
rect 20714 11064 20720 11076
rect 20119 11036 20300 11064
rect 20364 11036 20720 11064
rect 20119 11033 20131 11036
rect 20073 11027 20131 11033
rect 20272 11008 20300 11036
rect 20714 11024 20720 11036
rect 20772 11064 20778 11076
rect 21453 11067 21511 11073
rect 21453 11064 21465 11067
rect 20772 11036 21465 11064
rect 20772 11024 20778 11036
rect 21453 11033 21465 11036
rect 21499 11033 21511 11067
rect 21453 11027 21511 11033
rect 25130 11024 25136 11076
rect 25188 11064 25194 11076
rect 25884 11064 25912 11095
rect 29181 11067 29239 11073
rect 29181 11064 29193 11067
rect 25188 11036 25912 11064
rect 28750 11036 29193 11064
rect 25188 11024 25194 11036
rect 29181 11033 29193 11036
rect 29227 11033 29239 11067
rect 29181 11027 29239 11033
rect 29288 11008 29316 11095
rect 31202 11092 31208 11144
rect 31260 11092 31266 11144
rect 31389 11135 31447 11141
rect 31389 11101 31401 11135
rect 31435 11132 31447 11135
rect 31478 11132 31484 11144
rect 31435 11104 31484 11132
rect 31435 11101 31447 11104
rect 31389 11095 31447 11101
rect 31478 11092 31484 11104
rect 31536 11132 31542 11144
rect 31662 11132 31668 11144
rect 31536 11104 31668 11132
rect 31536 11092 31542 11104
rect 31662 11092 31668 11104
rect 31720 11092 31726 11144
rect 31220 11064 31248 11092
rect 31570 11064 31576 11076
rect 31220 11036 31576 11064
rect 31570 11024 31576 11036
rect 31628 11024 31634 11076
rect 18248 10968 18644 10996
rect 19408 10999 19466 11005
rect 19408 10965 19420 10999
rect 19454 10996 19466 10999
rect 20162 10996 20168 11008
rect 19454 10968 20168 10996
rect 19454 10965 19466 10968
rect 19408 10959 19466 10965
rect 20162 10956 20168 10968
rect 20220 10956 20226 11008
rect 20254 10956 20260 11008
rect 20312 10956 20318 11008
rect 25314 10956 25320 11008
rect 25372 10996 25378 11008
rect 25501 10999 25559 11005
rect 25501 10996 25513 10999
rect 25372 10968 25513 10996
rect 25372 10956 25378 10968
rect 25501 10965 25513 10968
rect 25547 10965 25559 10999
rect 25501 10959 25559 10965
rect 25958 10956 25964 11008
rect 26016 10956 26022 11008
rect 28258 10956 28264 11008
rect 28316 10996 28322 11008
rect 29270 10996 29276 11008
rect 28316 10968 29276 10996
rect 28316 10956 28322 10968
rect 29270 10956 29276 10968
rect 29328 10956 29334 11008
rect 31680 10996 31708 11092
rect 31772 11064 31800 11172
rect 31846 11092 31852 11144
rect 31904 11092 31910 11144
rect 32416 11141 32444 11308
rect 34057 11305 34069 11339
rect 34103 11336 34115 11339
rect 34330 11336 34336 11348
rect 34103 11308 34336 11336
rect 34103 11305 34115 11308
rect 34057 11299 34115 11305
rect 34330 11296 34336 11308
rect 34388 11296 34394 11348
rect 32493 11271 32551 11277
rect 32493 11237 32505 11271
rect 32539 11268 32551 11271
rect 32766 11268 32772 11280
rect 32539 11240 32772 11268
rect 32539 11237 32551 11240
rect 32493 11231 32551 11237
rect 32766 11228 32772 11240
rect 32824 11228 32830 11280
rect 34256 11240 35388 11268
rect 32582 11160 32588 11212
rect 32640 11160 32646 11212
rect 32953 11203 33011 11209
rect 32953 11169 32965 11203
rect 32999 11169 33011 11203
rect 32953 11163 33011 11169
rect 33413 11203 33471 11209
rect 33413 11169 33425 11203
rect 33459 11200 33471 11203
rect 33686 11200 33692 11212
rect 33459 11172 33692 11200
rect 33459 11169 33471 11172
rect 33413 11163 33471 11169
rect 32217 11135 32275 11141
rect 32217 11101 32229 11135
rect 32263 11101 32275 11135
rect 32217 11095 32275 11101
rect 32401 11135 32459 11141
rect 32401 11101 32413 11135
rect 32447 11101 32459 11135
rect 32401 11095 32459 11101
rect 32232 11064 32260 11095
rect 32490 11092 32496 11144
rect 32548 11132 32554 11144
rect 32676 11135 32734 11141
rect 32676 11132 32688 11135
rect 32548 11104 32688 11132
rect 32548 11092 32554 11104
rect 32676 11101 32688 11104
rect 32722 11101 32734 11135
rect 32676 11095 32734 11101
rect 32861 11135 32919 11141
rect 32861 11101 32873 11135
rect 32907 11101 32919 11135
rect 32861 11095 32919 11101
rect 31772 11036 32260 11064
rect 32306 11024 32312 11076
rect 32364 11064 32370 11076
rect 32876 11064 32904 11095
rect 32364 11036 32904 11064
rect 32968 11064 32996 11163
rect 33318 11092 33324 11144
rect 33376 11092 33382 11144
rect 33134 11064 33140 11076
rect 32968 11036 33140 11064
rect 32364 11024 32370 11036
rect 33134 11024 33140 11036
rect 33192 11024 33198 11076
rect 33428 10996 33456 11163
rect 33686 11160 33692 11172
rect 33744 11160 33750 11212
rect 34256 11144 34284 11240
rect 34330 11160 34336 11212
rect 34388 11200 34394 11212
rect 35250 11200 35256 11212
rect 34388 11172 34468 11200
rect 34388 11160 34394 11172
rect 34238 11092 34244 11144
rect 34296 11092 34302 11144
rect 34440 11064 34468 11172
rect 34624 11172 35256 11200
rect 34624 11144 34652 11172
rect 35250 11160 35256 11172
rect 35308 11160 35314 11212
rect 35360 11200 35388 11240
rect 36170 11200 36176 11212
rect 35360 11172 36176 11200
rect 36170 11160 36176 11172
rect 36228 11160 36234 11212
rect 34514 11092 34520 11144
rect 34572 11092 34578 11144
rect 34606 11092 34612 11144
rect 34664 11092 34670 11144
rect 34701 11135 34759 11141
rect 34701 11101 34713 11135
rect 34747 11101 34759 11135
rect 34701 11095 34759 11101
rect 34977 11135 35035 11141
rect 34977 11101 34989 11135
rect 35023 11132 35035 11135
rect 35066 11132 35072 11144
rect 35023 11104 35072 11132
rect 35023 11101 35035 11104
rect 34977 11095 35035 11101
rect 34716 11064 34744 11095
rect 35066 11092 35072 11104
rect 35124 11092 35130 11144
rect 34440 11036 34744 11064
rect 34793 11067 34851 11073
rect 34793 11033 34805 11067
rect 34839 11064 34851 11067
rect 35161 11067 35219 11073
rect 34839 11036 35112 11064
rect 34839 11033 34851 11036
rect 34793 11027 34851 11033
rect 31680 10968 33456 10996
rect 33594 10956 33600 11008
rect 33652 10996 33658 11008
rect 34425 10999 34483 11005
rect 34425 10996 34437 10999
rect 33652 10968 34437 10996
rect 33652 10956 33658 10968
rect 34425 10965 34437 10968
rect 34471 10996 34483 10999
rect 34698 10996 34704 11008
rect 34471 10968 34704 10996
rect 34471 10965 34483 10968
rect 34425 10959 34483 10965
rect 34698 10956 34704 10968
rect 34756 10956 34762 11008
rect 35084 10996 35112 11036
rect 35161 11033 35173 11067
rect 35207 11064 35219 11067
rect 35529 11067 35587 11073
rect 35529 11064 35541 11067
rect 35207 11036 35541 11064
rect 35207 11033 35219 11036
rect 35161 11027 35219 11033
rect 35529 11033 35541 11036
rect 35575 11033 35587 11067
rect 36814 11064 36820 11076
rect 36754 11036 36820 11064
rect 35529 11027 35587 11033
rect 36814 11024 36820 11036
rect 36872 11024 36878 11076
rect 35894 10996 35900 11008
rect 35084 10968 35900 10996
rect 35894 10956 35900 10968
rect 35952 10956 35958 11008
rect 36538 10956 36544 11008
rect 36596 10996 36602 11008
rect 37001 10999 37059 11005
rect 37001 10996 37013 10999
rect 36596 10968 37013 10996
rect 36596 10956 36602 10968
rect 37001 10965 37013 10968
rect 37047 10965 37059 10999
rect 37001 10959 37059 10965
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 18046 10752 18052 10804
rect 18104 10752 18110 10804
rect 18156 10764 18828 10792
rect 16853 10727 16911 10733
rect 16853 10693 16865 10727
rect 16899 10724 16911 10727
rect 17586 10724 17592 10736
rect 16899 10696 17592 10724
rect 16899 10693 16911 10696
rect 16853 10687 16911 10693
rect 17586 10684 17592 10696
rect 17644 10724 17650 10736
rect 18156 10724 18184 10764
rect 17644 10696 18184 10724
rect 17644 10684 17650 10696
rect 18230 10684 18236 10736
rect 18288 10684 18294 10736
rect 18322 10684 18328 10736
rect 18380 10684 18386 10736
rect 18414 10684 18420 10736
rect 18472 10684 18478 10736
rect 18555 10727 18613 10733
rect 18555 10693 18567 10727
rect 18601 10724 18613 10727
rect 18690 10724 18696 10736
rect 18601 10696 18696 10724
rect 18601 10693 18613 10696
rect 18555 10687 18613 10693
rect 18690 10684 18696 10696
rect 18748 10684 18754 10736
rect 18234 10681 18292 10684
rect 16482 10616 16488 10668
rect 16540 10665 16546 10668
rect 16540 10656 16551 10665
rect 17037 10659 17095 10665
rect 16540 10628 16585 10656
rect 16540 10619 16551 10628
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 16540 10616 16546 10619
rect 17052 10588 17080 10619
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 17313 10659 17371 10665
rect 17313 10656 17325 10659
rect 17184 10628 17325 10656
rect 17184 10616 17190 10628
rect 17313 10625 17325 10628
rect 17359 10625 17371 10659
rect 17313 10619 17371 10625
rect 17678 10616 17684 10668
rect 17736 10616 17742 10668
rect 18234 10647 18246 10681
rect 18280 10647 18292 10681
rect 18800 10665 18828 10764
rect 19058 10752 19064 10804
rect 19116 10792 19122 10804
rect 20714 10792 20720 10804
rect 19116 10764 20720 10792
rect 19116 10752 19122 10764
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 21821 10795 21879 10801
rect 21821 10761 21833 10795
rect 21867 10792 21879 10795
rect 22278 10792 22284 10804
rect 21867 10764 22284 10792
rect 21867 10761 21879 10764
rect 21821 10755 21879 10761
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 28350 10752 28356 10804
rect 28408 10752 28414 10804
rect 32950 10752 32956 10804
rect 33008 10752 33014 10804
rect 34514 10752 34520 10804
rect 34572 10792 34578 10804
rect 34993 10795 35051 10801
rect 34993 10792 35005 10795
rect 34572 10764 35005 10792
rect 34572 10752 34578 10764
rect 34993 10761 35005 10764
rect 35039 10792 35051 10795
rect 35039 10764 35112 10792
rect 35039 10761 35051 10764
rect 34993 10755 35051 10761
rect 19153 10727 19211 10733
rect 19153 10724 19165 10727
rect 18892 10696 19165 10724
rect 18234 10641 18292 10647
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10625 18843 10659
rect 18785 10619 18843 10625
rect 17696 10588 17724 10616
rect 17052 10560 17724 10588
rect 17957 10591 18015 10597
rect 17957 10557 17969 10591
rect 18003 10588 18015 10591
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18003 10560 18705 10588
rect 18003 10557 18015 10560
rect 17957 10551 18015 10557
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 17126 10480 17132 10532
rect 17184 10520 17190 10532
rect 17184 10492 17816 10520
rect 17184 10480 17190 10492
rect 16390 10412 16396 10464
rect 16448 10412 16454 10464
rect 17218 10412 17224 10464
rect 17276 10412 17282 10464
rect 17788 10452 17816 10492
rect 18892 10452 18920 10696
rect 19153 10693 19165 10696
rect 19199 10724 19211 10727
rect 19334 10724 19340 10736
rect 19199 10696 19340 10724
rect 19199 10693 19211 10696
rect 19153 10687 19211 10693
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 22462 10684 22468 10736
rect 22520 10684 22526 10736
rect 23658 10684 23664 10736
rect 23716 10684 23722 10736
rect 26694 10684 26700 10736
rect 26752 10724 26758 10736
rect 27065 10727 27123 10733
rect 26752 10696 27016 10724
rect 26752 10684 26758 10696
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10625 19303 10659
rect 19245 10619 19303 10625
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 19260 10588 19288 10619
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19484 10628 19717 10656
rect 19484 10616 19490 10628
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 19978 10616 19984 10668
rect 20036 10656 20042 10668
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 20036 10628 22017 10656
rect 20036 10616 20042 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22554 10616 22560 10668
rect 22612 10656 22618 10668
rect 22741 10659 22799 10665
rect 22741 10656 22753 10659
rect 22612 10628 22753 10656
rect 22612 10616 22618 10628
rect 22741 10625 22753 10628
rect 22787 10625 22799 10659
rect 22741 10619 22799 10625
rect 25314 10616 25320 10668
rect 25372 10656 25378 10668
rect 25777 10659 25835 10665
rect 25777 10656 25789 10659
rect 25372 10628 25789 10656
rect 25372 10616 25378 10628
rect 25777 10625 25789 10628
rect 25823 10625 25835 10659
rect 25777 10619 25835 10625
rect 25866 10616 25872 10668
rect 25924 10616 25930 10668
rect 25958 10616 25964 10668
rect 26016 10656 26022 10668
rect 26145 10659 26203 10665
rect 26145 10656 26157 10659
rect 26016 10628 26157 10656
rect 26016 10616 26022 10628
rect 26145 10625 26157 10628
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 26510 10616 26516 10668
rect 26568 10656 26574 10668
rect 26988 10665 27016 10696
rect 27065 10693 27077 10727
rect 27111 10724 27123 10727
rect 28166 10724 28172 10736
rect 27111 10696 28172 10724
rect 27111 10693 27123 10696
rect 27065 10687 27123 10693
rect 26605 10659 26663 10665
rect 26605 10656 26617 10659
rect 26568 10628 26617 10656
rect 26568 10616 26574 10628
rect 26605 10625 26617 10628
rect 26651 10656 26663 10659
rect 26973 10659 27031 10665
rect 26651 10628 26924 10656
rect 26651 10625 26663 10628
rect 26605 10619 26663 10625
rect 19208 10560 19288 10588
rect 19797 10591 19855 10597
rect 19208 10548 19214 10560
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 22097 10591 22155 10597
rect 22097 10588 22109 10591
rect 19843 10560 22109 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 22097 10557 22109 10560
rect 22143 10557 22155 10591
rect 22097 10551 22155 10557
rect 23017 10591 23075 10597
rect 23017 10557 23029 10591
rect 23063 10588 23075 10591
rect 24486 10588 24492 10600
rect 23063 10560 24492 10588
rect 23063 10557 23075 10560
rect 23017 10551 23075 10557
rect 19426 10480 19432 10532
rect 19484 10520 19490 10532
rect 19812 10520 19840 10551
rect 24486 10548 24492 10560
rect 24544 10548 24550 10600
rect 25498 10548 25504 10600
rect 25556 10548 25562 10600
rect 26694 10548 26700 10600
rect 26752 10588 26758 10600
rect 26789 10591 26847 10597
rect 26789 10588 26801 10591
rect 26752 10560 26801 10588
rect 26752 10548 26758 10560
rect 26789 10557 26801 10560
rect 26835 10557 26847 10591
rect 26896 10588 26924 10628
rect 26973 10625 26985 10659
rect 27019 10625 27031 10659
rect 26973 10619 27031 10625
rect 27154 10616 27160 10668
rect 27212 10616 27218 10668
rect 28000 10665 28028 10696
rect 28166 10684 28172 10696
rect 28224 10684 28230 10736
rect 28258 10684 28264 10736
rect 28316 10724 28322 10736
rect 28316 10696 28488 10724
rect 28316 10684 28322 10696
rect 27985 10659 28043 10665
rect 27985 10625 27997 10659
rect 28031 10625 28043 10659
rect 27985 10619 28043 10625
rect 28074 10616 28080 10668
rect 28132 10616 28138 10668
rect 28460 10665 28488 10696
rect 30466 10684 30472 10736
rect 30524 10684 30530 10736
rect 31018 10684 31024 10736
rect 31076 10684 31082 10736
rect 31478 10684 31484 10736
rect 31536 10684 31542 10736
rect 32674 10684 32680 10736
rect 32732 10724 32738 10736
rect 33410 10724 33416 10736
rect 32732 10696 33416 10724
rect 32732 10684 32738 10696
rect 33410 10684 33416 10696
rect 33468 10684 33474 10736
rect 34698 10684 34704 10736
rect 34756 10724 34762 10736
rect 34793 10727 34851 10733
rect 34793 10724 34805 10727
rect 34756 10696 34805 10724
rect 34756 10684 34762 10696
rect 34793 10693 34805 10696
rect 34839 10693 34851 10727
rect 35084 10724 35112 10764
rect 35158 10752 35164 10804
rect 35216 10752 35222 10804
rect 35434 10752 35440 10804
rect 35492 10752 35498 10804
rect 35894 10752 35900 10804
rect 35952 10792 35958 10804
rect 35989 10795 36047 10801
rect 35989 10792 36001 10795
rect 35952 10764 36001 10792
rect 35952 10752 35958 10764
rect 35989 10761 36001 10764
rect 36035 10761 36047 10795
rect 35989 10755 36047 10761
rect 36814 10752 36820 10804
rect 36872 10752 36878 10804
rect 35452 10724 35480 10752
rect 35084 10696 35480 10724
rect 34793 10687 34851 10693
rect 28445 10659 28503 10665
rect 28445 10625 28457 10659
rect 28491 10625 28503 10659
rect 28445 10619 28503 10625
rect 28994 10616 29000 10668
rect 29052 10656 29058 10668
rect 29457 10659 29515 10665
rect 29457 10656 29469 10659
rect 29052 10628 29469 10656
rect 29052 10616 29058 10628
rect 29457 10625 29469 10628
rect 29503 10625 29515 10659
rect 29457 10619 29515 10625
rect 27172 10588 27200 10616
rect 26896 10560 27200 10588
rect 29733 10591 29791 10597
rect 26789 10551 26847 10557
rect 29733 10557 29745 10591
rect 29779 10588 29791 10591
rect 31036 10588 31064 10684
rect 36262 10656 36268 10668
rect 36004 10628 36268 10656
rect 36004 10600 36032 10628
rect 36262 10616 36268 10628
rect 36320 10656 36326 10668
rect 36725 10659 36783 10665
rect 36725 10656 36737 10659
rect 36320 10628 36737 10656
rect 36320 10616 36326 10628
rect 36725 10625 36737 10628
rect 36771 10625 36783 10659
rect 36725 10619 36783 10625
rect 29779 10560 31064 10588
rect 29779 10557 29791 10560
rect 29733 10551 29791 10557
rect 35986 10548 35992 10600
rect 36044 10548 36050 10600
rect 36538 10548 36544 10600
rect 36596 10548 36602 10600
rect 25516 10520 25544 10548
rect 19484 10492 19840 10520
rect 24504 10492 25544 10520
rect 19484 10480 19490 10492
rect 17788 10424 18920 10452
rect 18966 10412 18972 10464
rect 19024 10412 19030 10464
rect 20070 10412 20076 10464
rect 20128 10412 20134 10464
rect 22373 10455 22431 10461
rect 22373 10421 22385 10455
rect 22419 10452 22431 10455
rect 23014 10452 23020 10464
rect 22419 10424 23020 10452
rect 22419 10421 22431 10424
rect 22373 10415 22431 10421
rect 23014 10412 23020 10424
rect 23072 10412 23078 10464
rect 24504 10461 24532 10492
rect 32858 10480 32864 10532
rect 32916 10520 32922 10532
rect 33045 10523 33103 10529
rect 33045 10520 33057 10523
rect 32916 10492 33057 10520
rect 32916 10480 32922 10492
rect 33045 10489 33057 10492
rect 33091 10520 33103 10523
rect 34422 10520 34428 10532
rect 33091 10492 34428 10520
rect 33091 10489 33103 10492
rect 33045 10483 33103 10489
rect 34422 10480 34428 10492
rect 34480 10520 34486 10532
rect 36556 10520 36584 10548
rect 34480 10492 36584 10520
rect 34480 10480 34486 10492
rect 24489 10455 24547 10461
rect 24489 10421 24501 10455
rect 24535 10421 24547 10455
rect 24489 10415 24547 10421
rect 24854 10412 24860 10464
rect 24912 10412 24918 10464
rect 25590 10412 25596 10464
rect 25648 10412 25654 10464
rect 26053 10455 26111 10461
rect 26053 10421 26065 10455
rect 26099 10452 26111 10455
rect 26326 10452 26332 10464
rect 26099 10424 26332 10452
rect 26099 10421 26111 10424
rect 26053 10415 26111 10421
rect 26326 10412 26332 10424
rect 26384 10412 26390 10464
rect 26418 10412 26424 10464
rect 26476 10412 26482 10464
rect 27798 10412 27804 10464
rect 27856 10412 27862 10464
rect 34790 10412 34796 10464
rect 34848 10452 34854 10464
rect 34977 10455 35035 10461
rect 34977 10452 34989 10455
rect 34848 10424 34989 10452
rect 34848 10412 34854 10424
rect 34977 10421 34989 10424
rect 35023 10421 35035 10455
rect 34977 10415 35035 10421
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 20162 10248 20168 10260
rect 17276 10220 20168 10248
rect 17276 10208 17282 10220
rect 18233 10183 18291 10189
rect 18233 10149 18245 10183
rect 18279 10149 18291 10183
rect 18233 10143 18291 10149
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10112 14979 10115
rect 18248 10112 18276 10143
rect 14967 10084 18276 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 16390 10044 16396 10056
rect 16054 10016 16396 10044
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 16758 10004 16764 10056
rect 16816 10044 16822 10056
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16816 10016 16865 10044
rect 16816 10004 16822 10016
rect 16853 10013 16865 10016
rect 16899 10044 16911 10047
rect 17494 10044 17500 10056
rect 16899 10016 17500 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10044 17647 10047
rect 17678 10044 17684 10056
rect 17635 10016 17684 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 17604 9976 17632 10007
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10044 18475 10047
rect 18690 10044 18696 10056
rect 18463 10016 18696 10044
rect 18463 10013 18475 10016
rect 18417 10007 18475 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 18800 10053 18828 10220
rect 20162 10208 20168 10220
rect 20220 10248 20226 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 20220 10220 20269 10248
rect 20220 10208 20226 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 20717 10251 20775 10257
rect 20717 10217 20729 10251
rect 20763 10248 20775 10251
rect 20806 10248 20812 10260
rect 20763 10220 20812 10248
rect 20763 10217 20775 10220
rect 20717 10211 20775 10217
rect 20806 10208 20812 10220
rect 20864 10208 20870 10260
rect 23658 10208 23664 10260
rect 23716 10208 23722 10260
rect 24486 10208 24492 10260
rect 24544 10208 24550 10260
rect 24854 10208 24860 10260
rect 24912 10208 24918 10260
rect 25222 10208 25228 10260
rect 25280 10208 25286 10260
rect 25590 10208 25596 10260
rect 25648 10208 25654 10260
rect 26510 10208 26516 10260
rect 26568 10208 26574 10260
rect 30466 10208 30472 10260
rect 30524 10208 30530 10260
rect 31386 10208 31392 10260
rect 31444 10248 31450 10260
rect 32674 10248 32680 10260
rect 31444 10220 32680 10248
rect 31444 10208 31450 10220
rect 32674 10208 32680 10220
rect 32732 10248 32738 10260
rect 33778 10248 33784 10260
rect 32732 10220 33784 10248
rect 32732 10208 32738 10220
rect 33778 10208 33784 10220
rect 33836 10248 33842 10260
rect 34238 10248 34244 10260
rect 33836 10220 34244 10248
rect 33836 10208 33842 10220
rect 34238 10208 34244 10220
rect 34296 10208 34302 10260
rect 19334 10140 19340 10192
rect 19392 10140 19398 10192
rect 19352 10112 19380 10140
rect 19978 10112 19984 10124
rect 19260 10084 19380 10112
rect 19444 10084 19984 10112
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10013 18843 10047
rect 18785 10007 18843 10013
rect 18874 10004 18880 10056
rect 18932 10004 18938 10056
rect 19058 10004 19064 10056
rect 19116 10004 19122 10056
rect 19260 10044 19288 10084
rect 19444 10053 19472 10084
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 20070 10072 20076 10124
rect 20128 10072 20134 10124
rect 20441 10115 20499 10121
rect 20441 10081 20453 10115
rect 20487 10112 20499 10115
rect 23014 10112 23020 10124
rect 20487 10084 23020 10112
rect 20487 10081 20499 10084
rect 20441 10075 20499 10081
rect 23014 10072 23020 10084
rect 23072 10072 23078 10124
rect 24872 10112 24900 10208
rect 25501 10183 25559 10189
rect 25501 10149 25513 10183
rect 25547 10180 25559 10183
rect 25608 10180 25636 10208
rect 25547 10152 25636 10180
rect 25547 10149 25559 10152
rect 25501 10143 25559 10149
rect 31404 10121 31432 10208
rect 33134 10180 33140 10192
rect 32324 10152 33140 10180
rect 25133 10115 25191 10121
rect 25133 10112 25145 10115
rect 24872 10084 25145 10112
rect 25133 10081 25145 10084
rect 25179 10081 25191 10115
rect 31389 10115 31447 10121
rect 25133 10075 25191 10081
rect 25516 10084 26188 10112
rect 19337 10047 19395 10053
rect 19337 10044 19349 10047
rect 19260 10016 19349 10044
rect 19337 10013 19349 10016
rect 19383 10013 19395 10047
rect 19337 10007 19395 10013
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10013 19579 10047
rect 20088 10044 20116 10072
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 20088 10016 20269 10044
rect 19521 10007 19579 10013
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 24673 10047 24731 10053
rect 24673 10013 24685 10047
rect 24719 10044 24731 10047
rect 25314 10044 25320 10056
rect 24719 10016 25320 10044
rect 24719 10013 24731 10016
rect 24673 10007 24731 10013
rect 16408 9948 17632 9976
rect 18141 9979 18199 9985
rect 16408 9917 16436 9948
rect 18141 9945 18153 9979
rect 18187 9976 18199 9979
rect 18509 9979 18567 9985
rect 18509 9976 18521 9979
rect 18187 9948 18521 9976
rect 18187 9945 18199 9948
rect 18141 9939 18199 9945
rect 18509 9945 18521 9948
rect 18555 9945 18567 9979
rect 18509 9939 18567 9945
rect 18601 9979 18659 9985
rect 18601 9945 18613 9979
rect 18647 9976 18659 9979
rect 18969 9979 19027 9985
rect 18969 9976 18981 9979
rect 18647 9948 18981 9976
rect 18647 9945 18659 9948
rect 18601 9939 18659 9945
rect 18969 9945 18981 9948
rect 19015 9945 19027 9979
rect 19536 9976 19564 10007
rect 18969 9939 19027 9945
rect 19352 9948 19564 9976
rect 19705 9979 19763 9985
rect 19352 9920 19380 9948
rect 19705 9945 19717 9979
rect 19751 9976 19763 9979
rect 20548 9976 20576 10007
rect 19751 9948 20576 9976
rect 23584 9976 23612 10007
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 25409 10047 25467 10053
rect 25409 10013 25421 10047
rect 25455 10013 25467 10047
rect 25409 10007 25467 10013
rect 23842 9976 23848 9988
rect 23584 9948 23848 9976
rect 19751 9945 19763 9948
rect 19705 9939 19763 9945
rect 23842 9936 23848 9948
rect 23900 9936 23906 9988
rect 24765 9979 24823 9985
rect 24765 9945 24777 9979
rect 24811 9945 24823 9979
rect 24765 9939 24823 9945
rect 16393 9911 16451 9917
rect 16393 9877 16405 9911
rect 16439 9877 16451 9911
rect 16393 9871 16451 9877
rect 17402 9868 17408 9920
rect 17460 9868 17466 9920
rect 19334 9868 19340 9920
rect 19392 9868 19398 9920
rect 24780 9908 24808 9939
rect 24854 9936 24860 9988
rect 24912 9936 24918 9988
rect 24946 9936 24952 9988
rect 25004 9985 25010 9988
rect 25004 9979 25033 9985
rect 25021 9945 25033 9979
rect 25004 9939 25033 9945
rect 25004 9936 25010 9939
rect 25130 9936 25136 9988
rect 25188 9976 25194 9988
rect 25424 9976 25452 10007
rect 25516 9988 25544 10084
rect 25590 10004 25596 10056
rect 25648 10004 25654 10056
rect 25682 10004 25688 10056
rect 25740 10004 25746 10056
rect 25774 10004 25780 10056
rect 25832 10004 25838 10056
rect 25869 10047 25927 10053
rect 25869 10013 25881 10047
rect 25915 10044 25927 10047
rect 26050 10044 26056 10056
rect 25915 10016 26056 10044
rect 25915 10013 25927 10016
rect 25869 10007 25927 10013
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 26160 10053 26188 10084
rect 31389 10081 31401 10115
rect 31435 10081 31447 10115
rect 31389 10075 31447 10081
rect 31570 10072 31576 10124
rect 31628 10112 31634 10124
rect 31938 10112 31944 10124
rect 31628 10084 31944 10112
rect 31628 10072 31634 10084
rect 31938 10072 31944 10084
rect 31996 10112 32002 10124
rect 32324 10112 32352 10152
rect 33134 10140 33140 10152
rect 33192 10140 33198 10192
rect 33410 10140 33416 10192
rect 33468 10180 33474 10192
rect 33468 10152 33916 10180
rect 33468 10140 33474 10152
rect 31996 10084 32352 10112
rect 31996 10072 32002 10084
rect 26145 10047 26203 10053
rect 26145 10013 26157 10047
rect 26191 10013 26203 10047
rect 26145 10007 26203 10013
rect 26694 10004 26700 10056
rect 26752 10004 26758 10056
rect 29270 10004 29276 10056
rect 29328 10044 29334 10056
rect 29733 10047 29791 10053
rect 29733 10044 29745 10047
rect 29328 10016 29745 10044
rect 29328 10004 29334 10016
rect 29733 10013 29745 10016
rect 29779 10044 29791 10047
rect 30282 10044 30288 10056
rect 29779 10016 30288 10044
rect 29779 10013 29791 10016
rect 29733 10007 29791 10013
rect 30282 10004 30288 10016
rect 30340 10044 30346 10056
rect 30377 10047 30435 10053
rect 30377 10044 30389 10047
rect 30340 10016 30389 10044
rect 30340 10004 30346 10016
rect 30377 10013 30389 10016
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 31110 10004 31116 10056
rect 31168 10044 31174 10056
rect 32324 10053 32352 10084
rect 32398 10072 32404 10124
rect 32456 10112 32462 10124
rect 32677 10115 32735 10121
rect 32677 10112 32689 10115
rect 32456 10084 32689 10112
rect 32456 10072 32462 10084
rect 32677 10081 32689 10084
rect 32723 10081 32735 10115
rect 33318 10112 33324 10124
rect 32677 10075 32735 10081
rect 32876 10084 33324 10112
rect 32876 10056 32904 10084
rect 33318 10072 33324 10084
rect 33376 10112 33382 10124
rect 33888 10121 33916 10152
rect 33781 10115 33839 10121
rect 33781 10112 33793 10115
rect 33376 10084 33793 10112
rect 33376 10072 33382 10084
rect 33781 10081 33793 10084
rect 33827 10081 33839 10115
rect 33781 10075 33839 10081
rect 33873 10115 33931 10121
rect 33873 10081 33885 10115
rect 33919 10112 33931 10115
rect 35250 10112 35256 10124
rect 33919 10084 35256 10112
rect 33919 10081 33931 10084
rect 33873 10075 33931 10081
rect 35250 10072 35256 10084
rect 35308 10072 35314 10124
rect 31297 10047 31355 10053
rect 31297 10044 31309 10047
rect 31168 10016 31309 10044
rect 31168 10004 31174 10016
rect 31297 10013 31309 10016
rect 31343 10013 31355 10047
rect 31297 10007 31355 10013
rect 32309 10047 32367 10053
rect 32309 10013 32321 10047
rect 32355 10013 32367 10047
rect 32309 10007 32367 10013
rect 32585 10047 32643 10053
rect 32585 10013 32597 10047
rect 32631 10044 32643 10047
rect 32858 10044 32864 10056
rect 32631 10016 32864 10044
rect 32631 10013 32643 10016
rect 32585 10007 32643 10013
rect 32858 10004 32864 10016
rect 32916 10004 32922 10056
rect 33134 10004 33140 10056
rect 33192 10044 33198 10056
rect 33597 10047 33655 10053
rect 33597 10044 33609 10047
rect 33192 10016 33609 10044
rect 33192 10004 33198 10016
rect 33597 10013 33609 10016
rect 33643 10013 33655 10047
rect 33597 10007 33655 10013
rect 33686 10004 33692 10056
rect 33744 10004 33750 10056
rect 34790 10004 34796 10056
rect 34848 10004 34854 10056
rect 35437 10047 35495 10053
rect 35437 10013 35449 10047
rect 35483 10013 35495 10047
rect 35437 10007 35495 10013
rect 25188 9948 25452 9976
rect 25188 9936 25194 9948
rect 25498 9936 25504 9988
rect 25556 9936 25562 9988
rect 25792 9976 25820 10004
rect 25961 9979 26019 9985
rect 25961 9976 25973 9979
rect 25792 9948 25973 9976
rect 25961 9945 25973 9948
rect 26007 9945 26019 9979
rect 25961 9939 26019 9945
rect 32493 9979 32551 9985
rect 32493 9945 32505 9979
rect 32539 9976 32551 9979
rect 33045 9979 33103 9985
rect 33045 9976 33057 9979
rect 32539 9948 33057 9976
rect 32539 9945 32551 9948
rect 32493 9939 32551 9945
rect 33045 9945 33057 9948
rect 33091 9976 33103 9979
rect 33704 9976 33732 10004
rect 33091 9948 33732 9976
rect 34808 9976 34836 10004
rect 35452 9976 35480 10007
rect 68462 10004 68468 10056
rect 68520 10004 68526 10056
rect 34808 9948 35480 9976
rect 33091 9945 33103 9948
rect 33045 9939 33103 9945
rect 26326 9908 26332 9920
rect 24780 9880 26332 9908
rect 26326 9868 26332 9880
rect 26384 9868 26390 9920
rect 28810 9868 28816 9920
rect 28868 9908 28874 9920
rect 29641 9911 29699 9917
rect 29641 9908 29653 9911
rect 28868 9880 29653 9908
rect 28868 9868 28874 9880
rect 29641 9877 29653 9880
rect 29687 9877 29699 9911
rect 29641 9871 29699 9877
rect 30926 9868 30932 9920
rect 30984 9868 30990 9920
rect 32582 9868 32588 9920
rect 32640 9868 32646 9920
rect 33410 9868 33416 9920
rect 33468 9868 33474 9920
rect 34698 9868 34704 9920
rect 34756 9868 34762 9920
rect 35526 9868 35532 9920
rect 35584 9868 35590 9920
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 17126 9664 17132 9716
rect 17184 9664 17190 9716
rect 17494 9664 17500 9716
rect 17552 9704 17558 9716
rect 17552 9676 17908 9704
rect 17552 9664 17558 9676
rect 15930 9596 15936 9648
rect 15988 9596 15994 9648
rect 17144 9636 17172 9664
rect 17880 9636 17908 9676
rect 18064 9676 19012 9704
rect 18064 9636 18092 9676
rect 17144 9608 17816 9636
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 14921 9503 14979 9509
rect 14921 9469 14933 9503
rect 14967 9500 14979 9503
rect 16669 9503 16727 9509
rect 16669 9500 16681 9503
rect 14967 9472 16681 9500
rect 14967 9469 14979 9472
rect 14921 9463 14979 9469
rect 16669 9469 16681 9472
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 16758 9460 16764 9512
rect 16816 9460 16822 9512
rect 16868 9500 16896 9531
rect 16942 9528 16948 9580
rect 17000 9528 17006 9580
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 17126 9528 17132 9580
rect 17184 9577 17190 9580
rect 17184 9571 17213 9577
rect 17201 9537 17213 9571
rect 17184 9531 17213 9537
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9568 17371 9571
rect 17402 9568 17408 9580
rect 17359 9540 17408 9568
rect 17359 9537 17371 9540
rect 17313 9531 17371 9537
rect 17184 9528 17190 9531
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 16868 9472 17448 9500
rect 14660 9364 14688 9460
rect 16393 9435 16451 9441
rect 16393 9401 16405 9435
rect 16439 9432 16451 9435
rect 16776 9432 16804 9460
rect 17420 9441 17448 9472
rect 16439 9404 16804 9432
rect 17405 9435 17463 9441
rect 16439 9401 16451 9404
rect 16393 9395 16451 9401
rect 17405 9401 17417 9435
rect 17451 9401 17463 9435
rect 17405 9395 17463 9401
rect 15562 9364 15568 9376
rect 14660 9336 15568 9364
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 17512 9364 17540 9608
rect 17586 9528 17592 9580
rect 17644 9528 17650 9580
rect 17788 9577 17816 9608
rect 17880 9608 18092 9636
rect 17880 9577 17908 9608
rect 18138 9596 18144 9648
rect 18196 9596 18202 9648
rect 18874 9645 18880 9648
rect 18845 9639 18880 9645
rect 18845 9636 18857 9639
rect 18248 9608 18857 9636
rect 17773 9571 17831 9577
rect 17773 9537 17785 9571
rect 17819 9537 17831 9571
rect 17773 9531 17831 9537
rect 17865 9571 17923 9577
rect 17865 9537 17877 9571
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18248 9568 18276 9608
rect 18845 9605 18857 9608
rect 18845 9599 18880 9605
rect 18874 9596 18880 9599
rect 18932 9596 18938 9648
rect 18984 9636 19012 9676
rect 23014 9664 23020 9716
rect 23072 9664 23078 9716
rect 24213 9707 24271 9713
rect 24213 9673 24225 9707
rect 24259 9704 24271 9707
rect 24946 9704 24952 9716
rect 24259 9676 24952 9704
rect 24259 9673 24271 9676
rect 24213 9667 24271 9673
rect 24946 9664 24952 9676
rect 25004 9704 25010 9716
rect 25222 9704 25228 9716
rect 25004 9676 25228 9704
rect 25004 9664 25010 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 25501 9707 25559 9713
rect 25501 9673 25513 9707
rect 25547 9704 25559 9707
rect 25682 9704 25688 9716
rect 25547 9676 25688 9704
rect 25547 9673 25559 9676
rect 25501 9667 25559 9673
rect 25682 9664 25688 9676
rect 25740 9664 25746 9716
rect 26145 9707 26203 9713
rect 26145 9673 26157 9707
rect 26191 9704 26203 9707
rect 26694 9704 26700 9716
rect 26191 9676 26700 9704
rect 26191 9673 26203 9676
rect 26145 9667 26203 9673
rect 26694 9664 26700 9676
rect 26752 9664 26758 9716
rect 27798 9664 27804 9716
rect 27856 9704 27862 9716
rect 27856 9676 29224 9704
rect 27856 9664 27862 9676
rect 19061 9639 19119 9645
rect 19061 9636 19073 9639
rect 18984 9608 19073 9636
rect 19061 9605 19073 9608
rect 19107 9636 19119 9639
rect 19426 9636 19432 9648
rect 19107 9608 19432 9636
rect 19107 9605 19119 9608
rect 19061 9599 19119 9605
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 20254 9596 20260 9648
rect 20312 9636 20318 9648
rect 20349 9639 20407 9645
rect 20349 9636 20361 9639
rect 20312 9608 20361 9636
rect 20312 9596 20318 9608
rect 20349 9605 20361 9608
rect 20395 9605 20407 9639
rect 20349 9599 20407 9605
rect 21266 9596 21272 9648
rect 21324 9636 21330 9648
rect 21913 9639 21971 9645
rect 21913 9636 21925 9639
rect 21324 9608 21925 9636
rect 21324 9596 21330 9608
rect 21913 9605 21925 9608
rect 21959 9605 21971 9639
rect 21913 9599 21971 9605
rect 24121 9639 24179 9645
rect 24121 9605 24133 9639
rect 24167 9636 24179 9639
rect 26234 9636 26240 9648
rect 24167 9608 26240 9636
rect 24167 9605 24179 9608
rect 24121 9599 24179 9605
rect 26234 9596 26240 9608
rect 26292 9636 26298 9648
rect 26418 9636 26424 9648
rect 26292 9608 26424 9636
rect 26292 9596 26298 9608
rect 26418 9596 26424 9608
rect 26476 9596 26482 9648
rect 26789 9639 26847 9645
rect 26789 9605 26801 9639
rect 26835 9636 26847 9639
rect 26835 9608 27200 9636
rect 26835 9605 26847 9608
rect 26789 9599 26847 9605
rect 27172 9580 27200 9608
rect 28810 9596 28816 9648
rect 28868 9596 28874 9648
rect 29196 9636 29224 9676
rect 31110 9664 31116 9716
rect 31168 9704 31174 9716
rect 31168 9676 32352 9704
rect 31168 9664 31174 9676
rect 29196 9608 29408 9636
rect 18012 9540 18276 9568
rect 18325 9571 18383 9577
rect 18012 9528 18018 9540
rect 18325 9537 18337 9571
rect 18371 9568 18383 9571
rect 18966 9568 18972 9580
rect 18371 9540 18972 9568
rect 18371 9537 18383 9540
rect 18325 9531 18383 9537
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 20530 9528 20536 9580
rect 20588 9528 20594 9580
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 20732 9540 21189 9568
rect 17678 9460 17684 9512
rect 17736 9500 17742 9512
rect 17736 9472 18552 9500
rect 17736 9460 17742 9472
rect 18524 9444 18552 9472
rect 18598 9460 18604 9512
rect 18656 9509 18662 9512
rect 18656 9500 18665 9509
rect 18656 9472 18701 9500
rect 18656 9463 18665 9472
rect 18656 9460 18662 9463
rect 18506 9392 18512 9444
rect 18564 9392 18570 9444
rect 18693 9435 18751 9441
rect 18693 9401 18705 9435
rect 18739 9432 18751 9435
rect 18739 9404 19380 9432
rect 18739 9401 18751 9404
rect 18693 9395 18751 9401
rect 19352 9376 19380 9404
rect 20732 9376 20760 9540
rect 21177 9537 21189 9540
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 21361 9571 21419 9577
rect 21361 9537 21373 9571
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 21082 9460 21088 9512
rect 21140 9500 21146 9512
rect 21376 9500 21404 9531
rect 21542 9528 21548 9580
rect 21600 9528 21606 9580
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 22066 9540 22661 9568
rect 21140 9472 21404 9500
rect 21140 9460 21146 9472
rect 21910 9460 21916 9512
rect 21968 9500 21974 9512
rect 22066 9500 22094 9540
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 22833 9571 22891 9577
rect 22833 9537 22845 9571
rect 22879 9537 22891 9571
rect 22833 9531 22891 9537
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9568 23351 9571
rect 23339 9540 23796 9568
rect 23339 9537 23351 9540
rect 23293 9531 23351 9537
rect 22465 9503 22523 9509
rect 22465 9500 22477 9503
rect 21968 9472 22094 9500
rect 22296 9472 22477 9500
rect 21968 9460 21974 9472
rect 20898 9392 20904 9444
rect 20956 9432 20962 9444
rect 21928 9432 21956 9460
rect 20956 9404 21956 9432
rect 20956 9392 20962 9404
rect 22296 9376 22324 9472
rect 22465 9469 22477 9472
rect 22511 9500 22523 9503
rect 22848 9500 22876 9531
rect 22511 9472 22876 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 23768 9441 23796 9540
rect 24762 9528 24768 9580
rect 24820 9528 24826 9580
rect 24946 9568 24952 9580
rect 24918 9528 24952 9568
rect 25004 9568 25010 9580
rect 25774 9568 25780 9580
rect 25004 9540 25780 9568
rect 25004 9528 25010 9540
rect 25774 9528 25780 9540
rect 25832 9528 25838 9580
rect 25866 9528 25872 9580
rect 25924 9568 25930 9580
rect 26329 9571 26387 9577
rect 26329 9568 26341 9571
rect 25924 9540 26341 9568
rect 25924 9528 25930 9540
rect 26329 9537 26341 9540
rect 26375 9537 26387 9571
rect 26329 9531 26387 9537
rect 27154 9528 27160 9580
rect 27212 9528 27218 9580
rect 29380 9577 29408 9608
rect 31202 9596 31208 9648
rect 31260 9596 31266 9648
rect 31938 9596 31944 9648
rect 31996 9596 32002 9648
rect 29365 9571 29423 9577
rect 29365 9537 29377 9571
rect 29411 9537 29423 9571
rect 29365 9531 29423 9537
rect 29546 9528 29552 9580
rect 29604 9528 29610 9580
rect 24394 9460 24400 9512
rect 24452 9500 24458 9512
rect 24918 9500 24946 9528
rect 25225 9503 25283 9509
rect 25225 9500 25237 9503
rect 24452 9472 24946 9500
rect 25056 9472 25237 9500
rect 24452 9460 24458 9472
rect 23753 9435 23811 9441
rect 23753 9401 23765 9435
rect 23799 9401 23811 9435
rect 25056 9432 25084 9472
rect 25225 9469 25237 9472
rect 25271 9500 25283 9503
rect 25958 9500 25964 9512
rect 25271 9472 25964 9500
rect 25271 9469 25283 9472
rect 25225 9463 25283 9469
rect 25958 9460 25964 9472
rect 26016 9460 26022 9512
rect 26418 9460 26424 9512
rect 26476 9460 26482 9512
rect 27525 9503 27583 9509
rect 27525 9469 27537 9503
rect 27571 9500 27583 9503
rect 27571 9472 27660 9500
rect 27571 9469 27583 9472
rect 27525 9463 27583 9469
rect 23753 9395 23811 9401
rect 24688 9404 25084 9432
rect 25133 9435 25191 9441
rect 24688 9376 24716 9404
rect 25133 9401 25145 9435
rect 25179 9432 25191 9435
rect 25179 9404 26556 9432
rect 25179 9401 25191 9404
rect 25133 9395 25191 9401
rect 26528 9376 26556 9404
rect 18598 9364 18604 9376
rect 17512 9336 18604 9364
rect 18598 9324 18604 9336
rect 18656 9364 18662 9376
rect 18877 9367 18935 9373
rect 18877 9364 18889 9367
rect 18656 9336 18889 9364
rect 18656 9324 18662 9336
rect 18877 9333 18889 9336
rect 18923 9333 18935 9367
rect 18877 9327 18935 9333
rect 19334 9324 19340 9376
rect 19392 9324 19398 9376
rect 20714 9324 20720 9376
rect 20772 9324 20778 9376
rect 20990 9324 20996 9376
rect 21048 9324 21054 9376
rect 22278 9324 22284 9376
rect 22336 9324 22342 9376
rect 23106 9324 23112 9376
rect 23164 9324 23170 9376
rect 24670 9324 24676 9376
rect 24728 9324 24734 9376
rect 25038 9324 25044 9376
rect 25096 9324 25102 9376
rect 26326 9324 26332 9376
rect 26384 9324 26390 9376
rect 26510 9324 26516 9376
rect 26568 9324 26574 9376
rect 27430 9324 27436 9376
rect 27488 9364 27494 9376
rect 27632 9364 27660 9472
rect 27798 9460 27804 9512
rect 27856 9460 27862 9512
rect 28994 9460 29000 9512
rect 29052 9500 29058 9512
rect 29917 9503 29975 9509
rect 29917 9500 29929 9503
rect 29052 9472 29929 9500
rect 29052 9460 29058 9472
rect 29917 9469 29929 9472
rect 29963 9469 29975 9503
rect 29917 9463 29975 9469
rect 30193 9503 30251 9509
rect 30193 9469 30205 9503
rect 30239 9500 30251 9503
rect 30742 9500 30748 9512
rect 30239 9472 30748 9500
rect 30239 9469 30251 9472
rect 30193 9463 30251 9469
rect 30742 9460 30748 9472
rect 30800 9460 30806 9512
rect 32324 9500 32352 9676
rect 32398 9664 32404 9716
rect 32456 9664 32462 9716
rect 32582 9704 32588 9716
rect 32508 9676 32588 9704
rect 32416 9577 32444 9664
rect 32508 9645 32536 9676
rect 32582 9664 32588 9676
rect 32640 9664 32646 9716
rect 32858 9664 32864 9716
rect 32916 9664 32922 9716
rect 33410 9704 33416 9716
rect 33336 9676 33416 9704
rect 32493 9639 32551 9645
rect 32493 9605 32505 9639
rect 32539 9605 32551 9639
rect 32493 9599 32551 9605
rect 32674 9596 32680 9648
rect 32732 9645 32738 9648
rect 32732 9639 32761 9645
rect 32749 9605 32761 9639
rect 32732 9599 32761 9605
rect 32732 9596 32738 9599
rect 32401 9571 32459 9577
rect 32401 9537 32413 9571
rect 32447 9537 32459 9571
rect 32401 9531 32459 9537
rect 32582 9528 32588 9580
rect 32640 9528 32646 9580
rect 32876 9577 32904 9664
rect 32861 9571 32919 9577
rect 32861 9537 32873 9571
rect 32907 9537 32919 9571
rect 33336 9574 33364 9676
rect 33410 9664 33416 9676
rect 33468 9664 33474 9716
rect 35250 9664 35256 9716
rect 35308 9704 35314 9716
rect 35713 9707 35771 9713
rect 35713 9704 35725 9707
rect 35308 9676 35725 9704
rect 35308 9664 35314 9676
rect 35713 9673 35725 9676
rect 35759 9673 35771 9707
rect 35713 9667 35771 9673
rect 33594 9596 33600 9648
rect 33652 9645 33658 9648
rect 33652 9639 33668 9645
rect 33656 9605 33668 9639
rect 33652 9599 33668 9605
rect 33652 9596 33658 9599
rect 34238 9596 34244 9648
rect 34296 9596 34302 9648
rect 35897 9639 35955 9645
rect 35897 9636 35909 9639
rect 35466 9608 35909 9636
rect 35897 9605 35909 9608
rect 35943 9605 35955 9639
rect 35897 9599 35955 9605
rect 33414 9577 33472 9583
rect 33414 9574 33426 9577
rect 33336 9546 33426 9574
rect 33414 9543 33426 9546
rect 33460 9543 33472 9577
rect 33414 9537 33472 9543
rect 33506 9571 33564 9577
rect 33506 9537 33518 9571
rect 33552 9568 33564 9571
rect 33715 9571 33773 9577
rect 33552 9540 33640 9568
rect 33552 9537 33564 9540
rect 32861 9531 32919 9537
rect 33506 9531 33564 9537
rect 32600 9500 32628 9528
rect 32324 9472 32628 9500
rect 29012 9364 29040 9460
rect 29273 9435 29331 9441
rect 29273 9401 29285 9435
rect 29319 9432 29331 9435
rect 29319 9404 29868 9432
rect 29319 9401 29331 9404
rect 29273 9395 29331 9401
rect 29840 9376 29868 9404
rect 27488 9336 29040 9364
rect 27488 9324 27494 9336
rect 29730 9324 29736 9376
rect 29788 9324 29794 9376
rect 29822 9324 29828 9376
rect 29880 9324 29886 9376
rect 32214 9324 32220 9376
rect 32272 9324 32278 9376
rect 33229 9367 33287 9373
rect 33229 9333 33241 9367
rect 33275 9364 33287 9367
rect 33410 9364 33416 9376
rect 33275 9336 33416 9364
rect 33275 9333 33287 9336
rect 33229 9327 33287 9333
rect 33410 9324 33416 9336
rect 33468 9324 33474 9376
rect 33612 9364 33640 9540
rect 33715 9537 33727 9571
rect 33761 9558 33773 9571
rect 33761 9537 33824 9558
rect 33715 9531 33824 9537
rect 33730 9530 33824 9531
rect 33796 9444 33824 9530
rect 33962 9528 33968 9580
rect 34020 9528 34026 9580
rect 35986 9528 35992 9580
rect 36044 9528 36050 9580
rect 33873 9503 33931 9509
rect 33873 9469 33885 9503
rect 33919 9500 33931 9503
rect 34698 9500 34704 9512
rect 33919 9472 34704 9500
rect 33919 9469 33931 9472
rect 33873 9463 33931 9469
rect 34698 9460 34704 9472
rect 34756 9460 34762 9512
rect 33778 9392 33784 9444
rect 33836 9392 33842 9444
rect 35526 9364 35532 9376
rect 33612 9336 35532 9364
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 15930 9120 15936 9172
rect 15988 9120 15994 9172
rect 16942 9120 16948 9172
rect 17000 9160 17006 9172
rect 17773 9163 17831 9169
rect 17773 9160 17785 9163
rect 17000 9132 17785 9160
rect 17000 9120 17006 9132
rect 17773 9129 17785 9132
rect 17819 9129 17831 9163
rect 17773 9123 17831 9129
rect 20070 9120 20076 9172
rect 20128 9160 20134 9172
rect 20257 9163 20315 9169
rect 20257 9160 20269 9163
rect 20128 9132 20269 9160
rect 20128 9120 20134 9132
rect 20257 9129 20269 9132
rect 20303 9129 20315 9163
rect 20257 9123 20315 9129
rect 20530 9120 20536 9172
rect 20588 9120 20594 9172
rect 20796 9163 20854 9169
rect 20796 9129 20808 9163
rect 20842 9160 20854 9163
rect 20990 9160 20996 9172
rect 20842 9132 20996 9160
rect 20842 9129 20854 9132
rect 20796 9123 20854 9129
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 22462 9160 22468 9172
rect 22066 9132 22468 9160
rect 17405 9095 17463 9101
rect 17405 9061 17417 9095
rect 17451 9092 17463 9095
rect 17954 9092 17960 9104
rect 17451 9064 17960 9092
rect 17451 9061 17463 9064
rect 17405 9055 17463 9061
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 18322 9052 18328 9104
rect 18380 9092 18386 9104
rect 19058 9092 19064 9104
rect 18380 9064 19064 9092
rect 18380 9052 18386 9064
rect 19058 9052 19064 9064
rect 19116 9092 19122 9104
rect 19981 9095 20039 9101
rect 19116 9064 19840 9092
rect 19116 9052 19122 9064
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 17678 9024 17684 9036
rect 17083 8996 17684 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 18693 9027 18751 9033
rect 18693 8993 18705 9027
rect 18739 9024 18751 9027
rect 18966 9024 18972 9036
rect 18739 8996 18972 9024
rect 18739 8993 18751 8996
rect 18693 8987 18751 8993
rect 18966 8984 18972 8996
rect 19024 9024 19030 9036
rect 19242 9024 19248 9036
rect 19024 8996 19248 9024
rect 19024 8984 19030 8996
rect 19242 8984 19248 8996
rect 19300 8984 19306 9036
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 16482 8956 16488 8968
rect 16071 8928 16488 8956
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 16482 8916 16488 8928
rect 16540 8956 16546 8968
rect 16758 8956 16764 8968
rect 16540 8928 16764 8956
rect 16540 8916 16546 8928
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8956 17279 8959
rect 17586 8956 17592 8968
rect 17267 8928 17592 8956
rect 17267 8925 17279 8928
rect 17221 8919 17279 8925
rect 17586 8916 17592 8928
rect 17644 8916 17650 8968
rect 19812 8965 19840 9064
rect 19981 9061 19993 9095
rect 20027 9092 20039 9095
rect 20548 9092 20576 9120
rect 20027 9064 20576 9092
rect 20027 9061 20039 9064
rect 19981 9055 20039 9061
rect 22066 9036 22094 9132
rect 22462 9120 22468 9132
rect 22520 9120 22526 9172
rect 24121 9163 24179 9169
rect 24121 9129 24133 9163
rect 24167 9160 24179 9163
rect 24394 9160 24400 9172
rect 24167 9132 24400 9160
rect 24167 9129 24179 9132
rect 24121 9123 24179 9129
rect 24394 9120 24400 9132
rect 24452 9120 24458 9172
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 24857 9163 24915 9169
rect 24857 9160 24869 9163
rect 24820 9132 24869 9160
rect 24820 9120 24826 9132
rect 24857 9129 24869 9132
rect 24903 9129 24915 9163
rect 24857 9123 24915 9129
rect 25501 9163 25559 9169
rect 25501 9129 25513 9163
rect 25547 9160 25559 9163
rect 25590 9160 25596 9172
rect 25547 9132 25596 9160
rect 25547 9129 25559 9132
rect 25501 9123 25559 9129
rect 25590 9120 25596 9132
rect 25648 9120 25654 9172
rect 25866 9120 25872 9172
rect 25924 9120 25930 9172
rect 26418 9120 26424 9172
rect 26476 9120 26482 9172
rect 26510 9120 26516 9172
rect 26568 9160 26574 9172
rect 26973 9163 27031 9169
rect 26568 9132 26832 9160
rect 26568 9120 26574 9132
rect 22278 9052 22284 9104
rect 22336 9052 22342 9104
rect 20533 9027 20591 9033
rect 20533 8993 20545 9027
rect 20579 9024 20591 9027
rect 22002 9024 22008 9036
rect 20579 8996 22008 9024
rect 20579 8993 20591 8996
rect 20533 8987 20591 8993
rect 22002 8984 22008 8996
rect 22060 9024 22094 9036
rect 22373 9027 22431 9033
rect 22373 9024 22385 9027
rect 22060 8996 22385 9024
rect 22060 8984 22066 8996
rect 22373 8993 22385 8996
rect 22419 8993 22431 9027
rect 22373 8987 22431 8993
rect 22649 9027 22707 9033
rect 22649 8993 22661 9027
rect 22695 9024 22707 9027
rect 23106 9024 23112 9036
rect 22695 8996 23112 9024
rect 22695 8993 22707 8996
rect 22649 8987 22707 8993
rect 23106 8984 23112 8996
rect 23164 8984 23170 9036
rect 25314 8984 25320 9036
rect 25372 8984 25378 9036
rect 25884 9024 25912 9120
rect 25700 8996 25912 9024
rect 25976 9064 26740 9092
rect 25700 8965 25728 8996
rect 25976 8968 26004 9064
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8925 18935 8959
rect 18877 8919 18935 8925
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8925 19855 8959
rect 19797 8919 19855 8925
rect 19981 8959 20039 8965
rect 19981 8925 19993 8959
rect 20027 8956 20039 8959
rect 25225 8959 25283 8965
rect 20027 8928 20392 8956
rect 20027 8925 20039 8928
rect 19981 8919 20039 8925
rect 17880 8888 17908 8919
rect 18892 8888 18920 8919
rect 17880 8860 18920 8888
rect 17126 8780 17132 8832
rect 17184 8820 17190 8832
rect 18690 8820 18696 8832
rect 17184 8792 18696 8820
rect 17184 8780 17190 8792
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 18892 8820 18920 8860
rect 19061 8891 19119 8897
rect 19061 8857 19073 8891
rect 19107 8888 19119 8891
rect 20225 8891 20283 8897
rect 20225 8888 20237 8891
rect 19107 8860 20237 8888
rect 19107 8857 19119 8860
rect 19061 8851 19119 8857
rect 19996 8832 20024 8860
rect 20225 8857 20237 8860
rect 20271 8857 20283 8891
rect 20225 8851 20283 8857
rect 19334 8820 19340 8832
rect 18892 8792 19340 8820
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 19978 8780 19984 8832
rect 20036 8780 20042 8832
rect 20073 8823 20131 8829
rect 20073 8789 20085 8823
rect 20119 8820 20131 8823
rect 20364 8820 20392 8928
rect 25225 8925 25237 8959
rect 25271 8956 25283 8959
rect 25685 8959 25743 8965
rect 25685 8956 25697 8959
rect 25271 8928 25697 8956
rect 25271 8925 25283 8928
rect 25225 8919 25283 8925
rect 25685 8925 25697 8928
rect 25731 8925 25743 8959
rect 25685 8919 25743 8925
rect 25777 8959 25835 8965
rect 25777 8925 25789 8959
rect 25823 8925 25835 8959
rect 25777 8919 25835 8925
rect 25869 8959 25927 8965
rect 25869 8925 25881 8959
rect 25915 8956 25927 8959
rect 25958 8956 25964 8968
rect 25915 8928 25964 8956
rect 25915 8925 25927 8928
rect 25869 8919 25927 8925
rect 20441 8891 20499 8897
rect 20441 8857 20453 8891
rect 20487 8888 20499 8891
rect 20898 8888 20904 8900
rect 20487 8860 20904 8888
rect 20487 8857 20499 8860
rect 20441 8851 20499 8857
rect 20898 8848 20904 8860
rect 20956 8848 20962 8900
rect 22646 8888 22652 8900
rect 22034 8860 22652 8888
rect 22646 8848 22652 8860
rect 22704 8848 22710 8900
rect 23658 8848 23664 8900
rect 23716 8848 23722 8900
rect 25792 8888 25820 8919
rect 25958 8916 25964 8928
rect 26016 8916 26022 8968
rect 26510 8916 26516 8968
rect 26568 8916 26574 8968
rect 26712 8965 26740 9064
rect 26605 8959 26663 8965
rect 26605 8925 26617 8959
rect 26651 8925 26663 8959
rect 26605 8919 26663 8925
rect 26697 8959 26755 8965
rect 26697 8925 26709 8959
rect 26743 8925 26755 8959
rect 26804 8956 26832 9132
rect 26973 9129 26985 9163
rect 27019 9129 27031 9163
rect 26973 9123 27031 9129
rect 26988 9092 27016 9123
rect 27154 9120 27160 9172
rect 27212 9160 27218 9172
rect 27525 9163 27583 9169
rect 27525 9160 27537 9163
rect 27212 9132 27537 9160
rect 27212 9120 27218 9132
rect 27525 9129 27537 9132
rect 27571 9129 27583 9163
rect 27525 9123 27583 9129
rect 27798 9120 27804 9172
rect 27856 9120 27862 9172
rect 27908 9132 29684 9160
rect 27908 9092 27936 9132
rect 29656 9104 29684 9132
rect 29730 9120 29736 9172
rect 29788 9120 29794 9172
rect 31113 9163 31171 9169
rect 31113 9129 31125 9163
rect 31159 9160 31171 9163
rect 31202 9160 31208 9172
rect 31159 9132 31208 9160
rect 31159 9129 31171 9132
rect 31113 9123 31171 9129
rect 31202 9120 31208 9132
rect 31260 9120 31266 9172
rect 33870 9160 33876 9172
rect 31312 9132 33876 9160
rect 26988 9064 27384 9092
rect 27356 9024 27384 9064
rect 27816 9064 27936 9092
rect 27816 9024 27844 9064
rect 29546 9052 29552 9104
rect 29604 9052 29610 9104
rect 29638 9052 29644 9104
rect 29696 9052 29702 9104
rect 29564 9024 29592 9052
rect 27356 8996 27844 9024
rect 28966 8996 29592 9024
rect 27065 8959 27123 8965
rect 27065 8956 27077 8959
rect 26804 8928 27077 8956
rect 26697 8919 26755 8925
rect 27065 8925 27077 8928
rect 27111 8925 27123 8959
rect 27065 8919 27123 8925
rect 26528 8888 26556 8916
rect 25792 8860 26556 8888
rect 26620 8888 26648 8919
rect 27356 8900 27384 8996
rect 28445 8959 28503 8965
rect 28445 8925 28457 8959
rect 28491 8956 28503 8959
rect 28537 8959 28595 8965
rect 28537 8956 28549 8959
rect 28491 8928 28549 8956
rect 28491 8925 28503 8928
rect 28445 8919 28503 8925
rect 28537 8925 28549 8928
rect 28583 8925 28595 8959
rect 28537 8919 28595 8925
rect 28721 8959 28779 8965
rect 28721 8925 28733 8959
rect 28767 8956 28779 8959
rect 28966 8956 28994 8996
rect 28767 8928 28994 8956
rect 29181 8959 29239 8965
rect 28767 8925 28779 8928
rect 28721 8919 28779 8925
rect 29181 8925 29193 8959
rect 29227 8956 29239 8959
rect 29549 8959 29607 8965
rect 29549 8956 29561 8959
rect 29227 8928 29561 8956
rect 29227 8925 29239 8928
rect 29181 8919 29239 8925
rect 29549 8925 29561 8928
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 26620 8860 27292 8888
rect 27264 8832 27292 8860
rect 27338 8848 27344 8900
rect 27396 8848 27402 8900
rect 27522 8848 27528 8900
rect 27580 8897 27586 8900
rect 27580 8891 27615 8897
rect 27603 8888 27615 8891
rect 28814 8891 28872 8897
rect 28814 8888 28826 8891
rect 27603 8860 28826 8888
rect 27603 8857 27615 8860
rect 27580 8851 27615 8857
rect 28814 8857 28826 8860
rect 28860 8857 28872 8891
rect 28814 8851 28872 8857
rect 27580 8848 27586 8851
rect 28902 8848 28908 8900
rect 28960 8848 28966 8900
rect 29043 8891 29101 8897
rect 29043 8857 29055 8891
rect 29089 8888 29101 8891
rect 29270 8888 29276 8900
rect 29089 8860 29276 8888
rect 29089 8857 29101 8860
rect 29043 8851 29101 8857
rect 29270 8848 29276 8860
rect 29328 8888 29334 8900
rect 29748 8888 29776 9120
rect 29822 8984 29828 9036
rect 29880 9024 29886 9036
rect 31312 9033 31340 9132
rect 33870 9120 33876 9132
rect 33928 9120 33934 9172
rect 33965 9163 34023 9169
rect 33965 9129 33977 9163
rect 34011 9160 34023 9163
rect 34790 9160 34796 9172
rect 34011 9132 34796 9160
rect 34011 9129 34023 9132
rect 33965 9123 34023 9129
rect 34790 9120 34796 9132
rect 34848 9120 34854 9172
rect 33413 9095 33471 9101
rect 33413 9061 33425 9095
rect 33459 9092 33471 9095
rect 33502 9092 33508 9104
rect 33459 9064 33508 9092
rect 33459 9061 33471 9064
rect 33413 9055 33471 9061
rect 33502 9052 33508 9064
rect 33560 9052 33566 9104
rect 33888 9092 33916 9120
rect 34606 9092 34612 9104
rect 33888 9064 34612 9092
rect 34606 9052 34612 9064
rect 34664 9052 34670 9104
rect 30101 9027 30159 9033
rect 30101 9024 30113 9027
rect 29880 8996 30113 9024
rect 29880 8984 29886 8996
rect 30101 8993 30113 8996
rect 30147 8993 30159 9027
rect 30101 8987 30159 8993
rect 31297 9027 31355 9033
rect 31297 8993 31309 9027
rect 31343 8993 31355 9027
rect 31297 8987 31355 8993
rect 31573 9027 31631 9033
rect 31573 8993 31585 9027
rect 31619 9024 31631 9027
rect 32214 9024 32220 9036
rect 31619 8996 32220 9024
rect 31619 8993 31631 8996
rect 31573 8987 31631 8993
rect 32214 8984 32220 8996
rect 32272 8984 32278 9036
rect 33318 8984 33324 9036
rect 33376 8984 33382 9036
rect 30650 8916 30656 8968
rect 30708 8956 30714 8968
rect 30837 8959 30895 8965
rect 30837 8956 30849 8959
rect 30708 8928 30849 8956
rect 30708 8916 30714 8928
rect 30837 8925 30849 8928
rect 30883 8925 30895 8959
rect 30837 8919 30895 8925
rect 31205 8959 31263 8965
rect 31205 8925 31217 8959
rect 31251 8925 31263 8959
rect 33336 8956 33364 8984
rect 33597 8959 33655 8965
rect 33597 8956 33609 8959
rect 33336 8928 33609 8956
rect 31205 8919 31263 8925
rect 33597 8925 33609 8928
rect 33643 8925 33655 8959
rect 33597 8919 33655 8925
rect 29328 8860 29776 8888
rect 29328 8848 29334 8860
rect 31220 8832 31248 8919
rect 33686 8916 33692 8968
rect 33744 8916 33750 8968
rect 32030 8848 32036 8900
rect 32088 8848 32094 8900
rect 33226 8848 33232 8900
rect 33284 8888 33290 8900
rect 33781 8891 33839 8897
rect 33781 8888 33793 8891
rect 33284 8860 33793 8888
rect 33284 8848 33290 8860
rect 33781 8857 33793 8860
rect 33827 8857 33839 8891
rect 33781 8851 33839 8857
rect 21542 8820 21548 8832
rect 20119 8792 21548 8820
rect 20119 8789 20131 8792
rect 20073 8783 20131 8789
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 27246 8780 27252 8832
rect 27304 8780 27310 8832
rect 27709 8823 27767 8829
rect 27709 8789 27721 8823
rect 27755 8820 27767 8823
rect 28258 8820 28264 8832
rect 27755 8792 28264 8820
rect 27755 8789 27767 8792
rect 27709 8783 27767 8789
rect 28258 8780 28264 8792
rect 28316 8780 28322 8832
rect 28534 8780 28540 8832
rect 28592 8820 28598 8832
rect 30285 8823 30343 8829
rect 30285 8820 30297 8823
rect 28592 8792 30297 8820
rect 28592 8780 28598 8792
rect 30285 8789 30297 8792
rect 30331 8789 30343 8823
rect 30285 8783 30343 8789
rect 31202 8780 31208 8832
rect 31260 8780 31266 8832
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 18690 8616 18696 8628
rect 17092 8588 18696 8616
rect 17092 8576 17098 8588
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 19058 8576 19064 8628
rect 19116 8616 19122 8628
rect 19321 8619 19379 8625
rect 19321 8616 19333 8619
rect 19116 8588 19333 8616
rect 19116 8576 19122 8588
rect 19321 8585 19333 8588
rect 19367 8616 19379 8619
rect 19705 8619 19763 8625
rect 19705 8616 19717 8619
rect 19367 8588 19717 8616
rect 19367 8585 19379 8588
rect 19321 8579 19379 8585
rect 19705 8585 19717 8588
rect 19751 8585 19763 8619
rect 19705 8579 19763 8585
rect 19978 8576 19984 8628
rect 20036 8576 20042 8628
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20128 8588 20576 8616
rect 20128 8576 20134 8588
rect 17126 8508 17132 8560
rect 17184 8508 17190 8560
rect 18524 8520 18644 8548
rect 18322 8440 18328 8492
rect 18380 8440 18386 8492
rect 18524 8489 18552 8520
rect 18485 8483 18552 8489
rect 18485 8449 18497 8483
rect 18531 8452 18552 8483
rect 18616 8479 18644 8520
rect 19150 8508 19156 8560
rect 19208 8508 19214 8560
rect 19521 8551 19579 8557
rect 19521 8548 19533 8551
rect 19306 8520 19533 8548
rect 18616 8473 18675 8479
rect 18531 8449 18543 8452
rect 18485 8443 18543 8449
rect 18616 8442 18629 8473
rect 18617 8439 18629 8442
rect 18663 8470 18675 8473
rect 18663 8442 18736 8470
rect 18663 8439 18675 8442
rect 18617 8433 18675 8439
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8412 17371 8415
rect 17586 8412 17592 8424
rect 17359 8384 17592 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 18506 8304 18512 8356
rect 18564 8304 18570 8356
rect 18708 8344 18736 8442
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 19058 8440 19064 8492
rect 19116 8440 19122 8492
rect 19168 8480 19196 8508
rect 19306 8480 19334 8520
rect 19521 8517 19533 8520
rect 19567 8517 19579 8551
rect 19521 8511 19579 8517
rect 19996 8548 20024 8576
rect 20548 8557 20576 8588
rect 20806 8576 20812 8628
rect 20864 8576 20870 8628
rect 20993 8619 21051 8625
rect 20993 8585 21005 8619
rect 21039 8616 21051 8619
rect 21082 8616 21088 8628
rect 21039 8588 21088 8616
rect 21039 8585 21051 8588
rect 20993 8579 21051 8585
rect 21082 8576 21088 8588
rect 21140 8576 21146 8628
rect 21266 8576 21272 8628
rect 21324 8576 21330 8628
rect 22646 8576 22652 8628
rect 22704 8576 22710 8628
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23658 8616 23664 8628
rect 23523 8588 23664 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 23842 8576 23848 8628
rect 23900 8576 23906 8628
rect 25038 8576 25044 8628
rect 25096 8616 25102 8628
rect 27065 8619 27123 8625
rect 27065 8616 27077 8619
rect 25096 8588 27077 8616
rect 25096 8576 25102 8588
rect 27065 8585 27077 8588
rect 27111 8585 27123 8619
rect 30650 8616 30656 8628
rect 27065 8579 27123 8585
rect 28000 8588 30656 8616
rect 20714 8557 20720 8560
rect 20441 8551 20499 8557
rect 20441 8548 20453 8551
rect 19996 8520 20453 8548
rect 19168 8452 19334 8480
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8480 19855 8483
rect 19996 8480 20024 8520
rect 20441 8517 20453 8520
rect 20487 8517 20499 8551
rect 20441 8511 20499 8517
rect 20533 8551 20591 8557
rect 20533 8517 20545 8551
rect 20579 8517 20591 8551
rect 20533 8511 20591 8517
rect 20671 8551 20720 8557
rect 20671 8517 20683 8551
rect 20717 8517 20720 8551
rect 20671 8511 20720 8517
rect 20714 8508 20720 8511
rect 20772 8508 20778 8560
rect 19843 8452 20024 8480
rect 20349 8483 20407 8489
rect 19843 8449 19855 8452
rect 19797 8443 19855 8449
rect 20349 8449 20361 8483
rect 20395 8449 20407 8483
rect 20824 8480 20852 8576
rect 20901 8483 20959 8489
rect 20901 8480 20913 8483
rect 20824 8452 20913 8480
rect 20349 8443 20407 8449
rect 20901 8449 20913 8452
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8480 21143 8483
rect 21284 8480 21312 8576
rect 21131 8452 21312 8480
rect 21131 8449 21143 8452
rect 21085 8443 21143 8449
rect 19076 8412 19104 8440
rect 18892 8384 19104 8412
rect 20364 8412 20392 8443
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22373 8483 22431 8489
rect 22373 8480 22385 8483
rect 21968 8452 22385 8480
rect 21968 8440 21974 8452
rect 22373 8449 22385 8452
rect 22419 8449 22431 8483
rect 22373 8443 22431 8449
rect 22738 8440 22744 8492
rect 22796 8480 22802 8492
rect 23385 8483 23443 8489
rect 23385 8480 23397 8483
rect 22796 8452 23397 8480
rect 22796 8440 22802 8452
rect 23385 8449 23397 8452
rect 23431 8480 23443 8483
rect 23860 8480 23888 8576
rect 24946 8508 24952 8560
rect 25004 8548 25010 8560
rect 25004 8520 26188 8548
rect 25004 8508 25010 8520
rect 23431 8452 23888 8480
rect 24857 8483 24915 8489
rect 23431 8449 23443 8452
rect 23385 8443 23443 8449
rect 24857 8449 24869 8483
rect 24903 8480 24915 8483
rect 25314 8480 25320 8492
rect 24903 8452 25320 8480
rect 24903 8449 24915 8452
rect 24857 8443 24915 8449
rect 25314 8440 25320 8452
rect 25372 8480 25378 8492
rect 26160 8489 26188 8520
rect 27246 8508 27252 8560
rect 27304 8548 27310 8560
rect 28000 8548 28028 8588
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 30742 8576 30748 8628
rect 30800 8576 30806 8628
rect 30926 8576 30932 8628
rect 30984 8576 30990 8628
rect 31573 8619 31631 8625
rect 31573 8585 31585 8619
rect 31619 8616 31631 8619
rect 32030 8616 32036 8628
rect 31619 8588 32036 8616
rect 31619 8585 31631 8588
rect 31573 8579 31631 8585
rect 32030 8576 32036 8588
rect 32088 8576 32094 8628
rect 27304 8520 28028 8548
rect 27304 8508 27310 8520
rect 27356 8489 27384 8520
rect 28000 8489 28028 8520
rect 28077 8551 28135 8557
rect 28077 8517 28089 8551
rect 28123 8548 28135 8551
rect 29270 8548 29276 8560
rect 28123 8520 28396 8548
rect 28123 8517 28135 8520
rect 28077 8511 28135 8517
rect 26145 8483 26203 8489
rect 25372 8452 25912 8480
rect 25372 8440 25378 8452
rect 20809 8415 20867 8421
rect 20364 8384 20576 8412
rect 18892 8344 18920 8384
rect 20548 8356 20576 8384
rect 20809 8381 20821 8415
rect 20855 8412 20867 8415
rect 21821 8415 21879 8421
rect 21821 8412 21833 8415
rect 20855 8384 21833 8412
rect 20855 8381 20867 8384
rect 20809 8375 20867 8381
rect 21821 8381 21833 8384
rect 21867 8381 21879 8415
rect 21821 8375 21879 8381
rect 24118 8372 24124 8424
rect 24176 8412 24182 8424
rect 24670 8412 24676 8424
rect 24176 8384 24676 8412
rect 24176 8372 24182 8384
rect 24670 8372 24676 8384
rect 24728 8372 24734 8424
rect 24765 8415 24823 8421
rect 24765 8381 24777 8415
rect 24811 8381 24823 8415
rect 24765 8375 24823 8381
rect 18708 8316 18920 8344
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 19610 8344 19616 8356
rect 19300 8316 19616 8344
rect 19300 8304 19306 8316
rect 19610 8304 19616 8316
rect 19668 8304 19674 8356
rect 20530 8304 20536 8356
rect 20588 8304 20594 8356
rect 24780 8344 24808 8375
rect 24946 8372 24952 8424
rect 25004 8372 25010 8424
rect 25777 8415 25835 8421
rect 25777 8381 25789 8415
rect 25823 8381 25835 8415
rect 25884 8412 25912 8452
rect 26145 8449 26157 8483
rect 26191 8449 26203 8483
rect 26145 8443 26203 8449
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8449 27491 8483
rect 27433 8443 27491 8449
rect 27985 8483 28043 8489
rect 27985 8449 27997 8483
rect 28031 8449 28043 8483
rect 27985 8443 28043 8449
rect 26329 8415 26387 8421
rect 26329 8412 26341 8415
rect 25884 8384 26341 8412
rect 25777 8375 25835 8381
rect 26329 8381 26341 8384
rect 26375 8381 26387 8415
rect 26329 8375 26387 8381
rect 25792 8344 25820 8375
rect 27154 8372 27160 8424
rect 27212 8412 27218 8424
rect 27448 8412 27476 8443
rect 28166 8440 28172 8492
rect 28224 8440 28230 8492
rect 28258 8440 28264 8492
rect 28316 8440 28322 8492
rect 28368 8480 28396 8520
rect 28644 8520 29276 8548
rect 28445 8483 28503 8489
rect 28445 8480 28457 8483
rect 28368 8452 28457 8480
rect 28445 8449 28457 8452
rect 28491 8449 28503 8483
rect 28445 8443 28503 8449
rect 28534 8440 28540 8492
rect 28592 8440 28598 8492
rect 28644 8489 28672 8520
rect 29270 8508 29276 8520
rect 29328 8508 29334 8560
rect 30190 8508 30196 8560
rect 30248 8508 30254 8560
rect 28629 8483 28687 8489
rect 28629 8449 28641 8483
rect 28675 8449 28687 8483
rect 28810 8480 28816 8492
rect 28629 8443 28687 8449
rect 28736 8452 28816 8480
rect 28736 8412 28764 8452
rect 28810 8440 28816 8452
rect 28868 8440 28874 8492
rect 28902 8440 28908 8492
rect 28960 8440 28966 8492
rect 30944 8489 30972 8576
rect 30929 8483 30987 8489
rect 30929 8449 30941 8483
rect 30975 8449 30987 8483
rect 30929 8443 30987 8449
rect 31481 8483 31539 8489
rect 31481 8449 31493 8483
rect 31527 8449 31539 8483
rect 31481 8443 31539 8449
rect 29181 8415 29239 8421
rect 29181 8412 29193 8415
rect 27212 8384 28764 8412
rect 28828 8384 29193 8412
rect 27212 8372 27218 8384
rect 25866 8344 25872 8356
rect 24780 8316 25872 8344
rect 25866 8304 25872 8316
rect 25924 8304 25930 8356
rect 28258 8304 28264 8356
rect 28316 8344 28322 8356
rect 28828 8353 28856 8384
rect 29181 8381 29193 8384
rect 29227 8381 29239 8415
rect 31202 8412 31208 8424
rect 29181 8375 29239 8381
rect 30300 8384 31208 8412
rect 28813 8347 28871 8353
rect 28316 8316 28764 8344
rect 28316 8304 28322 8316
rect 16666 8236 16672 8288
rect 16724 8236 16730 8288
rect 19058 8236 19064 8288
rect 19116 8236 19122 8288
rect 19150 8236 19156 8288
rect 19208 8236 19214 8288
rect 19334 8236 19340 8288
rect 19392 8236 19398 8288
rect 20162 8236 20168 8288
rect 20220 8236 20226 8288
rect 25130 8236 25136 8288
rect 25188 8236 25194 8288
rect 25222 8236 25228 8288
rect 25280 8236 25286 8288
rect 25958 8236 25964 8288
rect 26016 8236 26022 8288
rect 27338 8236 27344 8288
rect 27396 8236 27402 8288
rect 28736 8276 28764 8316
rect 28813 8313 28825 8347
rect 28859 8313 28871 8347
rect 28813 8307 28871 8313
rect 30300 8288 30328 8384
rect 31202 8372 31208 8384
rect 31260 8412 31266 8424
rect 31496 8412 31524 8443
rect 31260 8384 31524 8412
rect 31260 8372 31266 8384
rect 29178 8276 29184 8288
rect 28736 8248 29184 8276
rect 29178 8236 29184 8248
rect 29236 8236 29242 8288
rect 30282 8236 30288 8288
rect 30340 8236 30346 8288
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 17313 8075 17371 8081
rect 17313 8041 17325 8075
rect 17359 8072 17371 8075
rect 17586 8072 17592 8084
rect 17359 8044 17592 8072
rect 17359 8041 17371 8044
rect 17313 8035 17371 8041
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 19242 8072 19248 8084
rect 18564 8044 19248 8072
rect 18564 8032 18570 8044
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 28166 8032 28172 8084
rect 28224 8032 28230 8084
rect 29181 8075 29239 8081
rect 29181 8041 29193 8075
rect 29227 8072 29239 8075
rect 29546 8072 29552 8084
rect 29227 8044 29552 8072
rect 29227 8041 29239 8044
rect 29181 8035 29239 8041
rect 29546 8032 29552 8044
rect 29604 8032 29610 8084
rect 30190 8032 30196 8084
rect 30248 8032 30254 8084
rect 24762 7964 24768 8016
rect 24820 8004 24826 8016
rect 24820 7976 25912 8004
rect 24820 7964 24826 7976
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 15838 7936 15844 7948
rect 15620 7908 15844 7936
rect 15620 7896 15626 7908
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 19058 7936 19064 7948
rect 18340 7908 19064 7936
rect 18340 7877 18368 7908
rect 19058 7896 19064 7908
rect 19116 7936 19122 7948
rect 19705 7939 19763 7945
rect 19705 7936 19717 7939
rect 19116 7908 19717 7936
rect 19116 7896 19122 7908
rect 19705 7905 19717 7908
rect 19751 7905 19763 7939
rect 19705 7899 19763 7905
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 20070 7936 20076 7948
rect 19935 7908 20076 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 25041 7939 25099 7945
rect 25041 7905 25053 7939
rect 25087 7936 25099 7939
rect 25777 7939 25835 7945
rect 25777 7936 25789 7939
rect 25087 7908 25789 7936
rect 25087 7905 25099 7908
rect 25041 7899 25099 7905
rect 25777 7905 25789 7908
rect 25823 7905 25835 7939
rect 25777 7899 25835 7905
rect 25884 7936 25912 7976
rect 28184 7936 28212 8032
rect 25884 7908 26188 7936
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 15841 7803 15899 7809
rect 15841 7769 15853 7803
rect 15887 7800 15899 7803
rect 15930 7800 15936 7812
rect 15887 7772 15936 7800
rect 15887 7769 15899 7772
rect 15841 7763 15899 7769
rect 15930 7760 15936 7772
rect 15988 7760 15994 7812
rect 16850 7760 16856 7812
rect 16908 7760 16914 7812
rect 18064 7800 18092 7831
rect 18966 7828 18972 7880
rect 19024 7828 19030 7880
rect 19150 7828 19156 7880
rect 19208 7828 19214 7880
rect 19610 7828 19616 7880
rect 19668 7828 19674 7880
rect 21269 7871 21327 7877
rect 21269 7837 21281 7871
rect 21315 7868 21327 7871
rect 21818 7868 21824 7880
rect 21315 7840 21824 7868
rect 21315 7837 21327 7840
rect 21269 7831 21327 7837
rect 21818 7828 21824 7840
rect 21876 7868 21882 7880
rect 22738 7868 22744 7880
rect 21876 7840 22744 7868
rect 21876 7828 21882 7840
rect 22738 7828 22744 7840
rect 22796 7828 22802 7880
rect 24118 7828 24124 7880
rect 24176 7868 24182 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 24176 7840 24409 7868
rect 24176 7828 24182 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 25130 7828 25136 7880
rect 25188 7868 25194 7880
rect 25317 7871 25375 7877
rect 25317 7868 25329 7871
rect 25188 7840 25329 7868
rect 25188 7828 25194 7840
rect 25317 7837 25329 7840
rect 25363 7837 25375 7871
rect 25317 7831 25375 7837
rect 25501 7871 25559 7877
rect 25501 7837 25513 7871
rect 25547 7868 25559 7871
rect 25884 7868 25912 7908
rect 26160 7880 26188 7908
rect 27080 7908 28212 7936
rect 25547 7840 25912 7868
rect 25547 7837 25559 7840
rect 25501 7831 25559 7837
rect 26050 7828 26056 7880
rect 26108 7828 26114 7880
rect 26142 7828 26148 7880
rect 26200 7868 26206 7880
rect 26602 7868 26608 7880
rect 26200 7840 26608 7868
rect 26200 7828 26206 7840
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 27080 7877 27108 7908
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7868 27307 7871
rect 27522 7868 27528 7880
rect 27295 7840 27528 7868
rect 27295 7837 27307 7840
rect 27249 7831 27307 7837
rect 27522 7828 27528 7840
rect 27580 7828 27586 7880
rect 27890 7828 27896 7880
rect 27948 7828 27954 7880
rect 28184 7868 28212 7908
rect 28997 7871 29055 7877
rect 28997 7868 29009 7871
rect 28184 7840 29009 7868
rect 28997 7837 29009 7840
rect 29043 7837 29055 7871
rect 28997 7831 29055 7837
rect 29178 7828 29184 7880
rect 29236 7828 29242 7880
rect 30282 7828 30288 7880
rect 30340 7828 30346 7880
rect 19168 7800 19196 7828
rect 18064 7772 19196 7800
rect 25409 7803 25467 7809
rect 25409 7769 25421 7803
rect 25455 7769 25467 7803
rect 25409 7763 25467 7769
rect 17862 7692 17868 7744
rect 17920 7692 17926 7744
rect 18233 7735 18291 7741
rect 18233 7701 18245 7735
rect 18279 7732 18291 7735
rect 18417 7735 18475 7741
rect 18417 7732 18429 7735
rect 18279 7704 18429 7732
rect 18279 7701 18291 7704
rect 18233 7695 18291 7701
rect 18417 7701 18429 7704
rect 18463 7701 18475 7735
rect 18417 7695 18475 7701
rect 19242 7692 19248 7744
rect 19300 7692 19306 7744
rect 21174 7692 21180 7744
rect 21232 7692 21238 7744
rect 22830 7692 22836 7744
rect 22888 7692 22894 7744
rect 23658 7692 23664 7744
rect 23716 7732 23722 7744
rect 25133 7735 25191 7741
rect 25133 7732 25145 7735
rect 23716 7704 25145 7732
rect 23716 7692 23722 7704
rect 25133 7701 25145 7704
rect 25179 7701 25191 7735
rect 25424 7732 25452 7763
rect 25590 7760 25596 7812
rect 25648 7809 25654 7812
rect 25648 7803 25697 7809
rect 25648 7769 25651 7803
rect 25685 7800 25697 7803
rect 27908 7800 27936 7828
rect 25685 7772 27936 7800
rect 25685 7769 25697 7772
rect 25648 7763 25697 7769
rect 25648 7760 25654 7763
rect 29730 7760 29736 7812
rect 29788 7800 29794 7812
rect 30300 7800 30328 7828
rect 29788 7772 30328 7800
rect 29788 7760 29794 7772
rect 25961 7735 26019 7741
rect 25961 7732 25973 7735
rect 25424 7704 25973 7732
rect 25133 7695 25191 7701
rect 25961 7701 25973 7704
rect 26007 7701 26019 7735
rect 25961 7695 26019 7701
rect 27157 7735 27215 7741
rect 27157 7701 27169 7735
rect 27203 7732 27215 7735
rect 27798 7732 27804 7744
rect 27203 7704 27804 7732
rect 27203 7701 27215 7704
rect 27157 7695 27215 7701
rect 27798 7692 27804 7704
rect 27856 7692 27862 7744
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15988 7500 16037 7528
rect 15988 7488 15994 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16025 7491 16083 7497
rect 16666 7488 16672 7540
rect 16724 7488 16730 7540
rect 16761 7531 16819 7537
rect 16761 7497 16773 7531
rect 16807 7528 16819 7531
rect 16850 7528 16856 7540
rect 16807 7500 16856 7528
rect 16807 7497 16819 7500
rect 16761 7491 16819 7497
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 17862 7528 17868 7540
rect 17604 7500 17868 7528
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 16684 7392 16712 7488
rect 17604 7469 17632 7500
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18966 7488 18972 7540
rect 19024 7528 19030 7540
rect 19061 7531 19119 7537
rect 19061 7528 19073 7531
rect 19024 7500 19073 7528
rect 19024 7488 19030 7500
rect 19061 7497 19073 7500
rect 19107 7497 19119 7531
rect 19061 7491 19119 7497
rect 19242 7488 19248 7540
rect 19300 7488 19306 7540
rect 22002 7528 22008 7540
rect 19904 7500 22008 7528
rect 17589 7463 17647 7469
rect 17589 7429 17601 7463
rect 17635 7429 17647 7463
rect 17589 7423 17647 7429
rect 18322 7420 18328 7472
rect 18380 7420 18386 7472
rect 16255 7364 16712 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16816 7364 16865 7392
rect 16816 7352 16822 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 19260 7392 19288 7488
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 19260 7364 19349 7392
rect 16853 7355 16911 7361
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 19904 7401 19932 7500
rect 22002 7488 22008 7500
rect 22060 7528 22066 7540
rect 22060 7500 22140 7528
rect 22060 7488 22066 7500
rect 20162 7420 20168 7472
rect 20220 7420 20226 7472
rect 21174 7420 21180 7472
rect 21232 7420 21238 7472
rect 22112 7460 22140 7500
rect 23658 7488 23664 7540
rect 23716 7488 23722 7540
rect 24118 7488 24124 7540
rect 24176 7528 24182 7540
rect 25501 7531 25559 7537
rect 24176 7500 25176 7528
rect 24176 7488 24182 7500
rect 22186 7460 22192 7472
rect 21928 7432 22192 7460
rect 21928 7401 21956 7432
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 22830 7420 22836 7472
rect 22888 7420 22894 7472
rect 19889 7395 19947 7401
rect 19889 7392 19901 7395
rect 19852 7364 19901 7392
rect 19852 7352 19858 7364
rect 19889 7361 19901 7364
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 21913 7395 21971 7401
rect 21913 7361 21925 7395
rect 21959 7361 21971 7395
rect 21913 7355 21971 7361
rect 15838 7284 15844 7336
rect 15896 7324 15902 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 15896 7296 17325 7324
rect 15896 7284 15902 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 22189 7327 22247 7333
rect 22189 7293 22201 7327
rect 22235 7324 22247 7327
rect 23676 7324 23704 7488
rect 24213 7463 24271 7469
rect 24213 7429 24225 7463
rect 24259 7460 24271 7463
rect 24673 7463 24731 7469
rect 24673 7460 24685 7463
rect 24259 7432 24685 7460
rect 24259 7429 24271 7432
rect 24213 7423 24271 7429
rect 24673 7429 24685 7432
rect 24719 7429 24731 7463
rect 24673 7423 24731 7429
rect 24762 7420 24768 7472
rect 24820 7420 24826 7472
rect 25148 7469 25176 7500
rect 25501 7497 25513 7531
rect 25547 7528 25559 7531
rect 26050 7528 26056 7540
rect 25547 7500 26056 7528
rect 25547 7497 25559 7500
rect 25501 7491 25559 7497
rect 26050 7488 26056 7500
rect 26108 7528 26114 7540
rect 26789 7531 26847 7537
rect 26108 7500 26648 7528
rect 26108 7488 26114 7500
rect 25133 7463 25191 7469
rect 25133 7429 25145 7463
rect 25179 7429 25191 7463
rect 25133 7423 25191 7429
rect 25349 7463 25407 7469
rect 25349 7429 25361 7463
rect 25395 7460 25407 7463
rect 25958 7460 25964 7472
rect 25395 7432 25964 7460
rect 25395 7429 25407 7432
rect 25349 7423 25407 7429
rect 24946 7401 24952 7404
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7392 24179 7395
rect 24305 7395 24363 7401
rect 24167 7364 24256 7392
rect 24167 7361 24179 7364
rect 24121 7355 24179 7361
rect 22235 7296 23704 7324
rect 22235 7293 22247 7296
rect 22189 7287 22247 7293
rect 24228 7268 24256 7364
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 24581 7395 24639 7401
rect 24581 7361 24593 7395
rect 24627 7392 24639 7395
rect 24903 7395 24952 7401
rect 24627 7364 24808 7392
rect 24627 7361 24639 7364
rect 24581 7355 24639 7361
rect 24320 7324 24348 7355
rect 24780 7324 24808 7364
rect 24903 7361 24915 7395
rect 24949 7361 24952 7395
rect 24903 7355 24952 7361
rect 24946 7352 24952 7355
rect 25004 7352 25010 7404
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7392 25099 7395
rect 25222 7392 25228 7404
rect 25087 7364 25228 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 25593 7327 25651 7333
rect 25593 7324 25605 7327
rect 24320 7296 24624 7324
rect 24780 7296 25605 7324
rect 21637 7259 21695 7265
rect 21637 7225 21649 7259
rect 21683 7256 21695 7259
rect 21910 7256 21916 7268
rect 21683 7228 21916 7256
rect 21683 7225 21695 7228
rect 21637 7219 21695 7225
rect 21910 7216 21916 7228
rect 21968 7216 21974 7268
rect 23661 7259 23719 7265
rect 23661 7225 23673 7259
rect 23707 7256 23719 7259
rect 24118 7256 24124 7268
rect 23707 7228 24124 7256
rect 23707 7225 23719 7228
rect 23661 7219 23719 7225
rect 24118 7216 24124 7228
rect 24176 7216 24182 7268
rect 24210 7216 24216 7268
rect 24268 7256 24274 7268
rect 24596 7256 24624 7296
rect 25593 7293 25605 7296
rect 25639 7293 25651 7327
rect 25593 7287 25651 7293
rect 25700 7256 25728 7432
rect 25958 7420 25964 7432
rect 26016 7420 26022 7472
rect 25777 7395 25835 7401
rect 25777 7361 25789 7395
rect 25823 7392 25835 7395
rect 25866 7392 25872 7404
rect 25823 7364 25872 7392
rect 25823 7361 25835 7364
rect 25777 7355 25835 7361
rect 24268 7228 24532 7256
rect 24596 7228 25728 7256
rect 24268 7216 24274 7228
rect 19518 7148 19524 7200
rect 19576 7148 19582 7200
rect 24394 7148 24400 7200
rect 24452 7148 24458 7200
rect 24504 7188 24532 7228
rect 25317 7191 25375 7197
rect 25317 7188 25329 7191
rect 24504 7160 25329 7188
rect 25317 7157 25329 7160
rect 25363 7188 25375 7191
rect 25792 7188 25820 7355
rect 25866 7352 25872 7364
rect 25924 7352 25930 7404
rect 26620 7401 26648 7500
rect 26789 7497 26801 7531
rect 26835 7528 26847 7531
rect 27154 7528 27160 7540
rect 26835 7500 27160 7528
rect 26835 7497 26847 7500
rect 26789 7491 26847 7497
rect 27154 7488 27160 7500
rect 27212 7528 27218 7540
rect 27522 7528 27528 7540
rect 27212 7500 27528 7528
rect 27212 7488 27218 7500
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 27798 7420 27804 7472
rect 27856 7460 27862 7472
rect 28074 7460 28080 7472
rect 27856 7432 28080 7460
rect 27856 7420 27862 7432
rect 28074 7420 28080 7432
rect 28132 7460 28138 7472
rect 28169 7463 28227 7469
rect 28169 7460 28181 7463
rect 28132 7432 28181 7460
rect 28132 7420 28138 7432
rect 28169 7429 28181 7432
rect 28215 7429 28227 7463
rect 28169 7423 28227 7429
rect 26605 7395 26663 7401
rect 26605 7361 26617 7395
rect 26651 7361 26663 7395
rect 26605 7355 26663 7361
rect 26421 7327 26479 7333
rect 26421 7293 26433 7327
rect 26467 7324 26479 7327
rect 26510 7324 26516 7336
rect 26467 7296 26516 7324
rect 26467 7293 26479 7296
rect 26421 7287 26479 7293
rect 26510 7284 26516 7296
rect 26568 7284 26574 7336
rect 26620 7256 26648 7355
rect 27338 7352 27344 7404
rect 27396 7352 27402 7404
rect 27890 7352 27896 7404
rect 27948 7392 27954 7404
rect 27985 7395 28043 7401
rect 27985 7392 27997 7395
rect 27948 7364 27997 7392
rect 27948 7352 27954 7364
rect 27985 7361 27997 7364
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 27062 7284 27068 7336
rect 27120 7284 27126 7336
rect 27249 7327 27307 7333
rect 27249 7293 27261 7327
rect 27295 7324 27307 7327
rect 27798 7324 27804 7336
rect 27295 7296 27804 7324
rect 27295 7293 27307 7296
rect 27249 7287 27307 7293
rect 27798 7284 27804 7296
rect 27856 7284 27862 7336
rect 27982 7256 27988 7268
rect 26620 7228 27988 7256
rect 27982 7216 27988 7228
rect 28040 7216 28046 7268
rect 25363 7160 25820 7188
rect 27709 7191 27767 7197
rect 25363 7157 25375 7160
rect 25317 7151 25375 7157
rect 27709 7157 27721 7191
rect 27755 7188 27767 7191
rect 28166 7188 28172 7200
rect 27755 7160 28172 7188
rect 27755 7157 27767 7160
rect 27709 7151 27767 7157
rect 28166 7148 28172 7160
rect 28224 7148 28230 7200
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 16758 6944 16764 6996
rect 16816 6944 16822 6996
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 18417 6987 18475 6993
rect 18417 6984 18429 6987
rect 18380 6956 18429 6984
rect 18380 6944 18386 6956
rect 18417 6953 18429 6956
rect 18463 6953 18475 6987
rect 18417 6947 18475 6953
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 20054 6987 20112 6993
rect 20054 6984 20066 6987
rect 19576 6956 20066 6984
rect 19576 6944 19582 6956
rect 20054 6953 20066 6956
rect 20100 6953 20112 6987
rect 20054 6947 20112 6953
rect 22452 6987 22510 6993
rect 22452 6953 22464 6987
rect 22498 6984 22510 6987
rect 24394 6984 24400 6996
rect 22498 6956 24400 6984
rect 22498 6953 22510 6956
rect 22452 6947 22510 6953
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 27338 6944 27344 6996
rect 27396 6944 27402 6996
rect 16776 6916 16804 6944
rect 16776 6888 18368 6916
rect 18340 6789 18368 6888
rect 26712 6888 27568 6916
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 21545 6851 21603 6857
rect 21545 6848 21557 6851
rect 20128 6820 21557 6848
rect 20128 6808 20134 6820
rect 21545 6817 21557 6820
rect 21591 6817 21603 6851
rect 21545 6811 21603 6817
rect 22186 6808 22192 6860
rect 22244 6808 22250 6860
rect 24210 6808 24216 6860
rect 24268 6808 24274 6860
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 26712 6848 26740 6888
rect 26559 6820 26740 6848
rect 26789 6851 26847 6857
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 26789 6817 26801 6851
rect 26835 6848 26847 6851
rect 27430 6848 27436 6860
rect 26835 6820 27436 6848
rect 26835 6817 26847 6820
rect 26789 6811 26847 6817
rect 27430 6808 27436 6820
rect 27488 6808 27494 6860
rect 27540 6848 27568 6888
rect 28810 6876 28816 6928
rect 28868 6876 28874 6928
rect 28258 6848 28264 6860
rect 27540 6820 28264 6848
rect 28258 6808 28264 6820
rect 28316 6808 28322 6860
rect 28828 6848 28856 6876
rect 29181 6851 29239 6857
rect 29181 6848 29193 6851
rect 28828 6820 29193 6848
rect 29181 6817 29193 6820
rect 29227 6817 29239 6851
rect 29181 6811 29239 6817
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 19794 6740 19800 6792
rect 19852 6740 19858 6792
rect 21818 6740 21824 6792
rect 21876 6740 21882 6792
rect 23566 6740 23572 6792
rect 23624 6740 23630 6792
rect 26973 6783 27031 6789
rect 26973 6749 26985 6783
rect 27019 6749 27031 6783
rect 26973 6743 27031 6749
rect 21729 6715 21787 6721
rect 21729 6712 21741 6715
rect 21298 6684 21741 6712
rect 21729 6681 21741 6684
rect 21775 6681 21787 6715
rect 21729 6675 21787 6681
rect 26050 6672 26056 6724
rect 26108 6672 26114 6724
rect 26510 6672 26516 6724
rect 26568 6672 26574 6724
rect 26602 6672 26608 6724
rect 26660 6712 26666 6724
rect 26988 6712 27016 6743
rect 27154 6740 27160 6792
rect 27212 6740 27218 6792
rect 29730 6740 29736 6792
rect 29788 6740 29794 6792
rect 26660 6684 27016 6712
rect 26660 6672 26666 6684
rect 27706 6672 27712 6724
rect 27764 6672 27770 6724
rect 29641 6715 29699 6721
rect 29641 6712 29653 6715
rect 28934 6684 29653 6712
rect 29641 6681 29653 6684
rect 29687 6681 29699 6715
rect 29641 6675 29699 6681
rect 25041 6647 25099 6653
rect 25041 6613 25053 6647
rect 25087 6644 25099 6647
rect 26528 6644 26556 6672
rect 25087 6616 26556 6644
rect 25087 6613 25099 6616
rect 25041 6607 25099 6613
rect 29454 6604 29460 6656
rect 29512 6644 29518 6656
rect 29748 6644 29776 6740
rect 29512 6616 29776 6644
rect 29512 6604 29518 6616
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 23566 6400 23572 6452
rect 23624 6400 23630 6452
rect 23842 6400 23848 6452
rect 23900 6400 23906 6452
rect 26050 6400 26056 6452
rect 26108 6440 26114 6452
rect 26145 6443 26203 6449
rect 26145 6440 26157 6443
rect 26108 6412 26157 6440
rect 26108 6400 26114 6412
rect 26145 6409 26157 6412
rect 26191 6409 26203 6443
rect 26145 6403 26203 6409
rect 27706 6400 27712 6452
rect 27764 6440 27770 6452
rect 28353 6443 28411 6449
rect 28353 6440 28365 6443
rect 27764 6412 28365 6440
rect 27764 6400 27770 6412
rect 28353 6409 28365 6412
rect 28399 6409 28411 6443
rect 28353 6403 28411 6409
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6304 23719 6307
rect 23860 6304 23888 6400
rect 27798 6332 27804 6384
rect 27856 6372 27862 6384
rect 27893 6375 27951 6381
rect 27893 6372 27905 6375
rect 27856 6344 27905 6372
rect 27856 6332 27862 6344
rect 27893 6341 27905 6344
rect 27939 6341 27951 6375
rect 27893 6335 27951 6341
rect 27982 6332 27988 6384
rect 28040 6332 28046 6384
rect 28166 6332 28172 6384
rect 28224 6332 28230 6384
rect 23707 6276 23888 6304
rect 26053 6307 26111 6313
rect 23707 6273 23719 6276
rect 23661 6267 23719 6273
rect 26053 6273 26065 6307
rect 26099 6273 26111 6307
rect 26053 6267 26111 6273
rect 26068 6236 26096 6267
rect 26510 6264 26516 6316
rect 26568 6304 26574 6316
rect 26973 6307 27031 6313
rect 26973 6304 26985 6307
rect 26568 6276 26985 6304
rect 26568 6264 26574 6276
rect 26973 6273 26985 6276
rect 27019 6273 27031 6307
rect 26973 6267 27031 6273
rect 27617 6307 27675 6313
rect 27617 6273 27629 6307
rect 27663 6304 27675 6307
rect 27709 6307 27767 6313
rect 27709 6304 27721 6307
rect 27663 6276 27721 6304
rect 27663 6273 27675 6276
rect 27617 6267 27675 6273
rect 27709 6273 27721 6276
rect 27755 6273 27767 6307
rect 27709 6267 27767 6273
rect 28074 6264 28080 6316
rect 28132 6264 28138 6316
rect 28184 6304 28212 6332
rect 28537 6307 28595 6313
rect 28537 6304 28549 6307
rect 28184 6276 28549 6304
rect 28537 6273 28549 6276
rect 28583 6273 28595 6307
rect 28537 6267 28595 6273
rect 29454 6236 29460 6248
rect 26068 6208 29460 6236
rect 29454 6196 29460 6208
rect 29512 6196 29518 6248
rect 28258 6128 28264 6180
rect 28316 6128 28322 6180
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 13722 3516 13728 3528
rect 8444 3488 13728 3516
rect 8444 3476 8450 3488
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 20346 3000 20352 3052
rect 20404 3040 20410 3052
rect 43073 3043 43131 3049
rect 43073 3040 43085 3043
rect 20404 3012 43085 3040
rect 20404 3000 20410 3012
rect 43073 3009 43085 3012
rect 43119 3009 43131 3043
rect 43073 3003 43131 3009
rect 43254 2796 43260 2848
rect 43312 2796 43318 2848
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 26510 2388 26516 2440
rect 26568 2388 26574 2440
rect 43254 2388 43260 2440
rect 43312 2428 43318 2440
rect 43993 2431 44051 2437
rect 43993 2428 44005 2431
rect 43312 2400 44005 2428
rect 43312 2388 43318 2400
rect 43993 2397 44005 2400
rect 44039 2397 44051 2431
rect 43993 2391 44051 2397
rect 67634 2388 67640 2440
rect 67692 2388 67698 2440
rect 43806 2252 43812 2304
rect 43864 2292 43870 2304
rect 44269 2295 44327 2301
rect 44269 2292 44281 2295
rect 43864 2264 44281 2292
rect 43864 2252 43870 2264
rect 44269 2261 44281 2264
rect 44315 2261 44327 2295
rect 44269 2255 44327 2261
rect 67913 2295 67971 2301
rect 67913 2261 67925 2295
rect 67959 2292 67971 2295
rect 68002 2292 68008 2304
rect 67959 2264 68008 2292
rect 67959 2261 67971 2264
rect 67913 2255 67971 2261
rect 68002 2252 68008 2264
rect 68060 2252 68066 2304
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
<< via1 >>
rect 19574 67430 19626 67482
rect 19638 67430 19690 67482
rect 19702 67430 19754 67482
rect 19766 67430 19818 67482
rect 19830 67430 19882 67482
rect 50294 67430 50346 67482
rect 50358 67430 50410 67482
rect 50422 67430 50474 67482
rect 50486 67430 50538 67482
rect 50550 67430 50602 67482
rect 12992 67235 13044 67244
rect 12992 67201 13001 67235
rect 13001 67201 13035 67235
rect 13035 67201 13044 67235
rect 12992 67192 13044 67201
rect 30380 67235 30432 67244
rect 30380 67201 30389 67235
rect 30389 67201 30423 67235
rect 30423 67201 30432 67235
rect 30380 67192 30432 67201
rect 39396 67235 39448 67244
rect 39396 67201 39405 67235
rect 39405 67201 39439 67235
rect 39439 67201 39448 67235
rect 39396 67192 39448 67201
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 19574 66342 19626 66394
rect 19638 66342 19690 66394
rect 19702 66342 19754 66394
rect 19766 66342 19818 66394
rect 19830 66342 19882 66394
rect 50294 66342 50346 66394
rect 50358 66342 50410 66394
rect 50422 66342 50474 66394
rect 50486 66342 50538 66394
rect 50550 66342 50602 66394
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 19574 65254 19626 65306
rect 19638 65254 19690 65306
rect 19702 65254 19754 65306
rect 19766 65254 19818 65306
rect 19830 65254 19882 65306
rect 50294 65254 50346 65306
rect 50358 65254 50410 65306
rect 50422 65254 50474 65306
rect 50486 65254 50538 65306
rect 50550 65254 50602 65306
rect 1400 64991 1452 65000
rect 1400 64957 1409 64991
rect 1409 64957 1443 64991
rect 1443 64957 1452 64991
rect 1400 64948 1452 64957
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 34934 64710 34986 64762
rect 34998 64710 35050 64762
rect 35062 64710 35114 64762
rect 35126 64710 35178 64762
rect 35190 64710 35242 64762
rect 65654 64710 65706 64762
rect 65718 64710 65770 64762
rect 65782 64710 65834 64762
rect 65846 64710 65898 64762
rect 65910 64710 65962 64762
rect 19574 64166 19626 64218
rect 19638 64166 19690 64218
rect 19702 64166 19754 64218
rect 19766 64166 19818 64218
rect 19830 64166 19882 64218
rect 50294 64166 50346 64218
rect 50358 64166 50410 64218
rect 50422 64166 50474 64218
rect 50486 64166 50538 64218
rect 50550 64166 50602 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 34934 63622 34986 63674
rect 34998 63622 35050 63674
rect 35062 63622 35114 63674
rect 35126 63622 35178 63674
rect 35190 63622 35242 63674
rect 65654 63622 65706 63674
rect 65718 63622 65770 63674
rect 65782 63622 65834 63674
rect 65846 63622 65898 63674
rect 65910 63622 65962 63674
rect 19574 63078 19626 63130
rect 19638 63078 19690 63130
rect 19702 63078 19754 63130
rect 19766 63078 19818 63130
rect 19830 63078 19882 63130
rect 50294 63078 50346 63130
rect 50358 63078 50410 63130
rect 50422 63078 50474 63130
rect 50486 63078 50538 63130
rect 50550 63078 50602 63130
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 34934 62534 34986 62586
rect 34998 62534 35050 62586
rect 35062 62534 35114 62586
rect 35126 62534 35178 62586
rect 35190 62534 35242 62586
rect 65654 62534 65706 62586
rect 65718 62534 65770 62586
rect 65782 62534 65834 62586
rect 65846 62534 65898 62586
rect 65910 62534 65962 62586
rect 19574 61990 19626 62042
rect 19638 61990 19690 62042
rect 19702 61990 19754 62042
rect 19766 61990 19818 62042
rect 19830 61990 19882 62042
rect 50294 61990 50346 62042
rect 50358 61990 50410 62042
rect 50422 61990 50474 62042
rect 50486 61990 50538 62042
rect 50550 61990 50602 62042
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 65654 61446 65706 61498
rect 65718 61446 65770 61498
rect 65782 61446 65834 61498
rect 65846 61446 65898 61498
rect 65910 61446 65962 61498
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 65654 60358 65706 60410
rect 65718 60358 65770 60410
rect 65782 60358 65834 60410
rect 65846 60358 65898 60410
rect 65910 60358 65962 60410
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 65654 59270 65706 59322
rect 65718 59270 65770 59322
rect 65782 59270 65834 59322
rect 65846 59270 65898 59322
rect 65910 59270 65962 59322
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 65654 58182 65706 58234
rect 65718 58182 65770 58234
rect 65782 58182 65834 58234
rect 65846 58182 65898 58234
rect 65910 58182 65962 58234
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 68468 56151 68520 56160
rect 68468 56117 68477 56151
rect 68477 56117 68511 56151
rect 68511 56117 68520 56151
rect 68468 56108 68520 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 1768 46563 1820 46572
rect 1768 46529 1777 46563
rect 1777 46529 1811 46563
rect 1811 46529 1820 46563
rect 1768 46520 1820 46529
rect 940 46316 992 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 18236 37272 18288 37324
rect 940 37136 992 37188
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 21732 29112 21784 29164
rect 23940 29087 23992 29096
rect 23940 29053 23949 29087
rect 23949 29053 23983 29087
rect 23983 29053 23992 29087
rect 23940 29044 23992 29053
rect 21088 28951 21140 28960
rect 21088 28917 21097 28951
rect 21097 28917 21131 28951
rect 21131 28917 21140 28951
rect 21088 28908 21140 28917
rect 23296 28951 23348 28960
rect 23296 28917 23305 28951
rect 23305 28917 23339 28951
rect 23339 28917 23348 28951
rect 23296 28908 23348 28917
rect 23480 28908 23532 28960
rect 24860 28951 24912 28960
rect 24860 28917 24869 28951
rect 24869 28917 24903 28951
rect 24903 28917 24912 28951
rect 24860 28908 24912 28917
rect 25136 28908 25188 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 25412 28568 25464 28620
rect 17960 28364 18012 28416
rect 20352 28475 20404 28484
rect 20352 28441 20361 28475
rect 20361 28441 20395 28475
rect 20395 28441 20404 28475
rect 20352 28432 20404 28441
rect 21088 28432 21140 28484
rect 22100 28475 22152 28484
rect 22100 28441 22109 28475
rect 22109 28441 22143 28475
rect 22143 28441 22152 28475
rect 22100 28432 22152 28441
rect 22468 28475 22520 28484
rect 22468 28441 22477 28475
rect 22477 28441 22511 28475
rect 22511 28441 22520 28475
rect 22468 28432 22520 28441
rect 23480 28432 23532 28484
rect 24676 28475 24728 28484
rect 24676 28441 24685 28475
rect 24685 28441 24719 28475
rect 24719 28441 24728 28475
rect 24676 28432 24728 28441
rect 25136 28432 25188 28484
rect 25964 28432 26016 28484
rect 23940 28407 23992 28416
rect 23940 28373 23949 28407
rect 23949 28373 23983 28407
rect 23983 28373 23992 28407
rect 23940 28364 23992 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 20352 28160 20404 28212
rect 22468 28160 22520 28212
rect 21180 28067 21232 28076
rect 21180 28033 21189 28067
rect 21189 28033 21223 28067
rect 21223 28033 21232 28067
rect 21180 28024 21232 28033
rect 22100 27956 22152 28008
rect 22376 28067 22428 28076
rect 22376 28033 22385 28067
rect 22385 28033 22419 28067
rect 22419 28033 22428 28067
rect 22376 28024 22428 28033
rect 22468 28067 22520 28076
rect 22468 28033 22477 28067
rect 22477 28033 22511 28067
rect 22511 28033 22520 28067
rect 22468 28024 22520 28033
rect 22560 28067 22612 28076
rect 22560 28033 22569 28067
rect 22569 28033 22603 28067
rect 22603 28033 22612 28067
rect 22560 28024 22612 28033
rect 24860 28092 24912 28144
rect 25412 28092 25464 28144
rect 23296 28024 23348 28076
rect 68836 28024 68888 28076
rect 22652 27956 22704 28008
rect 25044 27956 25096 28008
rect 23572 27820 23624 27872
rect 23756 27863 23808 27872
rect 23756 27829 23765 27863
rect 23765 27829 23799 27863
rect 23799 27829 23808 27863
rect 23756 27820 23808 27829
rect 68284 27863 68336 27872
rect 68284 27829 68293 27863
rect 68293 27829 68327 27863
rect 68327 27829 68336 27863
rect 68284 27820 68336 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 22376 27616 22428 27668
rect 25044 27659 25096 27668
rect 25044 27625 25053 27659
rect 25053 27625 25087 27659
rect 25087 27625 25096 27659
rect 25044 27616 25096 27625
rect 22652 27548 22704 27600
rect 24216 27548 24268 27600
rect 22100 27480 22152 27532
rect 22928 27480 22980 27532
rect 23756 27480 23808 27532
rect 25412 27548 25464 27600
rect 20996 27455 21048 27464
rect 20996 27421 21005 27455
rect 21005 27421 21039 27455
rect 21039 27421 21048 27455
rect 20996 27412 21048 27421
rect 23388 27455 23440 27464
rect 23388 27421 23397 27455
rect 23397 27421 23431 27455
rect 23431 27421 23440 27455
rect 23388 27412 23440 27421
rect 23572 27412 23624 27464
rect 23296 27344 23348 27396
rect 23940 27344 23992 27396
rect 20628 27276 20680 27328
rect 21272 27276 21324 27328
rect 21640 27276 21692 27328
rect 22560 27276 22612 27328
rect 23020 27276 23072 27328
rect 24768 27387 24820 27396
rect 24768 27353 24777 27387
rect 24777 27353 24811 27387
rect 24811 27353 24820 27387
rect 24768 27344 24820 27353
rect 25044 27344 25096 27396
rect 25320 27455 25372 27464
rect 25320 27421 25329 27455
rect 25329 27421 25363 27455
rect 25363 27421 25372 27455
rect 25320 27412 25372 27421
rect 25412 27455 25464 27464
rect 25412 27421 25421 27455
rect 25421 27421 25455 27455
rect 25455 27421 25464 27455
rect 25412 27412 25464 27421
rect 26056 27412 26108 27464
rect 26608 27344 26660 27396
rect 28632 27344 28684 27396
rect 30564 27412 30616 27464
rect 25780 27276 25832 27328
rect 27712 27276 27764 27328
rect 29368 27319 29420 27328
rect 29368 27285 29377 27319
rect 29377 27285 29411 27319
rect 29411 27285 29420 27319
rect 29368 27276 29420 27285
rect 29552 27319 29604 27328
rect 29552 27285 29561 27319
rect 29561 27285 29595 27319
rect 29595 27285 29604 27319
rect 29552 27276 29604 27285
rect 30288 27319 30340 27328
rect 30288 27285 30297 27319
rect 30297 27285 30331 27319
rect 30331 27285 30340 27319
rect 30288 27276 30340 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 20628 27072 20680 27124
rect 18788 27004 18840 27056
rect 17868 26979 17920 26988
rect 17868 26945 17877 26979
rect 17877 26945 17911 26979
rect 17911 26945 17920 26979
rect 17868 26936 17920 26945
rect 20812 26936 20864 26988
rect 19800 26868 19852 26920
rect 19708 26775 19760 26784
rect 19708 26741 19717 26775
rect 19717 26741 19751 26775
rect 19751 26741 19760 26775
rect 19708 26732 19760 26741
rect 20352 26911 20404 26920
rect 20352 26877 20361 26911
rect 20361 26877 20395 26911
rect 20395 26877 20404 26911
rect 20352 26868 20404 26877
rect 20996 27072 21048 27124
rect 21272 27072 21324 27124
rect 22468 27072 22520 27124
rect 22744 27072 22796 27124
rect 22928 27072 22980 27124
rect 23296 27072 23348 27124
rect 21640 27047 21692 27056
rect 21640 27013 21649 27047
rect 21649 27013 21683 27047
rect 21683 27013 21692 27047
rect 21640 27004 21692 27013
rect 23572 27004 23624 27056
rect 20444 26800 20496 26852
rect 20260 26732 20312 26784
rect 20536 26775 20588 26784
rect 20536 26741 20545 26775
rect 20545 26741 20579 26775
rect 20579 26741 20588 26775
rect 20536 26732 20588 26741
rect 22836 26936 22888 26988
rect 23480 26979 23532 26988
rect 23480 26945 23489 26979
rect 23489 26945 23523 26979
rect 23523 26945 23532 26979
rect 23480 26936 23532 26945
rect 22652 26868 22704 26920
rect 22928 26800 22980 26852
rect 23388 26843 23440 26852
rect 23388 26809 23397 26843
rect 23397 26809 23431 26843
rect 23431 26809 23440 26843
rect 23388 26800 23440 26809
rect 22836 26775 22888 26784
rect 22836 26741 22845 26775
rect 22845 26741 22879 26775
rect 22879 26741 22888 26775
rect 22836 26732 22888 26741
rect 23664 26868 23716 26920
rect 24676 27115 24728 27124
rect 24676 27081 24685 27115
rect 24685 27081 24719 27115
rect 24719 27081 24728 27115
rect 24676 27072 24728 27081
rect 24768 27115 24820 27124
rect 24768 27081 24777 27115
rect 24777 27081 24811 27115
rect 24811 27081 24820 27115
rect 24768 27072 24820 27081
rect 26608 27072 26660 27124
rect 28632 27115 28684 27124
rect 28632 27081 28641 27115
rect 28641 27081 28675 27115
rect 28675 27081 28684 27115
rect 28632 27072 28684 27081
rect 29552 27072 29604 27124
rect 30288 27072 30340 27124
rect 24216 27047 24268 27056
rect 24216 27013 24233 27047
rect 24233 27013 24268 27047
rect 24216 27004 24268 27013
rect 25504 27004 25556 27056
rect 25964 27004 26016 27056
rect 24308 26979 24360 26988
rect 24308 26945 24317 26979
rect 24317 26945 24351 26979
rect 24351 26945 24360 26979
rect 24308 26936 24360 26945
rect 25044 26936 25096 26988
rect 25596 26979 25648 26988
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 23848 26775 23900 26784
rect 23848 26741 23857 26775
rect 23857 26741 23891 26775
rect 23891 26741 23900 26775
rect 23848 26732 23900 26741
rect 25320 26868 25372 26920
rect 25504 26800 25556 26852
rect 27160 26868 27212 26920
rect 27436 26868 27488 26920
rect 27712 26979 27764 26988
rect 27712 26945 27721 26979
rect 27721 26945 27755 26979
rect 27755 26945 27764 26979
rect 27712 26936 27764 26945
rect 28816 26979 28868 26988
rect 28816 26945 28825 26979
rect 28825 26945 28859 26979
rect 28859 26945 28868 26979
rect 28816 26936 28868 26945
rect 32956 27004 33008 27056
rect 32404 26936 32456 26988
rect 29736 26732 29788 26784
rect 30288 26732 30340 26784
rect 31484 26732 31536 26784
rect 33784 26732 33836 26784
rect 34060 26775 34112 26784
rect 34060 26741 34069 26775
rect 34069 26741 34103 26775
rect 34103 26741 34112 26775
rect 34060 26732 34112 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 18328 26528 18380 26580
rect 18788 26571 18840 26580
rect 18788 26537 18797 26571
rect 18797 26537 18831 26571
rect 18831 26537 18840 26571
rect 18788 26528 18840 26537
rect 19708 26528 19760 26580
rect 19800 26571 19852 26580
rect 19800 26537 19809 26571
rect 19809 26537 19843 26571
rect 19843 26537 19852 26571
rect 19800 26528 19852 26537
rect 19340 26460 19392 26512
rect 10416 26256 10468 26308
rect 12440 26299 12492 26308
rect 12440 26265 12449 26299
rect 12449 26265 12483 26299
rect 12483 26265 12492 26299
rect 12440 26256 12492 26265
rect 18236 26367 18288 26376
rect 18236 26333 18245 26367
rect 18245 26333 18279 26367
rect 18279 26333 18288 26367
rect 18236 26324 18288 26333
rect 20444 26528 20496 26580
rect 20536 26528 20588 26580
rect 20812 26528 20864 26580
rect 21640 26528 21692 26580
rect 22744 26571 22796 26580
rect 22744 26537 22753 26571
rect 22753 26537 22787 26571
rect 22787 26537 22796 26571
rect 22744 26528 22796 26537
rect 23480 26528 23532 26580
rect 25504 26528 25556 26580
rect 27436 26571 27488 26580
rect 27436 26537 27445 26571
rect 27445 26537 27479 26571
rect 27479 26537 27488 26571
rect 27436 26528 27488 26537
rect 27712 26528 27764 26580
rect 28540 26571 28592 26580
rect 28540 26537 28549 26571
rect 28549 26537 28583 26571
rect 28583 26537 28592 26571
rect 28540 26528 28592 26537
rect 28816 26528 28868 26580
rect 23296 26460 23348 26512
rect 20260 26367 20312 26376
rect 20260 26333 20269 26367
rect 20269 26333 20303 26367
rect 20303 26333 20312 26367
rect 21180 26392 21232 26444
rect 21272 26392 21324 26444
rect 20260 26324 20312 26333
rect 21548 26367 21600 26376
rect 21548 26333 21557 26367
rect 21557 26333 21591 26367
rect 21591 26333 21600 26367
rect 21548 26324 21600 26333
rect 21640 26324 21692 26376
rect 20076 26256 20128 26308
rect 13820 26188 13872 26240
rect 13912 26231 13964 26240
rect 13912 26197 13921 26231
rect 13921 26197 13955 26231
rect 13955 26197 13964 26231
rect 13912 26188 13964 26197
rect 16212 26188 16264 26240
rect 19432 26188 19484 26240
rect 22008 26367 22060 26376
rect 22008 26333 22017 26367
rect 22017 26333 22051 26367
rect 22051 26333 22060 26367
rect 22008 26324 22060 26333
rect 22192 26324 22244 26376
rect 23664 26392 23716 26444
rect 25412 26435 25464 26444
rect 25412 26401 25421 26435
rect 25421 26401 25455 26435
rect 25455 26401 25464 26435
rect 25412 26392 25464 26401
rect 22468 26256 22520 26308
rect 22744 26256 22796 26308
rect 25320 26324 25372 26376
rect 25596 26324 25648 26376
rect 27068 26324 27120 26376
rect 27804 26324 27856 26376
rect 29736 26367 29788 26376
rect 29736 26333 29745 26367
rect 29745 26333 29779 26367
rect 29779 26333 29788 26367
rect 29736 26324 29788 26333
rect 30472 26392 30524 26444
rect 34060 26528 34112 26580
rect 31484 26367 31536 26376
rect 28080 26256 28132 26308
rect 29368 26256 29420 26308
rect 21824 26188 21876 26240
rect 23112 26188 23164 26240
rect 24952 26231 25004 26240
rect 24952 26197 24961 26231
rect 24961 26197 24995 26231
rect 24995 26197 25004 26231
rect 24952 26188 25004 26197
rect 27712 26188 27764 26240
rect 27896 26188 27948 26240
rect 28724 26231 28776 26240
rect 28724 26197 28733 26231
rect 28733 26197 28767 26231
rect 28767 26197 28776 26231
rect 28724 26188 28776 26197
rect 29276 26188 29328 26240
rect 31484 26333 31493 26367
rect 31493 26333 31527 26367
rect 31527 26333 31536 26367
rect 31484 26324 31536 26333
rect 31760 26367 31812 26376
rect 31760 26333 31769 26367
rect 31769 26333 31803 26367
rect 31803 26333 31812 26367
rect 31760 26324 31812 26333
rect 32404 26435 32456 26444
rect 32404 26401 32413 26435
rect 32413 26401 32447 26435
rect 32447 26401 32456 26435
rect 32404 26392 32456 26401
rect 32956 26435 33008 26444
rect 32956 26401 32965 26435
rect 32965 26401 32999 26435
rect 32999 26401 33008 26435
rect 32956 26392 33008 26401
rect 33048 26435 33100 26444
rect 33048 26401 33057 26435
rect 33057 26401 33091 26435
rect 33091 26401 33100 26435
rect 33048 26392 33100 26401
rect 33876 26392 33928 26444
rect 30748 26299 30800 26308
rect 30748 26265 30757 26299
rect 30757 26265 30791 26299
rect 30791 26265 30800 26299
rect 30748 26256 30800 26265
rect 30932 26256 30984 26308
rect 30472 26188 30524 26240
rect 31208 26188 31260 26240
rect 32680 26324 32732 26376
rect 32864 26367 32916 26376
rect 32864 26333 32873 26367
rect 32873 26333 32907 26367
rect 32907 26333 32916 26367
rect 32864 26324 32916 26333
rect 31760 26188 31812 26240
rect 32220 26188 32272 26240
rect 32680 26188 32732 26240
rect 33324 26299 33376 26308
rect 33324 26265 33333 26299
rect 33333 26265 33367 26299
rect 33367 26265 33376 26299
rect 33324 26256 33376 26265
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 16304 25916 16356 25968
rect 19340 25984 19392 26036
rect 19432 25916 19484 25968
rect 21180 26027 21232 26036
rect 21180 25993 21189 26027
rect 21189 25993 21223 26027
rect 21223 25993 21232 26027
rect 21180 25984 21232 25993
rect 21548 25984 21600 26036
rect 22008 25984 22060 26036
rect 22652 26027 22704 26036
rect 22652 25993 22661 26027
rect 22661 25993 22695 26027
rect 22695 25993 22704 26027
rect 22652 25984 22704 25993
rect 25504 25984 25556 26036
rect 28540 25984 28592 26036
rect 30472 25984 30524 26036
rect 20352 25916 20404 25968
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 13820 25848 13872 25900
rect 17960 25848 18012 25900
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 12808 25823 12860 25832
rect 12808 25789 12817 25823
rect 12817 25789 12851 25823
rect 12851 25789 12860 25823
rect 12808 25780 12860 25789
rect 13912 25780 13964 25832
rect 14280 25823 14332 25832
rect 14280 25789 14289 25823
rect 14289 25789 14323 25823
rect 14323 25789 14332 25823
rect 14280 25780 14332 25789
rect 21548 25891 21600 25900
rect 21548 25857 21557 25891
rect 21557 25857 21591 25891
rect 21591 25857 21600 25891
rect 21548 25848 21600 25857
rect 21824 25891 21876 25900
rect 21824 25857 21833 25891
rect 21833 25857 21867 25891
rect 21867 25857 21876 25891
rect 21824 25848 21876 25857
rect 21916 25848 21968 25900
rect 12440 25712 12492 25764
rect 22100 25848 22152 25900
rect 22744 25891 22796 25900
rect 22744 25857 22753 25891
rect 22753 25857 22787 25891
rect 22787 25857 22796 25891
rect 22744 25848 22796 25857
rect 23848 25848 23900 25900
rect 24768 25891 24820 25900
rect 24768 25857 24777 25891
rect 24777 25857 24811 25891
rect 24811 25857 24820 25891
rect 24768 25848 24820 25857
rect 24952 25891 25004 25900
rect 24952 25857 24961 25891
rect 24961 25857 24995 25891
rect 24995 25857 25004 25891
rect 24952 25848 25004 25857
rect 25136 25891 25188 25900
rect 25136 25857 25145 25891
rect 25145 25857 25179 25891
rect 25179 25857 25188 25891
rect 25136 25848 25188 25857
rect 27068 25916 27120 25968
rect 26240 25848 26292 25900
rect 25044 25823 25096 25832
rect 25044 25789 25053 25823
rect 25053 25789 25087 25823
rect 25087 25789 25096 25823
rect 25044 25780 25096 25789
rect 25320 25780 25372 25832
rect 15752 25687 15804 25696
rect 15752 25653 15761 25687
rect 15761 25653 15795 25687
rect 15795 25653 15804 25687
rect 15752 25644 15804 25653
rect 22192 25644 22244 25696
rect 25596 25755 25648 25764
rect 25596 25721 25605 25755
rect 25605 25721 25639 25755
rect 25639 25721 25648 25755
rect 25596 25712 25648 25721
rect 27436 25848 27488 25900
rect 27620 25891 27672 25900
rect 27620 25857 27629 25891
rect 27629 25857 27663 25891
rect 27663 25857 27672 25891
rect 27620 25848 27672 25857
rect 27712 25891 27764 25900
rect 27712 25857 27721 25891
rect 27721 25857 27755 25891
rect 27755 25857 27764 25891
rect 27712 25848 27764 25857
rect 27896 25848 27948 25900
rect 29184 25891 29236 25900
rect 29184 25857 29193 25891
rect 29193 25857 29227 25891
rect 29227 25857 29236 25891
rect 29184 25848 29236 25857
rect 31208 25891 31260 25900
rect 31208 25857 31217 25891
rect 31217 25857 31251 25891
rect 31251 25857 31260 25891
rect 31208 25848 31260 25857
rect 31484 25848 31536 25900
rect 29920 25823 29972 25832
rect 29920 25789 29929 25823
rect 29929 25789 29963 25823
rect 29963 25789 29972 25823
rect 29920 25780 29972 25789
rect 30564 25780 30616 25832
rect 31116 25823 31168 25832
rect 31116 25789 31125 25823
rect 31125 25789 31159 25823
rect 31159 25789 31168 25823
rect 31116 25780 31168 25789
rect 27160 25712 27212 25764
rect 23204 25644 23256 25696
rect 24032 25644 24084 25696
rect 25320 25687 25372 25696
rect 25320 25653 25329 25687
rect 25329 25653 25363 25687
rect 25363 25653 25372 25687
rect 25320 25644 25372 25653
rect 26700 25687 26752 25696
rect 26700 25653 26709 25687
rect 26709 25653 26743 25687
rect 26743 25653 26752 25687
rect 26700 25644 26752 25653
rect 27804 25644 27856 25696
rect 28816 25712 28868 25764
rect 29276 25644 29328 25696
rect 29368 25687 29420 25696
rect 29368 25653 29377 25687
rect 29377 25653 29411 25687
rect 29411 25653 29420 25687
rect 29368 25644 29420 25653
rect 30656 25644 30708 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 12716 25440 12768 25492
rect 14280 25440 14332 25492
rect 16304 25483 16356 25492
rect 16304 25449 16313 25483
rect 16313 25449 16347 25483
rect 16347 25449 16356 25483
rect 16304 25440 16356 25449
rect 12624 25372 12676 25424
rect 9772 25304 9824 25356
rect 10416 25304 10468 25356
rect 10968 25304 11020 25356
rect 13360 25279 13412 25288
rect 13360 25245 13369 25279
rect 13369 25245 13403 25279
rect 13403 25245 13412 25279
rect 13360 25236 13412 25245
rect 14004 25304 14056 25356
rect 13912 25236 13964 25288
rect 15752 25304 15804 25356
rect 17960 25304 18012 25356
rect 19064 25304 19116 25356
rect 16028 25279 16080 25288
rect 16028 25245 16037 25279
rect 16037 25245 16071 25279
rect 16071 25245 16080 25279
rect 16028 25236 16080 25245
rect 11152 25168 11204 25220
rect 16672 25279 16724 25288
rect 16672 25245 16681 25279
rect 16681 25245 16715 25279
rect 16715 25245 16724 25279
rect 16672 25236 16724 25245
rect 18696 25279 18748 25288
rect 18696 25245 18705 25279
rect 18705 25245 18739 25279
rect 18739 25245 18748 25279
rect 18696 25236 18748 25245
rect 22836 25440 22888 25492
rect 23296 25440 23348 25492
rect 23572 25483 23624 25492
rect 23572 25449 23581 25483
rect 23581 25449 23615 25483
rect 23615 25449 23624 25483
rect 23572 25440 23624 25449
rect 24768 25440 24820 25492
rect 27620 25440 27672 25492
rect 29276 25483 29328 25492
rect 29276 25449 29285 25483
rect 29285 25449 29319 25483
rect 29319 25449 29328 25483
rect 29276 25440 29328 25449
rect 29368 25440 29420 25492
rect 22284 25304 22336 25356
rect 22744 25372 22796 25424
rect 16212 25168 16264 25220
rect 16580 25168 16632 25220
rect 17960 25168 18012 25220
rect 19432 25168 19484 25220
rect 19984 25168 20036 25220
rect 21456 25168 21508 25220
rect 11980 25100 12032 25152
rect 12164 25143 12216 25152
rect 12164 25109 12173 25143
rect 12173 25109 12207 25143
rect 12207 25109 12216 25143
rect 12164 25100 12216 25109
rect 12440 25100 12492 25152
rect 16488 25100 16540 25152
rect 18052 25143 18104 25152
rect 18052 25109 18061 25143
rect 18061 25109 18095 25143
rect 18095 25109 18104 25143
rect 18052 25100 18104 25109
rect 20812 25100 20864 25152
rect 22560 25211 22612 25220
rect 22560 25177 22569 25211
rect 22569 25177 22603 25211
rect 22603 25177 22612 25211
rect 22560 25168 22612 25177
rect 22652 25211 22704 25220
rect 22652 25177 22661 25211
rect 22661 25177 22695 25211
rect 22695 25177 22704 25211
rect 22652 25168 22704 25177
rect 23296 25279 23348 25288
rect 23296 25245 23305 25279
rect 23305 25245 23339 25279
rect 23339 25245 23348 25279
rect 23296 25236 23348 25245
rect 24216 25236 24268 25288
rect 27896 25372 27948 25424
rect 24860 25304 24912 25356
rect 26056 25347 26108 25356
rect 26056 25313 26065 25347
rect 26065 25313 26099 25347
rect 26099 25313 26108 25347
rect 26056 25304 26108 25313
rect 27712 25347 27764 25356
rect 27712 25313 27721 25347
rect 27721 25313 27755 25347
rect 27755 25313 27764 25347
rect 27712 25304 27764 25313
rect 28080 25304 28132 25356
rect 25044 25236 25096 25288
rect 25320 25279 25372 25288
rect 25320 25245 25324 25279
rect 25324 25245 25358 25279
rect 25358 25245 25372 25279
rect 25320 25236 25372 25245
rect 25596 25279 25648 25288
rect 25596 25245 25641 25279
rect 25641 25245 25648 25279
rect 25596 25236 25648 25245
rect 25780 25279 25832 25288
rect 25780 25245 25789 25279
rect 25789 25245 25823 25279
rect 25823 25245 25832 25279
rect 25780 25236 25832 25245
rect 26700 25236 26752 25288
rect 27804 25279 27856 25288
rect 27804 25245 27813 25279
rect 27813 25245 27847 25279
rect 27847 25245 27856 25279
rect 27804 25236 27856 25245
rect 28724 25304 28776 25356
rect 23020 25100 23072 25152
rect 23664 25211 23716 25220
rect 23664 25177 23673 25211
rect 23673 25177 23707 25211
rect 23707 25177 23716 25211
rect 23664 25168 23716 25177
rect 25412 25211 25464 25220
rect 25412 25177 25421 25211
rect 25421 25177 25455 25211
rect 25455 25177 25464 25211
rect 25412 25168 25464 25177
rect 25504 25211 25556 25220
rect 25504 25177 25513 25211
rect 25513 25177 25547 25211
rect 25547 25177 25556 25211
rect 25504 25168 25556 25177
rect 28816 25279 28868 25288
rect 28816 25245 28825 25279
rect 28825 25245 28859 25279
rect 28859 25245 28868 25279
rect 28816 25236 28868 25245
rect 30932 25372 30984 25424
rect 30380 25236 30432 25288
rect 31208 25279 31260 25288
rect 31208 25245 31217 25279
rect 31217 25245 31251 25279
rect 31251 25245 31260 25279
rect 31208 25236 31260 25245
rect 33784 25236 33836 25288
rect 35532 25236 35584 25288
rect 37280 25236 37332 25288
rect 27712 25100 27764 25152
rect 29092 25100 29144 25152
rect 31484 25211 31536 25220
rect 31484 25177 31493 25211
rect 31493 25177 31527 25211
rect 31527 25177 31536 25211
rect 31484 25168 31536 25177
rect 31852 25168 31904 25220
rect 30748 25100 30800 25152
rect 31760 25100 31812 25152
rect 33324 25168 33376 25220
rect 32128 25143 32180 25152
rect 32128 25109 32153 25143
rect 32153 25109 32180 25143
rect 32128 25100 32180 25109
rect 32312 25143 32364 25152
rect 32312 25109 32321 25143
rect 32321 25109 32355 25143
rect 32355 25109 32364 25143
rect 32312 25100 32364 25109
rect 36176 25143 36228 25152
rect 36176 25109 36185 25143
rect 36185 25109 36219 25143
rect 36219 25109 36228 25143
rect 36176 25100 36228 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 11152 24939 11204 24948
rect 11152 24905 11161 24939
rect 11161 24905 11195 24939
rect 11195 24905 11204 24939
rect 11152 24896 11204 24905
rect 11980 24939 12032 24948
rect 11980 24905 11989 24939
rect 11989 24905 12023 24939
rect 12023 24905 12032 24939
rect 11980 24896 12032 24905
rect 12164 24896 12216 24948
rect 14004 24896 14056 24948
rect 16028 24896 16080 24948
rect 16580 24896 16632 24948
rect 16672 24896 16724 24948
rect 19432 24939 19484 24948
rect 19432 24905 19441 24939
rect 19441 24905 19475 24939
rect 19475 24905 19484 24939
rect 19432 24896 19484 24905
rect 19984 24896 20036 24948
rect 22560 24896 22612 24948
rect 22652 24896 22704 24948
rect 23112 24896 23164 24948
rect 9312 24828 9364 24880
rect 10140 24760 10192 24812
rect 11244 24828 11296 24880
rect 11152 24760 11204 24812
rect 7932 24556 7984 24608
rect 9864 24692 9916 24744
rect 11520 24692 11572 24744
rect 9588 24624 9640 24676
rect 10784 24556 10836 24608
rect 11980 24556 12032 24608
rect 12808 24828 12860 24880
rect 13820 24760 13872 24812
rect 14280 24803 14332 24812
rect 14280 24769 14314 24803
rect 14314 24769 14332 24803
rect 14280 24760 14332 24769
rect 16304 24803 16356 24812
rect 16304 24769 16313 24803
rect 16313 24769 16347 24803
rect 16347 24769 16356 24803
rect 16304 24760 16356 24769
rect 24952 24896 25004 24948
rect 25412 24939 25464 24948
rect 25412 24905 25421 24939
rect 25421 24905 25455 24939
rect 25455 24905 25464 24939
rect 25412 24896 25464 24905
rect 25504 24896 25556 24948
rect 29092 24896 29144 24948
rect 30748 24896 30800 24948
rect 31208 24896 31260 24948
rect 32220 24939 32272 24948
rect 32220 24905 32229 24939
rect 32229 24905 32263 24939
rect 32263 24905 32272 24939
rect 32220 24896 32272 24905
rect 32312 24896 32364 24948
rect 33324 24896 33376 24948
rect 16764 24760 16816 24812
rect 18052 24760 18104 24812
rect 19248 24803 19300 24812
rect 19248 24769 19257 24803
rect 19257 24769 19291 24803
rect 19291 24769 19300 24803
rect 19248 24760 19300 24769
rect 20812 24760 20864 24812
rect 21548 24760 21600 24812
rect 21732 24760 21784 24812
rect 22100 24760 22152 24812
rect 12624 24556 12676 24608
rect 12900 24599 12952 24608
rect 12900 24565 12909 24599
rect 12909 24565 12943 24599
rect 12943 24565 12952 24599
rect 12900 24556 12952 24565
rect 20168 24692 20220 24744
rect 20536 24735 20588 24744
rect 20536 24701 20545 24735
rect 20545 24701 20579 24735
rect 20579 24701 20588 24735
rect 20536 24692 20588 24701
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 23572 24828 23624 24880
rect 24584 24828 24636 24880
rect 22376 24760 22428 24769
rect 25780 24803 25832 24812
rect 25780 24769 25789 24803
rect 25789 24769 25823 24803
rect 25823 24769 25832 24803
rect 25780 24760 25832 24769
rect 27620 24760 27672 24812
rect 28080 24760 28132 24812
rect 31852 24828 31904 24880
rect 28724 24760 28776 24812
rect 30656 24760 30708 24812
rect 30932 24760 30984 24812
rect 15752 24624 15804 24676
rect 16672 24556 16724 24608
rect 18696 24624 18748 24676
rect 23572 24667 23624 24676
rect 23572 24633 23581 24667
rect 23581 24633 23615 24667
rect 23615 24633 23624 24667
rect 23572 24624 23624 24633
rect 18144 24599 18196 24608
rect 18144 24565 18153 24599
rect 18153 24565 18187 24599
rect 18187 24565 18196 24599
rect 18144 24556 18196 24565
rect 19892 24599 19944 24608
rect 19892 24565 19901 24599
rect 19901 24565 19935 24599
rect 19935 24565 19944 24599
rect 19892 24556 19944 24565
rect 20720 24556 20772 24608
rect 21916 24599 21968 24608
rect 21916 24565 21925 24599
rect 21925 24565 21959 24599
rect 21959 24565 21968 24599
rect 21916 24556 21968 24565
rect 23296 24556 23348 24608
rect 28172 24692 28224 24744
rect 31116 24692 31168 24744
rect 29184 24624 29236 24676
rect 32220 24760 32272 24812
rect 32496 24803 32548 24812
rect 32496 24769 32505 24803
rect 32505 24769 32539 24803
rect 32539 24769 32548 24803
rect 32496 24760 32548 24769
rect 32588 24803 32640 24812
rect 32588 24769 32597 24803
rect 32597 24769 32631 24803
rect 32631 24769 32640 24803
rect 32588 24760 32640 24769
rect 33784 24760 33836 24812
rect 34336 24760 34388 24812
rect 34520 24803 34572 24812
rect 34520 24769 34554 24803
rect 34554 24769 34572 24803
rect 34520 24760 34572 24769
rect 36176 24828 36228 24880
rect 31852 24692 31904 24744
rect 32588 24624 32640 24676
rect 24676 24556 24728 24608
rect 28080 24599 28132 24608
rect 28080 24565 28089 24599
rect 28089 24565 28123 24599
rect 28123 24565 28132 24599
rect 28080 24556 28132 24565
rect 29552 24599 29604 24608
rect 29552 24565 29561 24599
rect 29561 24565 29595 24599
rect 29595 24565 29604 24599
rect 29552 24556 29604 24565
rect 31760 24556 31812 24608
rect 32496 24556 32548 24608
rect 35992 24556 36044 24608
rect 36084 24556 36136 24608
rect 37924 24599 37976 24608
rect 37924 24565 37933 24599
rect 37933 24565 37967 24599
rect 37967 24565 37976 24599
rect 37924 24556 37976 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 9312 24352 9364 24404
rect 9864 24352 9916 24404
rect 12808 24352 12860 24404
rect 12900 24352 12952 24404
rect 14004 24352 14056 24404
rect 14280 24352 14332 24404
rect 16764 24352 16816 24404
rect 18144 24352 18196 24404
rect 19248 24352 19300 24404
rect 10324 24284 10376 24336
rect 9956 24191 10008 24200
rect 9956 24157 9965 24191
rect 9965 24157 9999 24191
rect 9999 24157 10008 24191
rect 9956 24148 10008 24157
rect 10508 24148 10560 24200
rect 8852 24012 8904 24064
rect 10600 24055 10652 24064
rect 10600 24021 10609 24055
rect 10609 24021 10643 24055
rect 10643 24021 10652 24055
rect 10600 24012 10652 24021
rect 10784 24080 10836 24132
rect 11244 24191 11296 24200
rect 11244 24157 11253 24191
rect 11253 24157 11287 24191
rect 11287 24157 11296 24191
rect 11244 24148 11296 24157
rect 11336 24191 11388 24200
rect 11336 24157 11345 24191
rect 11345 24157 11379 24191
rect 11379 24157 11388 24191
rect 11336 24148 11388 24157
rect 11520 24191 11572 24200
rect 11520 24157 11529 24191
rect 11529 24157 11563 24191
rect 11563 24157 11572 24191
rect 11520 24148 11572 24157
rect 12624 24216 12676 24268
rect 13084 24191 13136 24200
rect 13084 24157 13093 24191
rect 13093 24157 13127 24191
rect 13127 24157 13136 24191
rect 13084 24148 13136 24157
rect 15752 24216 15804 24268
rect 11152 24012 11204 24064
rect 11244 24012 11296 24064
rect 12900 24123 12952 24132
rect 12900 24089 12909 24123
rect 12909 24089 12943 24123
rect 12943 24089 12952 24123
rect 12900 24080 12952 24089
rect 15936 24148 15988 24200
rect 16580 24191 16632 24200
rect 16580 24157 16589 24191
rect 16589 24157 16623 24191
rect 16623 24157 16632 24191
rect 16580 24148 16632 24157
rect 19064 24259 19116 24268
rect 19064 24225 19073 24259
rect 19073 24225 19107 24259
rect 19107 24225 19116 24259
rect 19064 24216 19116 24225
rect 20812 24352 20864 24404
rect 21916 24284 21968 24336
rect 22192 24284 22244 24336
rect 24584 24352 24636 24404
rect 30564 24395 30616 24404
rect 30564 24361 30573 24395
rect 30573 24361 30607 24395
rect 30607 24361 30616 24395
rect 30564 24352 30616 24361
rect 30932 24352 30984 24404
rect 32128 24352 32180 24404
rect 29920 24284 29972 24336
rect 33140 24352 33192 24404
rect 34520 24352 34572 24404
rect 37280 24395 37332 24404
rect 37280 24361 37289 24395
rect 37289 24361 37323 24395
rect 37323 24361 37332 24395
rect 37280 24352 37332 24361
rect 37924 24352 37976 24404
rect 21456 24216 21508 24268
rect 17500 24080 17552 24132
rect 18512 24080 18564 24132
rect 19892 24080 19944 24132
rect 13176 24012 13228 24064
rect 14740 24055 14792 24064
rect 14740 24021 14749 24055
rect 14749 24021 14783 24055
rect 14783 24021 14792 24055
rect 14740 24012 14792 24021
rect 15384 24012 15436 24064
rect 16672 24055 16724 24064
rect 16672 24021 16681 24055
rect 16681 24021 16715 24055
rect 16715 24021 16724 24055
rect 16672 24012 16724 24021
rect 17224 24012 17276 24064
rect 20076 24055 20128 24064
rect 20076 24021 20085 24055
rect 20085 24021 20119 24055
rect 20119 24021 20128 24055
rect 20076 24012 20128 24021
rect 21732 24012 21784 24064
rect 22192 24148 22244 24200
rect 22652 24191 22704 24200
rect 22652 24157 22661 24191
rect 22661 24157 22695 24191
rect 22695 24157 22704 24191
rect 22652 24148 22704 24157
rect 27620 24216 27672 24268
rect 28080 24216 28132 24268
rect 29276 24216 29328 24268
rect 31852 24216 31904 24268
rect 22284 24123 22336 24132
rect 22284 24089 22293 24123
rect 22293 24089 22327 24123
rect 22327 24089 22336 24123
rect 22284 24080 22336 24089
rect 25688 24148 25740 24200
rect 27344 24191 27396 24200
rect 27344 24157 27353 24191
rect 27353 24157 27387 24191
rect 27387 24157 27396 24191
rect 27344 24148 27396 24157
rect 27988 24148 28040 24200
rect 28172 24148 28224 24200
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 32496 24216 32548 24268
rect 30196 24148 30248 24200
rect 32220 24191 32272 24200
rect 32220 24157 32229 24191
rect 32229 24157 32263 24191
rect 32263 24157 32272 24191
rect 32220 24148 32272 24157
rect 32312 24148 32364 24200
rect 32864 24191 32916 24200
rect 32864 24157 32873 24191
rect 32873 24157 32907 24191
rect 32907 24157 32916 24191
rect 32864 24148 32916 24157
rect 32956 24191 33008 24200
rect 32956 24157 32965 24191
rect 32965 24157 32999 24191
rect 32999 24157 33008 24191
rect 32956 24148 33008 24157
rect 34336 24148 34388 24200
rect 35164 24191 35216 24200
rect 35164 24157 35173 24191
rect 35173 24157 35207 24191
rect 35207 24157 35216 24191
rect 35164 24148 35216 24157
rect 35532 24148 35584 24200
rect 35992 24148 36044 24200
rect 36360 24191 36412 24200
rect 36360 24157 36369 24191
rect 36369 24157 36403 24191
rect 36403 24157 36412 24191
rect 36360 24148 36412 24157
rect 37096 24148 37148 24200
rect 32588 24080 32640 24132
rect 34060 24080 34112 24132
rect 22928 24055 22980 24064
rect 22928 24021 22937 24055
rect 22937 24021 22971 24055
rect 22971 24021 22980 24055
rect 22928 24012 22980 24021
rect 25320 24055 25372 24064
rect 25320 24021 25329 24055
rect 25329 24021 25363 24055
rect 25363 24021 25372 24055
rect 25320 24012 25372 24021
rect 26976 24055 27028 24064
rect 26976 24021 26985 24055
rect 26985 24021 27019 24055
rect 27019 24021 27028 24055
rect 26976 24012 27028 24021
rect 27896 24055 27948 24064
rect 27896 24021 27905 24055
rect 27905 24021 27939 24055
rect 27939 24021 27948 24055
rect 27896 24012 27948 24021
rect 28540 24055 28592 24064
rect 28540 24021 28549 24055
rect 28549 24021 28583 24055
rect 28583 24021 28592 24055
rect 28540 24012 28592 24021
rect 32680 24055 32732 24064
rect 32680 24021 32689 24055
rect 32689 24021 32723 24055
rect 32723 24021 32732 24055
rect 32680 24012 32732 24021
rect 33048 24055 33100 24064
rect 33048 24021 33057 24055
rect 33057 24021 33091 24055
rect 33091 24021 33100 24055
rect 33048 24012 33100 24021
rect 36452 24055 36504 24064
rect 36452 24021 36461 24055
rect 36461 24021 36495 24055
rect 36495 24021 36504 24055
rect 36452 24012 36504 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 9956 23808 10008 23860
rect 10048 23808 10100 23860
rect 10508 23851 10560 23860
rect 10508 23817 10517 23851
rect 10517 23817 10551 23851
rect 10551 23817 10560 23851
rect 10508 23808 10560 23817
rect 10600 23808 10652 23860
rect 8944 23740 8996 23792
rect 11336 23808 11388 23860
rect 11980 23808 12032 23860
rect 11520 23783 11572 23792
rect 11520 23749 11529 23783
rect 11529 23749 11563 23783
rect 11563 23749 11572 23783
rect 11520 23740 11572 23749
rect 10324 23715 10376 23724
rect 10324 23681 10333 23715
rect 10333 23681 10367 23715
rect 10367 23681 10376 23715
rect 10324 23672 10376 23681
rect 10508 23672 10560 23724
rect 11060 23672 11112 23724
rect 7932 23647 7984 23656
rect 7932 23613 7941 23647
rect 7941 23613 7975 23647
rect 7975 23613 7984 23647
rect 7932 23604 7984 23613
rect 9956 23536 10008 23588
rect 11336 23715 11388 23724
rect 11336 23681 11345 23715
rect 11345 23681 11379 23715
rect 11379 23681 11388 23715
rect 12900 23851 12952 23860
rect 12900 23817 12909 23851
rect 12909 23817 12943 23851
rect 12943 23817 12952 23851
rect 12900 23808 12952 23817
rect 16304 23808 16356 23860
rect 17960 23808 18012 23860
rect 18512 23851 18564 23860
rect 18512 23817 18521 23851
rect 18521 23817 18555 23851
rect 18555 23817 18564 23851
rect 18512 23808 18564 23817
rect 20536 23808 20588 23860
rect 24308 23808 24360 23860
rect 25320 23808 25372 23860
rect 25688 23851 25740 23860
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 26976 23808 27028 23860
rect 27344 23808 27396 23860
rect 28172 23808 28224 23860
rect 28540 23808 28592 23860
rect 32680 23808 32732 23860
rect 13360 23740 13412 23792
rect 11336 23672 11388 23681
rect 12992 23672 13044 23724
rect 13084 23672 13136 23724
rect 12532 23647 12584 23656
rect 12532 23613 12541 23647
rect 12541 23613 12575 23647
rect 12575 23613 12584 23647
rect 12532 23604 12584 23613
rect 13268 23604 13320 23656
rect 17224 23604 17276 23656
rect 17500 23672 17552 23724
rect 16948 23536 17000 23588
rect 11612 23468 11664 23520
rect 14372 23468 14424 23520
rect 15936 23468 15988 23520
rect 18052 23715 18104 23724
rect 18052 23681 18061 23715
rect 18061 23681 18095 23715
rect 18095 23681 18104 23715
rect 18052 23672 18104 23681
rect 19064 23672 19116 23724
rect 18604 23604 18656 23656
rect 20260 23672 20312 23724
rect 18328 23536 18380 23588
rect 19432 23536 19484 23588
rect 22744 23715 22796 23724
rect 22744 23681 22753 23715
rect 22753 23681 22787 23715
rect 22787 23681 22796 23715
rect 22744 23672 22796 23681
rect 23388 23672 23440 23724
rect 22468 23604 22520 23656
rect 22652 23647 22704 23656
rect 22652 23613 22661 23647
rect 22661 23613 22695 23647
rect 22695 23613 22704 23647
rect 22652 23604 22704 23613
rect 22836 23604 22888 23656
rect 25044 23604 25096 23656
rect 25228 23604 25280 23656
rect 25780 23672 25832 23724
rect 26516 23715 26568 23724
rect 26516 23681 26525 23715
rect 26525 23681 26559 23715
rect 26559 23681 26568 23715
rect 26516 23672 26568 23681
rect 26884 23604 26936 23656
rect 32956 23740 33008 23792
rect 35164 23808 35216 23860
rect 34152 23715 34204 23724
rect 34152 23681 34161 23715
rect 34161 23681 34195 23715
rect 34195 23681 34204 23715
rect 34152 23672 34204 23681
rect 36268 23740 36320 23792
rect 36360 23672 36412 23724
rect 36544 23715 36596 23724
rect 36544 23681 36553 23715
rect 36553 23681 36587 23715
rect 36587 23681 36596 23715
rect 36544 23672 36596 23681
rect 37096 23672 37148 23724
rect 27712 23604 27764 23656
rect 29092 23647 29144 23656
rect 29092 23613 29101 23647
rect 29101 23613 29135 23647
rect 29135 23613 29144 23647
rect 29092 23604 29144 23613
rect 30564 23604 30616 23656
rect 30932 23604 30984 23656
rect 33048 23604 33100 23656
rect 33876 23604 33928 23656
rect 27160 23536 27212 23588
rect 27528 23536 27580 23588
rect 30196 23579 30248 23588
rect 30196 23545 30205 23579
rect 30205 23545 30239 23579
rect 30239 23545 30248 23579
rect 30196 23536 30248 23545
rect 32588 23536 32640 23588
rect 34060 23536 34112 23588
rect 36084 23647 36136 23656
rect 36084 23613 36093 23647
rect 36093 23613 36127 23647
rect 36127 23613 36136 23647
rect 36084 23604 36136 23613
rect 36728 23604 36780 23656
rect 36820 23647 36872 23656
rect 36820 23613 36829 23647
rect 36829 23613 36863 23647
rect 36863 23613 36872 23647
rect 36820 23604 36872 23613
rect 36360 23536 36412 23588
rect 36636 23579 36688 23588
rect 36636 23545 36645 23579
rect 36645 23545 36679 23579
rect 36679 23545 36688 23579
rect 36636 23536 36688 23545
rect 18420 23468 18472 23520
rect 19984 23468 20036 23520
rect 23296 23468 23348 23520
rect 24584 23468 24636 23520
rect 25596 23511 25648 23520
rect 25596 23477 25605 23511
rect 25605 23477 25639 23511
rect 25639 23477 25648 23511
rect 25596 23468 25648 23477
rect 26700 23511 26752 23520
rect 26700 23477 26709 23511
rect 26709 23477 26743 23511
rect 26743 23477 26752 23511
rect 26700 23468 26752 23477
rect 30472 23511 30524 23520
rect 30472 23477 30481 23511
rect 30481 23477 30515 23511
rect 30515 23477 30524 23511
rect 30472 23468 30524 23477
rect 37280 23468 37332 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 8944 23264 8996 23316
rect 11060 23264 11112 23316
rect 11612 23196 11664 23248
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 13176 23264 13228 23316
rect 14924 23264 14976 23316
rect 16580 23264 16632 23316
rect 16672 23196 16724 23248
rect 17132 23239 17184 23248
rect 17132 23205 17141 23239
rect 17141 23205 17175 23239
rect 17175 23205 17184 23239
rect 17132 23196 17184 23205
rect 11888 23128 11940 23180
rect 12532 23128 12584 23180
rect 12808 23103 12860 23112
rect 12808 23069 12817 23103
rect 12817 23069 12851 23103
rect 12851 23069 12860 23103
rect 12808 23060 12860 23069
rect 8852 22992 8904 23044
rect 10600 22992 10652 23044
rect 11336 23035 11388 23044
rect 10692 22967 10744 22976
rect 10692 22933 10701 22967
rect 10701 22933 10735 22967
rect 10735 22933 10744 22967
rect 10692 22924 10744 22933
rect 11336 23001 11363 23035
rect 11363 23001 11388 23035
rect 11336 22992 11388 23001
rect 11888 22992 11940 23044
rect 13820 23128 13872 23180
rect 14096 23128 14148 23180
rect 14556 23171 14608 23180
rect 14556 23137 14565 23171
rect 14565 23137 14599 23171
rect 14599 23137 14608 23171
rect 14556 23128 14608 23137
rect 13176 23103 13228 23112
rect 13176 23069 13185 23103
rect 13185 23069 13219 23103
rect 13219 23069 13228 23103
rect 13176 23060 13228 23069
rect 14372 23103 14424 23112
rect 14372 23069 14381 23103
rect 14381 23069 14415 23103
rect 14415 23069 14424 23103
rect 14372 23060 14424 23069
rect 15936 23060 15988 23112
rect 16120 23103 16172 23112
rect 16120 23069 16129 23103
rect 16129 23069 16163 23103
rect 16163 23069 16172 23103
rect 16120 23060 16172 23069
rect 17500 23171 17552 23180
rect 17500 23137 17509 23171
rect 17509 23137 17543 23171
rect 17543 23137 17552 23171
rect 17500 23128 17552 23137
rect 18052 23264 18104 23316
rect 20260 23264 20312 23316
rect 25228 23264 25280 23316
rect 25780 23264 25832 23316
rect 27712 23264 27764 23316
rect 27896 23264 27948 23316
rect 28356 23264 28408 23316
rect 27620 23239 27672 23248
rect 27620 23205 27629 23239
rect 27629 23205 27663 23239
rect 27663 23205 27672 23239
rect 27620 23196 27672 23205
rect 29552 23264 29604 23316
rect 30932 23307 30984 23316
rect 30932 23273 30941 23307
rect 30941 23273 30975 23307
rect 30975 23273 30984 23307
rect 30932 23264 30984 23273
rect 31484 23264 31536 23316
rect 32864 23264 32916 23316
rect 32956 23307 33008 23316
rect 32956 23273 32965 23307
rect 32965 23273 32999 23307
rect 32999 23273 33008 23307
rect 32956 23264 33008 23273
rect 35348 23264 35400 23316
rect 35532 23264 35584 23316
rect 36636 23264 36688 23316
rect 17224 23060 17276 23112
rect 17592 23060 17644 23112
rect 18420 23103 18472 23112
rect 18420 23069 18429 23103
rect 18429 23069 18463 23103
rect 18463 23069 18472 23103
rect 18420 23060 18472 23069
rect 12532 22967 12584 22976
rect 12532 22933 12541 22967
rect 12541 22933 12575 22967
rect 12575 22933 12584 22967
rect 12532 22924 12584 22933
rect 12716 22967 12768 22976
rect 12716 22933 12725 22967
rect 12725 22933 12759 22967
rect 12759 22933 12768 22967
rect 12716 22924 12768 22933
rect 12900 22924 12952 22976
rect 14280 22967 14332 22976
rect 14280 22933 14295 22967
rect 14295 22933 14329 22967
rect 14329 22933 14332 22967
rect 14280 22924 14332 22933
rect 14832 23035 14884 23044
rect 14832 23001 14866 23035
rect 14866 23001 14884 23035
rect 14832 22992 14884 23001
rect 22836 23060 22888 23112
rect 23112 23060 23164 23112
rect 24124 23103 24176 23112
rect 24124 23069 24133 23103
rect 24133 23069 24167 23103
rect 24167 23069 24176 23103
rect 24124 23060 24176 23069
rect 24676 23060 24728 23112
rect 26056 23103 26108 23112
rect 26056 23069 26065 23103
rect 26065 23069 26099 23103
rect 26099 23069 26108 23103
rect 26056 23060 26108 23069
rect 26700 23060 26752 23112
rect 15016 22924 15068 22976
rect 23020 22992 23072 23044
rect 25596 22992 25648 23044
rect 29092 23128 29144 23180
rect 32220 23171 32272 23180
rect 32220 23137 32229 23171
rect 32229 23137 32263 23171
rect 32263 23137 32272 23171
rect 32220 23128 32272 23137
rect 32404 23128 32456 23180
rect 36544 23196 36596 23248
rect 31208 23103 31260 23112
rect 31208 23069 31217 23103
rect 31217 23069 31251 23103
rect 31251 23069 31260 23103
rect 31208 23060 31260 23069
rect 32312 23060 32364 23112
rect 28080 22992 28132 23044
rect 28264 23035 28316 23044
rect 28264 23001 28273 23035
rect 28273 23001 28307 23035
rect 28307 23001 28316 23035
rect 28264 22992 28316 23001
rect 29368 22992 29420 23044
rect 33232 23060 33284 23112
rect 32864 22992 32916 23044
rect 36452 23128 36504 23180
rect 34152 23103 34204 23112
rect 15200 22924 15252 22976
rect 16120 22924 16172 22976
rect 17776 22967 17828 22976
rect 17776 22933 17785 22967
rect 17785 22933 17819 22967
rect 17819 22933 17828 22967
rect 17776 22924 17828 22933
rect 19340 22924 19392 22976
rect 23296 22967 23348 22976
rect 23296 22933 23305 22967
rect 23305 22933 23339 22967
rect 23339 22933 23348 22967
rect 23296 22924 23348 22933
rect 28356 22924 28408 22976
rect 29184 22924 29236 22976
rect 31024 22967 31076 22976
rect 31024 22933 31033 22967
rect 31033 22933 31067 22967
rect 31067 22933 31076 22967
rect 31024 22924 31076 22933
rect 32588 22967 32640 22976
rect 32588 22933 32623 22967
rect 32623 22933 32640 22967
rect 34152 23069 34161 23103
rect 34161 23069 34195 23103
rect 34195 23069 34204 23103
rect 34152 23060 34204 23069
rect 34428 23060 34480 23112
rect 34244 23035 34296 23044
rect 34244 23001 34253 23035
rect 34253 23001 34287 23035
rect 34287 23001 34296 23035
rect 34244 22992 34296 23001
rect 36084 23103 36136 23112
rect 36084 23069 36093 23103
rect 36093 23069 36127 23103
rect 36127 23069 36136 23103
rect 36084 23060 36136 23069
rect 36176 23060 36228 23112
rect 36728 23128 36780 23180
rect 36268 22992 36320 23044
rect 36636 23060 36688 23112
rect 37280 23103 37332 23112
rect 37280 23069 37314 23103
rect 37314 23069 37332 23103
rect 37280 23060 37332 23069
rect 35440 22967 35492 22976
rect 32588 22924 32640 22933
rect 35440 22933 35467 22967
rect 35467 22933 35492 22967
rect 35440 22924 35492 22933
rect 35532 22924 35584 22976
rect 38384 22967 38436 22976
rect 38384 22933 38393 22967
rect 38393 22933 38427 22967
rect 38427 22933 38436 22967
rect 38384 22924 38436 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 10048 22720 10100 22772
rect 10692 22720 10744 22772
rect 11336 22720 11388 22772
rect 11612 22720 11664 22772
rect 13176 22720 13228 22772
rect 13268 22763 13320 22772
rect 13268 22729 13277 22763
rect 13277 22729 13311 22763
rect 13311 22729 13320 22763
rect 13268 22720 13320 22729
rect 14280 22720 14332 22772
rect 14832 22720 14884 22772
rect 15016 22720 15068 22772
rect 17132 22720 17184 22772
rect 22744 22720 22796 22772
rect 23296 22720 23348 22772
rect 23388 22720 23440 22772
rect 8944 22652 8996 22704
rect 10324 22652 10376 22704
rect 7932 22627 7984 22636
rect 7932 22593 7941 22627
rect 7941 22593 7975 22627
rect 7975 22593 7984 22627
rect 7932 22584 7984 22593
rect 9864 22584 9916 22636
rect 9956 22627 10008 22636
rect 9956 22593 9965 22627
rect 9965 22593 9999 22627
rect 9999 22593 10008 22627
rect 9956 22584 10008 22593
rect 10600 22584 10652 22636
rect 10876 22627 10928 22636
rect 10876 22593 10885 22627
rect 10885 22593 10919 22627
rect 10919 22593 10928 22627
rect 10876 22584 10928 22593
rect 11152 22584 11204 22636
rect 12440 22584 12492 22636
rect 12900 22627 12952 22636
rect 12900 22593 12909 22627
rect 12909 22593 12943 22627
rect 12943 22593 12952 22627
rect 12900 22584 12952 22593
rect 11612 22559 11664 22568
rect 11612 22525 11621 22559
rect 11621 22525 11655 22559
rect 11655 22525 11664 22559
rect 11612 22516 11664 22525
rect 10140 22448 10192 22500
rect 12164 22516 12216 22568
rect 12900 22423 12952 22432
rect 12900 22389 12909 22423
rect 12909 22389 12943 22423
rect 12943 22389 12952 22423
rect 12900 22380 12952 22389
rect 14556 22584 14608 22636
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 16672 22652 16724 22704
rect 17592 22627 17644 22636
rect 17592 22593 17601 22627
rect 17601 22593 17635 22627
rect 17635 22593 17644 22627
rect 17592 22584 17644 22593
rect 19064 22652 19116 22704
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 19432 22627 19484 22636
rect 19432 22593 19441 22627
rect 19441 22593 19475 22627
rect 19475 22593 19484 22627
rect 19432 22584 19484 22593
rect 19708 22559 19760 22568
rect 19708 22525 19717 22559
rect 19717 22525 19751 22559
rect 19751 22525 19760 22559
rect 19708 22516 19760 22525
rect 20076 22584 20128 22636
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 20720 22584 20772 22593
rect 21088 22584 21140 22636
rect 21732 22584 21784 22636
rect 23020 22695 23072 22704
rect 23020 22661 23049 22695
rect 23049 22661 23072 22695
rect 23020 22652 23072 22661
rect 23204 22584 23256 22636
rect 23848 22720 23900 22772
rect 24124 22720 24176 22772
rect 24308 22763 24360 22772
rect 24308 22729 24317 22763
rect 24317 22729 24351 22763
rect 24351 22729 24360 22763
rect 24308 22720 24360 22729
rect 25136 22720 25188 22772
rect 24768 22652 24820 22704
rect 26056 22652 26108 22704
rect 28356 22720 28408 22772
rect 29368 22763 29420 22772
rect 29368 22729 29377 22763
rect 29377 22729 29411 22763
rect 29411 22729 29420 22763
rect 29368 22720 29420 22729
rect 24216 22584 24268 22636
rect 24676 22584 24728 22636
rect 20904 22516 20956 22568
rect 29092 22584 29144 22636
rect 16672 22423 16724 22432
rect 16672 22389 16681 22423
rect 16681 22389 16715 22423
rect 16715 22389 16724 22423
rect 16672 22380 16724 22389
rect 16948 22380 17000 22432
rect 23664 22491 23716 22500
rect 23664 22457 23673 22491
rect 23673 22457 23707 22491
rect 23707 22457 23716 22491
rect 23664 22448 23716 22457
rect 26332 22516 26384 22568
rect 28816 22559 28868 22568
rect 28816 22525 28825 22559
rect 28825 22525 28859 22559
rect 28859 22525 28868 22559
rect 28816 22516 28868 22525
rect 29276 22584 29328 22636
rect 30656 22720 30708 22772
rect 32220 22720 32272 22772
rect 26424 22448 26476 22500
rect 20720 22380 20772 22432
rect 21364 22423 21416 22432
rect 21364 22389 21373 22423
rect 21373 22389 21407 22423
rect 21407 22389 21416 22423
rect 21364 22380 21416 22389
rect 25504 22380 25556 22432
rect 30472 22584 30524 22636
rect 31024 22584 31076 22636
rect 30380 22559 30432 22568
rect 30380 22525 30389 22559
rect 30389 22525 30423 22559
rect 30423 22525 30432 22559
rect 30380 22516 30432 22525
rect 34244 22720 34296 22772
rect 36084 22720 36136 22772
rect 38384 22720 38436 22772
rect 33324 22584 33376 22636
rect 33876 22652 33928 22704
rect 34336 22652 34388 22704
rect 34520 22584 34572 22636
rect 32956 22516 33008 22568
rect 35624 22516 35676 22568
rect 38016 22652 38068 22704
rect 35348 22448 35400 22500
rect 32128 22423 32180 22432
rect 32128 22389 32137 22423
rect 32137 22389 32171 22423
rect 32171 22389 32180 22423
rect 32128 22380 32180 22389
rect 32404 22380 32456 22432
rect 32588 22380 32640 22432
rect 35256 22423 35308 22432
rect 35256 22389 35265 22423
rect 35265 22389 35299 22423
rect 35299 22389 35308 22423
rect 35256 22380 35308 22389
rect 35992 22380 36044 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 8944 22176 8996 22228
rect 9956 22176 10008 22228
rect 12164 22176 12216 22228
rect 12440 22108 12492 22160
rect 12900 22176 12952 22228
rect 15476 22219 15528 22228
rect 15476 22185 15485 22219
rect 15485 22185 15519 22219
rect 15519 22185 15528 22219
rect 15476 22176 15528 22185
rect 16948 22219 17000 22228
rect 16948 22185 16957 22219
rect 16957 22185 16991 22219
rect 16991 22185 17000 22219
rect 16948 22176 17000 22185
rect 19064 22176 19116 22228
rect 19248 22176 19300 22228
rect 19708 22176 19760 22228
rect 25504 22176 25556 22228
rect 26424 22219 26476 22228
rect 26424 22185 26433 22219
rect 26433 22185 26467 22219
rect 26467 22185 26476 22219
rect 26424 22176 26476 22185
rect 13084 22108 13136 22160
rect 18788 22108 18840 22160
rect 22836 22108 22888 22160
rect 8852 21972 8904 22024
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 10876 21972 10928 22024
rect 12532 21972 12584 22024
rect 11704 21904 11756 21956
rect 13360 22040 13412 22092
rect 15200 22040 15252 22092
rect 19248 22040 19300 22092
rect 13268 21972 13320 22024
rect 16580 22015 16632 22024
rect 16580 21981 16598 22015
rect 16598 21981 16632 22015
rect 16580 21972 16632 21981
rect 17592 22015 17644 22024
rect 17592 21981 17601 22015
rect 17601 21981 17635 22015
rect 17635 21981 17644 22015
rect 17592 21972 17644 21981
rect 10508 21836 10560 21888
rect 11152 21836 11204 21888
rect 11980 21836 12032 21888
rect 12440 21836 12492 21888
rect 13544 21836 13596 21888
rect 14004 21836 14056 21888
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 18052 21972 18104 22024
rect 17960 21836 18012 21888
rect 18420 22015 18472 22024
rect 18420 21981 18429 22015
rect 18429 21981 18463 22015
rect 18463 21981 18472 22015
rect 18420 21972 18472 21981
rect 23848 22040 23900 22092
rect 19156 21904 19208 21956
rect 20720 22015 20772 22024
rect 20720 21981 20729 22015
rect 20729 21981 20763 22015
rect 20763 21981 20772 22015
rect 20720 21972 20772 21981
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 24308 21972 24360 22024
rect 24400 22015 24452 22024
rect 24400 21981 24409 22015
rect 24409 21981 24443 22015
rect 24443 21981 24452 22015
rect 24400 21972 24452 21981
rect 26884 22108 26936 22160
rect 29368 22176 29420 22228
rect 31208 22176 31260 22228
rect 30380 22040 30432 22092
rect 20260 21904 20312 21956
rect 21272 21904 21324 21956
rect 22836 21904 22888 21956
rect 23388 21904 23440 21956
rect 24216 21947 24268 21956
rect 24216 21913 24225 21947
rect 24225 21913 24259 21947
rect 24259 21913 24268 21947
rect 24216 21904 24268 21913
rect 24676 21947 24728 21956
rect 24676 21913 24685 21947
rect 24685 21913 24719 21947
rect 24719 21913 24728 21947
rect 24676 21904 24728 21913
rect 18696 21836 18748 21888
rect 19064 21879 19116 21888
rect 19064 21845 19073 21879
rect 19073 21845 19107 21879
rect 19107 21845 19116 21879
rect 19064 21836 19116 21845
rect 22100 21836 22152 21888
rect 24492 21879 24544 21888
rect 24492 21845 24501 21879
rect 24501 21845 24535 21879
rect 24535 21845 24544 21879
rect 24492 21836 24544 21845
rect 25688 21879 25740 21888
rect 25688 21845 25697 21879
rect 25697 21845 25731 21879
rect 25731 21845 25740 21879
rect 25688 21836 25740 21845
rect 26700 21879 26752 21888
rect 26700 21845 26709 21879
rect 26709 21845 26743 21879
rect 26743 21845 26752 21879
rect 26700 21836 26752 21845
rect 27804 22015 27856 22024
rect 27804 21981 27813 22015
rect 27813 21981 27847 22015
rect 27847 21981 27856 22015
rect 27804 21972 27856 21981
rect 28172 21972 28224 22024
rect 32496 22176 32548 22228
rect 33232 22219 33284 22228
rect 33232 22185 33241 22219
rect 33241 22185 33275 22219
rect 33275 22185 33284 22219
rect 33232 22176 33284 22185
rect 33876 22108 33928 22160
rect 34520 22108 34572 22160
rect 34796 22108 34848 22160
rect 35532 22108 35584 22160
rect 36176 22176 36228 22228
rect 38016 22219 38068 22228
rect 36544 22108 36596 22160
rect 38016 22185 38025 22219
rect 38025 22185 38059 22219
rect 38059 22185 38068 22219
rect 38016 22176 38068 22185
rect 29460 21904 29512 21956
rect 27160 21836 27212 21888
rect 27988 21879 28040 21888
rect 27988 21845 27997 21879
rect 27997 21845 28031 21879
rect 28031 21845 28040 21879
rect 27988 21836 28040 21845
rect 28448 21836 28500 21888
rect 33324 22015 33376 22024
rect 33324 21981 33333 22015
rect 33333 21981 33367 22015
rect 33367 21981 33376 22015
rect 33324 21972 33376 21981
rect 34428 22040 34480 22092
rect 35164 22083 35216 22092
rect 35164 22049 35173 22083
rect 35173 22049 35207 22083
rect 35207 22049 35216 22083
rect 35164 22040 35216 22049
rect 35624 22083 35676 22092
rect 35624 22049 35633 22083
rect 35633 22049 35667 22083
rect 35667 22049 35676 22083
rect 35624 22040 35676 22049
rect 35900 22040 35952 22092
rect 36636 22083 36688 22092
rect 36636 22049 36645 22083
rect 36645 22049 36679 22083
rect 36679 22049 36688 22083
rect 36636 22040 36688 22049
rect 32128 21947 32180 21956
rect 32128 21913 32162 21947
rect 32162 21913 32180 21947
rect 32128 21904 32180 21913
rect 33048 21904 33100 21956
rect 31852 21836 31904 21888
rect 34796 21972 34848 22024
rect 35440 22009 35492 22024
rect 35440 21975 35446 22009
rect 35446 21975 35480 22009
rect 35480 21975 35492 22009
rect 35440 21972 35492 21975
rect 36728 21972 36780 22024
rect 35992 21947 36044 21956
rect 35992 21913 36019 21947
rect 36019 21913 36044 21947
rect 35992 21904 36044 21913
rect 35808 21879 35860 21888
rect 35808 21845 35817 21879
rect 35817 21845 35851 21879
rect 35851 21845 35860 21879
rect 35808 21836 35860 21845
rect 36268 21879 36320 21888
rect 36268 21845 36277 21879
rect 36277 21845 36311 21879
rect 36311 21845 36320 21879
rect 36268 21836 36320 21845
rect 36912 21947 36964 21956
rect 36912 21913 36946 21947
rect 36946 21913 36964 21947
rect 36912 21904 36964 21913
rect 36820 21836 36872 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 10324 21632 10376 21684
rect 10784 21632 10836 21684
rect 9864 21496 9916 21548
rect 10876 21496 10928 21548
rect 11152 21539 11204 21548
rect 11152 21505 11161 21539
rect 11161 21505 11195 21539
rect 11195 21505 11204 21539
rect 11152 21496 11204 21505
rect 11980 21632 12032 21684
rect 13912 21632 13964 21684
rect 14924 21632 14976 21684
rect 18420 21632 18472 21684
rect 19340 21632 19392 21684
rect 23112 21632 23164 21684
rect 26332 21632 26384 21684
rect 27988 21632 28040 21684
rect 28816 21632 28868 21684
rect 29460 21675 29512 21684
rect 29460 21641 29469 21675
rect 29469 21641 29503 21675
rect 29503 21641 29512 21675
rect 29460 21632 29512 21641
rect 11888 21607 11940 21616
rect 11888 21573 11897 21607
rect 11897 21573 11931 21607
rect 11931 21573 11940 21607
rect 11888 21564 11940 21573
rect 19156 21564 19208 21616
rect 11336 21428 11388 21480
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 12256 21496 12308 21548
rect 12716 21496 12768 21548
rect 13360 21539 13412 21548
rect 13360 21505 13369 21539
rect 13369 21505 13403 21539
rect 13403 21505 13412 21539
rect 13360 21496 13412 21505
rect 13912 21496 13964 21548
rect 14740 21496 14792 21548
rect 14096 21428 14148 21480
rect 17684 21539 17736 21548
rect 17684 21505 17693 21539
rect 17693 21505 17727 21539
rect 17727 21505 17736 21539
rect 17684 21496 17736 21505
rect 20904 21607 20956 21616
rect 20904 21573 20913 21607
rect 20913 21573 20947 21607
rect 20947 21573 20956 21607
rect 20904 21564 20956 21573
rect 26240 21564 26292 21616
rect 18052 21428 18104 21480
rect 10876 21360 10928 21412
rect 11888 21360 11940 21412
rect 16028 21360 16080 21412
rect 8484 21335 8536 21344
rect 8484 21301 8493 21335
rect 8493 21301 8527 21335
rect 8527 21301 8536 21335
rect 8484 21292 8536 21301
rect 11152 21292 11204 21344
rect 14280 21292 14332 21344
rect 17316 21335 17368 21344
rect 17316 21301 17325 21335
rect 17325 21301 17359 21335
rect 17359 21301 17368 21335
rect 17316 21292 17368 21301
rect 18236 21335 18288 21344
rect 18236 21301 18245 21335
rect 18245 21301 18279 21335
rect 18279 21301 18288 21335
rect 18236 21292 18288 21301
rect 19340 21292 19392 21344
rect 23940 21496 23992 21548
rect 24676 21496 24728 21548
rect 20720 21471 20772 21480
rect 20720 21437 20729 21471
rect 20729 21437 20763 21471
rect 20763 21437 20772 21471
rect 20720 21428 20772 21437
rect 22836 21428 22888 21480
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 24492 21428 24544 21480
rect 25228 21428 25280 21480
rect 25412 21496 25464 21548
rect 25596 21539 25648 21548
rect 25596 21505 25605 21539
rect 25605 21505 25639 21539
rect 25639 21505 25648 21539
rect 25596 21496 25648 21505
rect 25688 21496 25740 21548
rect 27712 21564 27764 21616
rect 26240 21428 26292 21480
rect 26424 21471 26476 21480
rect 26424 21437 26433 21471
rect 26433 21437 26467 21471
rect 26467 21437 26476 21471
rect 26424 21428 26476 21437
rect 29184 21496 29236 21548
rect 33876 21564 33928 21616
rect 35348 21632 35400 21684
rect 36268 21632 36320 21684
rect 35440 21607 35492 21616
rect 35440 21573 35449 21607
rect 35449 21573 35483 21607
rect 35483 21573 35492 21607
rect 35440 21564 35492 21573
rect 36728 21607 36780 21616
rect 36728 21573 36737 21607
rect 36737 21573 36771 21607
rect 36771 21573 36780 21607
rect 36728 21564 36780 21573
rect 29276 21471 29328 21480
rect 29276 21437 29285 21471
rect 29285 21437 29319 21471
rect 29319 21437 29328 21471
rect 29276 21428 29328 21437
rect 29368 21428 29420 21480
rect 34244 21496 34296 21548
rect 36636 21539 36688 21548
rect 36636 21505 36645 21539
rect 36645 21505 36679 21539
rect 36679 21505 36688 21539
rect 36636 21496 36688 21505
rect 32036 21428 32088 21480
rect 33048 21428 33100 21480
rect 23388 21360 23440 21412
rect 24216 21360 24268 21412
rect 25596 21360 25648 21412
rect 26608 21360 26660 21412
rect 36912 21403 36964 21412
rect 36912 21369 36921 21403
rect 36921 21369 36955 21403
rect 36955 21369 36964 21403
rect 36912 21360 36964 21369
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 20996 21335 21048 21344
rect 20996 21301 21005 21335
rect 21005 21301 21039 21335
rect 21039 21301 21048 21335
rect 20996 21292 21048 21301
rect 23480 21292 23532 21344
rect 25780 21335 25832 21344
rect 25780 21301 25789 21335
rect 25789 21301 25823 21335
rect 25823 21301 25832 21335
rect 25780 21292 25832 21301
rect 28724 21335 28776 21344
rect 28724 21301 28733 21335
rect 28733 21301 28767 21335
rect 28767 21301 28776 21335
rect 28724 21292 28776 21301
rect 30196 21292 30248 21344
rect 35348 21292 35400 21344
rect 35716 21292 35768 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 17960 21088 18012 21140
rect 20996 21088 21048 21140
rect 10324 20952 10376 21004
rect 10600 20952 10652 21004
rect 10968 20995 11020 21004
rect 10968 20961 10977 20995
rect 10977 20961 11011 20995
rect 11011 20961 11020 20995
rect 10968 20952 11020 20961
rect 9588 20884 9640 20936
rect 11060 20927 11112 20936
rect 11060 20893 11069 20927
rect 11069 20893 11103 20927
rect 11103 20893 11112 20927
rect 11060 20884 11112 20893
rect 11336 20927 11388 20936
rect 11336 20893 11345 20927
rect 11345 20893 11379 20927
rect 11379 20893 11388 20927
rect 11336 20884 11388 20893
rect 11888 20927 11940 20936
rect 11888 20893 11897 20927
rect 11897 20893 11931 20927
rect 11931 20893 11940 20927
rect 11888 20884 11940 20893
rect 14096 20995 14148 21004
rect 14096 20961 14105 20995
rect 14105 20961 14139 20995
rect 14139 20961 14148 20995
rect 14096 20952 14148 20961
rect 14280 20952 14332 21004
rect 12072 20927 12124 20936
rect 12072 20893 12081 20927
rect 12081 20893 12115 20927
rect 12115 20893 12124 20927
rect 12072 20884 12124 20893
rect 12256 20927 12308 20936
rect 12256 20893 12265 20927
rect 12265 20893 12299 20927
rect 12299 20893 12308 20927
rect 12256 20884 12308 20893
rect 8852 20816 8904 20868
rect 9404 20816 9456 20868
rect 8668 20791 8720 20800
rect 8668 20757 8677 20791
rect 8677 20757 8711 20791
rect 8711 20757 8720 20791
rect 8668 20748 8720 20757
rect 10784 20816 10836 20868
rect 11428 20859 11480 20868
rect 11428 20825 11437 20859
rect 11437 20825 11471 20859
rect 11471 20825 11480 20859
rect 11428 20816 11480 20825
rect 11796 20748 11848 20800
rect 13268 20884 13320 20936
rect 13360 20927 13412 20936
rect 13360 20893 13369 20927
rect 13369 20893 13403 20927
rect 13403 20893 13412 20927
rect 13360 20884 13412 20893
rect 17316 20927 17368 20936
rect 17316 20893 17334 20927
rect 17334 20893 17368 20927
rect 17316 20884 17368 20893
rect 12532 20859 12584 20868
rect 12532 20825 12541 20859
rect 12541 20825 12575 20859
rect 12575 20825 12584 20859
rect 12532 20816 12584 20825
rect 14832 20816 14884 20868
rect 19156 20884 19208 20936
rect 20260 20884 20312 20936
rect 21548 20884 21600 20936
rect 22928 20884 22980 20936
rect 18236 20816 18288 20868
rect 20076 20816 20128 20868
rect 22468 20816 22520 20868
rect 23112 20859 23164 20868
rect 23112 20825 23146 20859
rect 23146 20825 23164 20859
rect 23112 20816 23164 20825
rect 24216 21131 24268 21140
rect 24216 21097 24225 21131
rect 24225 21097 24259 21131
rect 24259 21097 24268 21131
rect 24216 21088 24268 21097
rect 25412 21088 25464 21140
rect 27804 21131 27856 21140
rect 27804 21097 27813 21131
rect 27813 21097 27847 21131
rect 27847 21097 27856 21131
rect 27804 21088 27856 21097
rect 28724 21088 28776 21140
rect 29276 21088 29328 21140
rect 29368 21131 29420 21140
rect 29368 21097 29377 21131
rect 29377 21097 29411 21131
rect 29411 21097 29420 21131
rect 29368 21088 29420 21097
rect 29552 21088 29604 21140
rect 30196 21131 30248 21140
rect 30196 21097 30205 21131
rect 30205 21097 30239 21131
rect 30239 21097 30248 21131
rect 30196 21088 30248 21097
rect 23940 20952 23992 21004
rect 29184 21020 29236 21072
rect 24676 20927 24728 20936
rect 24676 20893 24685 20927
rect 24685 20893 24719 20927
rect 24719 20893 24728 20927
rect 24676 20884 24728 20893
rect 25780 20884 25832 20936
rect 26240 20884 26292 20936
rect 26700 20927 26752 20936
rect 26700 20893 26734 20927
rect 26734 20893 26752 20927
rect 26700 20884 26752 20893
rect 28448 20816 28500 20868
rect 28816 20884 28868 20936
rect 15936 20748 15988 20800
rect 17316 20748 17368 20800
rect 17408 20748 17460 20800
rect 19340 20791 19392 20800
rect 19340 20757 19349 20791
rect 19349 20757 19383 20791
rect 19383 20757 19392 20791
rect 19340 20748 19392 20757
rect 20904 20791 20956 20800
rect 20904 20757 20913 20791
rect 20913 20757 20947 20791
rect 20947 20757 20956 20791
rect 20904 20748 20956 20757
rect 22376 20791 22428 20800
rect 22376 20757 22385 20791
rect 22385 20757 22419 20791
rect 22419 20757 22428 20791
rect 22376 20748 22428 20757
rect 24400 20791 24452 20800
rect 24400 20757 24409 20791
rect 24409 20757 24443 20791
rect 24443 20757 24452 20791
rect 24400 20748 24452 20757
rect 25228 20748 25280 20800
rect 27896 20791 27948 20800
rect 27896 20757 27905 20791
rect 27905 20757 27939 20791
rect 27939 20757 27948 20791
rect 27896 20748 27948 20757
rect 29276 20748 29328 20800
rect 34244 21131 34296 21140
rect 34244 21097 34253 21131
rect 34253 21097 34287 21131
rect 34287 21097 34296 21131
rect 34244 21088 34296 21097
rect 33140 21020 33192 21072
rect 33876 21020 33928 21072
rect 35900 21088 35952 21140
rect 32036 20884 32088 20936
rect 33876 20927 33928 20936
rect 33876 20893 33885 20927
rect 33885 20893 33919 20927
rect 33919 20893 33928 20927
rect 33876 20884 33928 20893
rect 35348 20952 35400 21004
rect 35440 20952 35492 21004
rect 32128 20816 32180 20868
rect 37188 20927 37240 20936
rect 37188 20893 37197 20927
rect 37197 20893 37231 20927
rect 37231 20893 37240 20927
rect 37188 20884 37240 20893
rect 30104 20748 30156 20800
rect 30472 20748 30524 20800
rect 30564 20791 30616 20800
rect 30564 20757 30573 20791
rect 30573 20757 30607 20791
rect 30607 20757 30616 20791
rect 30564 20748 30616 20757
rect 32864 20791 32916 20800
rect 32864 20757 32873 20791
rect 32873 20757 32907 20791
rect 32907 20757 32916 20791
rect 32864 20748 32916 20757
rect 35072 20748 35124 20800
rect 35348 20859 35400 20868
rect 35348 20825 35383 20859
rect 35383 20825 35400 20859
rect 35348 20816 35400 20825
rect 35532 20816 35584 20868
rect 35716 20816 35768 20868
rect 38660 20884 38712 20936
rect 37832 20791 37884 20800
rect 37832 20757 37841 20791
rect 37841 20757 37875 20791
rect 37875 20757 37884 20791
rect 37832 20748 37884 20757
rect 37924 20791 37976 20800
rect 37924 20757 37933 20791
rect 37933 20757 37967 20791
rect 37967 20757 37976 20791
rect 37924 20748 37976 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 11060 20544 11112 20596
rect 11428 20544 11480 20596
rect 11704 20587 11756 20596
rect 11704 20553 11713 20587
rect 11713 20553 11747 20587
rect 11747 20553 11756 20587
rect 11704 20544 11756 20553
rect 12072 20544 12124 20596
rect 14832 20544 14884 20596
rect 14924 20544 14976 20596
rect 8484 20476 8536 20528
rect 8668 20476 8720 20528
rect 11244 20519 11296 20528
rect 11244 20485 11253 20519
rect 11253 20485 11287 20519
rect 11287 20485 11296 20519
rect 11244 20476 11296 20485
rect 10324 20408 10376 20460
rect 7932 20383 7984 20392
rect 7932 20349 7941 20383
rect 7941 20349 7975 20383
rect 7975 20349 7984 20383
rect 7932 20340 7984 20349
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 11060 20272 11112 20324
rect 11704 20408 11756 20460
rect 12624 20476 12676 20528
rect 11888 20340 11940 20392
rect 13268 20408 13320 20460
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 13912 20451 13964 20460
rect 13912 20417 13921 20451
rect 13921 20417 13955 20451
rect 13955 20417 13964 20451
rect 13912 20408 13964 20417
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 16028 20451 16080 20460
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 17592 20544 17644 20596
rect 18052 20544 18104 20596
rect 20720 20544 20772 20596
rect 22376 20544 22428 20596
rect 23112 20544 23164 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 26424 20544 26476 20596
rect 27712 20587 27764 20596
rect 27712 20553 27721 20587
rect 27721 20553 27755 20587
rect 27755 20553 27764 20587
rect 27712 20544 27764 20553
rect 29184 20544 29236 20596
rect 17316 20476 17368 20528
rect 15292 20340 15344 20392
rect 12256 20204 12308 20256
rect 13268 20247 13320 20256
rect 13268 20213 13277 20247
rect 13277 20213 13311 20247
rect 13311 20213 13320 20247
rect 13268 20204 13320 20213
rect 14096 20247 14148 20256
rect 14096 20213 14105 20247
rect 14105 20213 14139 20247
rect 14139 20213 14148 20247
rect 14096 20204 14148 20213
rect 14648 20204 14700 20256
rect 15200 20247 15252 20256
rect 15200 20213 15209 20247
rect 15209 20213 15243 20247
rect 15243 20213 15252 20247
rect 15200 20204 15252 20213
rect 17960 20451 18012 20460
rect 17960 20417 17969 20451
rect 17969 20417 18003 20451
rect 18003 20417 18012 20451
rect 17960 20408 18012 20417
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 19340 20408 19392 20460
rect 20260 20451 20312 20460
rect 20260 20417 20269 20451
rect 20269 20417 20303 20451
rect 20303 20417 20312 20451
rect 20260 20408 20312 20417
rect 20904 20408 20956 20460
rect 22928 20476 22980 20528
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 23388 20451 23440 20460
rect 23388 20417 23397 20451
rect 23397 20417 23431 20451
rect 23431 20417 23440 20451
rect 23388 20408 23440 20417
rect 23480 20451 23532 20460
rect 23480 20417 23489 20451
rect 23489 20417 23523 20451
rect 23523 20417 23532 20451
rect 23480 20408 23532 20417
rect 24400 20408 24452 20460
rect 26240 20476 26292 20528
rect 28448 20519 28500 20528
rect 28448 20485 28457 20519
rect 28457 20485 28491 20519
rect 28491 20485 28500 20519
rect 28448 20476 28500 20485
rect 21180 20340 21232 20392
rect 21364 20315 21416 20324
rect 21364 20281 21373 20315
rect 21373 20281 21407 20315
rect 21407 20281 21416 20315
rect 21364 20272 21416 20281
rect 22376 20272 22428 20324
rect 24216 20340 24268 20392
rect 27896 20408 27948 20460
rect 29276 20408 29328 20460
rect 18512 20204 18564 20256
rect 22192 20204 22244 20256
rect 22836 20204 22888 20256
rect 28816 20340 28868 20392
rect 30104 20451 30156 20460
rect 30104 20417 30113 20451
rect 30113 20417 30147 20451
rect 30147 20417 30156 20451
rect 30104 20408 30156 20417
rect 30564 20408 30616 20460
rect 30472 20272 30524 20324
rect 31392 20451 31444 20460
rect 31392 20417 31401 20451
rect 31401 20417 31435 20451
rect 31435 20417 31444 20451
rect 31392 20408 31444 20417
rect 32128 20587 32180 20596
rect 32128 20553 32137 20587
rect 32137 20553 32171 20587
rect 32171 20553 32180 20587
rect 32128 20544 32180 20553
rect 35348 20544 35400 20596
rect 35440 20544 35492 20596
rect 37188 20544 37240 20596
rect 38660 20587 38712 20596
rect 38660 20553 38669 20587
rect 38669 20553 38703 20587
rect 38703 20553 38712 20587
rect 38660 20544 38712 20553
rect 33140 20476 33192 20528
rect 32864 20408 32916 20460
rect 34520 20408 34572 20460
rect 35072 20451 35124 20460
rect 35072 20417 35089 20451
rect 35089 20417 35123 20451
rect 35123 20417 35124 20451
rect 35624 20476 35676 20528
rect 35072 20408 35124 20417
rect 35348 20408 35400 20460
rect 35532 20451 35584 20460
rect 35532 20417 35541 20451
rect 35541 20417 35575 20451
rect 35575 20417 35584 20451
rect 35532 20408 35584 20417
rect 35808 20451 35860 20460
rect 35808 20417 35820 20451
rect 35820 20417 35854 20451
rect 35854 20417 35860 20451
rect 35808 20408 35860 20417
rect 36084 20451 36136 20460
rect 36084 20417 36093 20451
rect 36093 20417 36127 20451
rect 36127 20417 36136 20451
rect 36084 20408 36136 20417
rect 36176 20451 36228 20460
rect 36176 20417 36185 20451
rect 36185 20417 36219 20451
rect 36219 20417 36228 20451
rect 36176 20408 36228 20417
rect 23388 20204 23440 20256
rect 23756 20204 23808 20256
rect 24308 20204 24360 20256
rect 28540 20247 28592 20256
rect 28540 20213 28549 20247
rect 28549 20213 28583 20247
rect 28583 20213 28592 20247
rect 28540 20204 28592 20213
rect 29092 20204 29144 20256
rect 32680 20204 32732 20256
rect 36728 20408 36780 20460
rect 37832 20476 37884 20528
rect 37924 20408 37976 20460
rect 37280 20383 37332 20392
rect 37280 20349 37289 20383
rect 37289 20349 37323 20383
rect 37323 20349 37332 20383
rect 37280 20340 37332 20349
rect 32864 20204 32916 20256
rect 33692 20204 33744 20256
rect 35900 20204 35952 20256
rect 37188 20204 37240 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 9588 20043 9640 20052
rect 9588 20009 9597 20043
rect 9597 20009 9631 20043
rect 9631 20009 9640 20043
rect 9588 20000 9640 20009
rect 15200 20000 15252 20052
rect 16028 20000 16080 20052
rect 20076 20000 20128 20052
rect 21364 20000 21416 20052
rect 22468 20043 22520 20052
rect 22468 20009 22477 20043
rect 22477 20009 22511 20043
rect 22511 20009 22520 20043
rect 22468 20000 22520 20009
rect 22560 20043 22612 20052
rect 22560 20009 22569 20043
rect 22569 20009 22603 20043
rect 22603 20009 22612 20043
rect 22560 20000 22612 20009
rect 23020 20043 23072 20052
rect 23020 20009 23029 20043
rect 23029 20009 23063 20043
rect 23063 20009 23072 20043
rect 23020 20000 23072 20009
rect 23940 20000 23992 20052
rect 28540 20000 28592 20052
rect 29092 20043 29144 20052
rect 29092 20009 29101 20043
rect 29101 20009 29135 20043
rect 29135 20009 29144 20043
rect 29092 20000 29144 20009
rect 29368 20000 29420 20052
rect 30472 20000 30524 20052
rect 32772 20000 32824 20052
rect 10876 19864 10928 19916
rect 12532 19864 12584 19916
rect 22284 19932 22336 19984
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 12256 19796 12308 19848
rect 20260 19796 20312 19848
rect 20720 19839 20772 19848
rect 20720 19805 20729 19839
rect 20729 19805 20763 19839
rect 20763 19805 20772 19839
rect 20720 19796 20772 19805
rect 1768 19660 1820 19712
rect 11152 19728 11204 19780
rect 11612 19728 11664 19780
rect 12992 19771 13044 19780
rect 12992 19737 13001 19771
rect 13001 19737 13035 19771
rect 13035 19737 13044 19771
rect 12992 19728 13044 19737
rect 14096 19728 14148 19780
rect 15568 19728 15620 19780
rect 16304 19728 16356 19780
rect 16212 19660 16264 19712
rect 19984 19728 20036 19780
rect 21088 19796 21140 19848
rect 22192 19839 22244 19848
rect 22192 19805 22201 19839
rect 22201 19805 22235 19839
rect 22235 19805 22244 19839
rect 22192 19796 22244 19805
rect 22376 19796 22428 19848
rect 22468 19796 22520 19848
rect 24032 19932 24084 19984
rect 25228 19907 25280 19916
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 26240 19864 26292 19916
rect 27528 19907 27580 19916
rect 27528 19873 27537 19907
rect 27537 19873 27571 19907
rect 27571 19873 27580 19907
rect 27528 19864 27580 19873
rect 23296 19796 23348 19848
rect 23572 19839 23624 19848
rect 23572 19805 23581 19839
rect 23581 19805 23615 19839
rect 23615 19805 23624 19839
rect 23572 19796 23624 19805
rect 23756 19839 23808 19848
rect 23756 19805 23765 19839
rect 23765 19805 23799 19839
rect 23799 19805 23808 19839
rect 23756 19796 23808 19805
rect 23940 19796 23992 19848
rect 29736 19932 29788 19984
rect 29276 19839 29328 19848
rect 29276 19805 29285 19839
rect 29285 19805 29319 19839
rect 29319 19805 29328 19839
rect 29276 19796 29328 19805
rect 29368 19839 29420 19848
rect 29368 19805 29377 19839
rect 29377 19805 29411 19839
rect 29411 19805 29420 19839
rect 29368 19796 29420 19805
rect 35348 20000 35400 20052
rect 35440 20000 35492 20052
rect 36084 20000 36136 20052
rect 37188 20000 37240 20052
rect 35256 19864 35308 19916
rect 36176 19864 36228 19916
rect 37004 19864 37056 19916
rect 32036 19839 32088 19848
rect 32036 19805 32045 19839
rect 32045 19805 32079 19839
rect 32079 19805 32088 19839
rect 32036 19796 32088 19805
rect 22652 19728 22704 19780
rect 32864 19728 32916 19780
rect 32956 19728 33008 19780
rect 33692 19771 33744 19780
rect 20904 19660 20956 19712
rect 24584 19703 24636 19712
rect 24584 19669 24593 19703
rect 24593 19669 24627 19703
rect 24627 19669 24636 19703
rect 24584 19660 24636 19669
rect 30104 19660 30156 19712
rect 30564 19660 30616 19712
rect 32772 19660 32824 19712
rect 33692 19737 33701 19771
rect 33701 19737 33735 19771
rect 33735 19737 33744 19771
rect 33692 19728 33744 19737
rect 33416 19703 33468 19712
rect 33416 19669 33425 19703
rect 33425 19669 33459 19703
rect 33459 19669 33468 19703
rect 35900 19796 35952 19848
rect 34612 19728 34664 19780
rect 34888 19703 34940 19712
rect 33416 19660 33468 19669
rect 34888 19669 34897 19703
rect 34897 19669 34931 19703
rect 34931 19669 34940 19703
rect 34888 19660 34940 19669
rect 35164 19660 35216 19712
rect 35532 19703 35584 19712
rect 35532 19669 35559 19703
rect 35559 19669 35584 19703
rect 35532 19660 35584 19669
rect 35624 19660 35676 19712
rect 37004 19660 37056 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 11612 19456 11664 19508
rect 12992 19456 13044 19508
rect 14648 19388 14700 19440
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 14280 19320 14332 19372
rect 16212 19456 16264 19508
rect 16304 19456 16356 19508
rect 18512 19499 18564 19508
rect 18512 19465 18521 19499
rect 18521 19465 18555 19499
rect 18555 19465 18564 19499
rect 18512 19456 18564 19465
rect 20996 19456 21048 19508
rect 16304 19363 16356 19372
rect 16304 19329 16313 19363
rect 16313 19329 16347 19363
rect 16347 19329 16356 19363
rect 16304 19320 16356 19329
rect 17316 19363 17368 19372
rect 17316 19329 17350 19363
rect 17350 19329 17368 19363
rect 17316 19320 17368 19329
rect 19800 19320 19852 19372
rect 21548 19388 21600 19440
rect 29736 19456 29788 19508
rect 30656 19456 30708 19508
rect 31852 19456 31904 19508
rect 32772 19499 32824 19508
rect 32772 19465 32781 19499
rect 32781 19465 32815 19499
rect 32815 19465 32824 19499
rect 32772 19456 32824 19465
rect 32956 19456 33008 19508
rect 19984 19320 20036 19372
rect 11060 19252 11112 19304
rect 14096 19252 14148 19304
rect 14464 19116 14516 19168
rect 20628 19320 20680 19372
rect 20904 19320 20956 19372
rect 21180 19363 21232 19372
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 21272 19320 21324 19372
rect 21640 19363 21692 19372
rect 21640 19329 21649 19363
rect 21649 19329 21683 19363
rect 21683 19329 21692 19363
rect 21640 19320 21692 19329
rect 22284 19388 22336 19440
rect 22928 19320 22980 19372
rect 23296 19320 23348 19372
rect 24584 19320 24636 19372
rect 26516 19388 26568 19440
rect 28080 19388 28132 19440
rect 25688 19363 25740 19372
rect 25688 19329 25722 19363
rect 25722 19329 25740 19363
rect 25688 19320 25740 19329
rect 29920 19363 29972 19372
rect 29920 19329 29929 19363
rect 29929 19329 29963 19363
rect 29963 19329 29972 19363
rect 29920 19320 29972 19329
rect 30288 19320 30340 19372
rect 30104 19295 30156 19304
rect 30104 19261 30113 19295
rect 30113 19261 30147 19295
rect 30147 19261 30156 19295
rect 30104 19252 30156 19261
rect 20720 19184 20772 19236
rect 21180 19184 21232 19236
rect 27252 19184 27304 19236
rect 31392 19388 31444 19440
rect 31668 19431 31720 19440
rect 31668 19397 31697 19431
rect 31697 19397 31720 19431
rect 31668 19388 31720 19397
rect 17408 19116 17460 19168
rect 18420 19159 18472 19168
rect 18420 19125 18429 19159
rect 18429 19125 18463 19159
rect 18463 19125 18472 19159
rect 18420 19116 18472 19125
rect 20904 19116 20956 19168
rect 21272 19116 21324 19168
rect 23480 19116 23532 19168
rect 23940 19159 23992 19168
rect 23940 19125 23949 19159
rect 23949 19125 23983 19159
rect 23983 19125 23992 19159
rect 23940 19116 23992 19125
rect 26056 19116 26108 19168
rect 26884 19116 26936 19168
rect 27712 19159 27764 19168
rect 27712 19125 27721 19159
rect 27721 19125 27755 19159
rect 27755 19125 27764 19159
rect 27712 19116 27764 19125
rect 33416 19388 33468 19440
rect 34520 19388 34572 19440
rect 35072 19388 35124 19440
rect 31944 19363 31996 19372
rect 31944 19329 31953 19363
rect 31953 19329 31987 19363
rect 31987 19329 31996 19363
rect 31944 19320 31996 19329
rect 32680 19320 32732 19372
rect 33140 19320 33192 19372
rect 35256 19431 35308 19440
rect 35256 19397 35265 19431
rect 35265 19397 35299 19431
rect 35299 19397 35308 19431
rect 35256 19388 35308 19397
rect 37004 19499 37056 19508
rect 37004 19465 37013 19499
rect 37013 19465 37047 19499
rect 37047 19465 37056 19499
rect 37004 19456 37056 19465
rect 35532 19363 35584 19372
rect 35532 19329 35541 19363
rect 35541 19329 35575 19363
rect 35575 19329 35584 19363
rect 35532 19320 35584 19329
rect 34612 19295 34664 19304
rect 34612 19261 34621 19295
rect 34621 19261 34655 19295
rect 34655 19261 34664 19295
rect 34612 19252 34664 19261
rect 35072 19252 35124 19304
rect 37280 19320 37332 19372
rect 30748 19116 30800 19168
rect 32680 19116 32732 19168
rect 34796 19159 34848 19168
rect 34796 19125 34805 19159
rect 34805 19125 34839 19159
rect 34839 19125 34848 19159
rect 34796 19116 34848 19125
rect 34888 19116 34940 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 12624 18776 12676 18828
rect 9496 18708 9548 18760
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 11060 18751 11112 18760
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 14280 18912 14332 18964
rect 14096 18844 14148 18896
rect 18604 18912 18656 18964
rect 19800 18912 19852 18964
rect 21916 18912 21968 18964
rect 23572 18912 23624 18964
rect 23664 18912 23716 18964
rect 15568 18819 15620 18828
rect 15568 18785 15577 18819
rect 15577 18785 15611 18819
rect 15611 18785 15620 18819
rect 15568 18776 15620 18785
rect 13452 18640 13504 18692
rect 9496 18615 9548 18624
rect 9496 18581 9505 18615
rect 9505 18581 9539 18615
rect 9539 18581 9548 18615
rect 9496 18572 9548 18581
rect 10140 18572 10192 18624
rect 10968 18615 11020 18624
rect 10968 18581 10977 18615
rect 10977 18581 11011 18615
rect 11011 18581 11020 18615
rect 10968 18572 11020 18581
rect 12164 18615 12216 18624
rect 12164 18581 12173 18615
rect 12173 18581 12207 18615
rect 12207 18581 12216 18615
rect 12164 18572 12216 18581
rect 13084 18572 13136 18624
rect 13176 18615 13228 18624
rect 13176 18581 13185 18615
rect 13185 18581 13219 18615
rect 13219 18581 13228 18615
rect 13176 18572 13228 18581
rect 13728 18572 13780 18624
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 18420 18776 18472 18828
rect 20444 18776 20496 18828
rect 17408 18751 17460 18760
rect 17408 18717 17417 18751
rect 17417 18717 17451 18751
rect 17451 18717 17460 18751
rect 17408 18708 17460 18717
rect 17868 18708 17920 18760
rect 18052 18751 18104 18760
rect 18052 18717 18061 18751
rect 18061 18717 18095 18751
rect 18095 18717 18104 18751
rect 18052 18708 18104 18717
rect 18512 18708 18564 18760
rect 20260 18751 20312 18760
rect 20260 18717 20269 18751
rect 20269 18717 20303 18751
rect 20303 18717 20312 18751
rect 20260 18708 20312 18717
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 17960 18572 18012 18624
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 19340 18572 19392 18624
rect 20168 18572 20220 18624
rect 20444 18683 20496 18692
rect 20444 18649 20479 18683
rect 20479 18649 20496 18683
rect 20444 18640 20496 18649
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 22100 18819 22152 18828
rect 22100 18785 22109 18819
rect 22109 18785 22143 18819
rect 22143 18785 22152 18819
rect 22100 18776 22152 18785
rect 22284 18819 22336 18828
rect 22284 18785 22293 18819
rect 22293 18785 22327 18819
rect 22327 18785 22336 18819
rect 22284 18776 22336 18785
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 22836 18708 22888 18760
rect 22652 18640 22704 18692
rect 22100 18572 22152 18624
rect 23204 18751 23256 18760
rect 23204 18717 23213 18751
rect 23213 18717 23247 18751
rect 23247 18717 23256 18751
rect 23204 18708 23256 18717
rect 23388 18751 23440 18760
rect 23388 18717 23397 18751
rect 23397 18717 23431 18751
rect 23431 18717 23440 18751
rect 23388 18708 23440 18717
rect 25044 18776 25096 18828
rect 25596 18912 25648 18964
rect 25688 18912 25740 18964
rect 29920 18912 29972 18964
rect 28724 18887 28776 18896
rect 28724 18853 28733 18887
rect 28733 18853 28767 18887
rect 28767 18853 28776 18887
rect 28724 18844 28776 18853
rect 27712 18776 27764 18828
rect 28816 18776 28868 18828
rect 25596 18708 25648 18760
rect 26608 18751 26660 18760
rect 26608 18717 26617 18751
rect 26617 18717 26651 18751
rect 26651 18717 26660 18751
rect 26608 18708 26660 18717
rect 25872 18640 25924 18692
rect 28080 18708 28132 18760
rect 27068 18572 27120 18624
rect 29184 18708 29236 18760
rect 31392 18912 31444 18964
rect 29644 18640 29696 18692
rect 30564 18844 30616 18896
rect 30840 18844 30892 18896
rect 31760 18912 31812 18964
rect 33968 18912 34020 18964
rect 34612 18912 34664 18964
rect 34980 18887 35032 18896
rect 34980 18853 34989 18887
rect 34989 18853 35023 18887
rect 35023 18853 35032 18887
rect 34980 18844 35032 18853
rect 36728 18844 36780 18896
rect 30748 18819 30800 18828
rect 30748 18785 30757 18819
rect 30757 18785 30791 18819
rect 30791 18785 30800 18819
rect 30748 18776 30800 18785
rect 31668 18776 31720 18828
rect 32588 18819 32640 18828
rect 32588 18785 32597 18819
rect 32597 18785 32631 18819
rect 32631 18785 32640 18819
rect 32588 18776 32640 18785
rect 32956 18819 33008 18828
rect 32956 18785 32965 18819
rect 32965 18785 32999 18819
rect 32999 18785 33008 18819
rect 32956 18776 33008 18785
rect 32680 18708 32732 18760
rect 29736 18572 29788 18624
rect 30288 18683 30340 18692
rect 30288 18649 30297 18683
rect 30297 18649 30331 18683
rect 30331 18649 30340 18683
rect 30288 18640 30340 18649
rect 34796 18751 34848 18760
rect 34796 18717 34805 18751
rect 34805 18717 34839 18751
rect 34839 18717 34848 18751
rect 34796 18708 34848 18717
rect 37188 18751 37240 18760
rect 37188 18717 37197 18751
rect 37197 18717 37231 18751
rect 37231 18717 37240 18751
rect 37188 18708 37240 18717
rect 38292 18640 38344 18692
rect 36636 18572 36688 18624
rect 37004 18615 37056 18624
rect 37004 18581 37013 18615
rect 37013 18581 37047 18615
rect 37047 18581 37056 18615
rect 37004 18572 37056 18581
rect 38476 18572 38528 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 7932 18368 7984 18420
rect 9496 18300 9548 18352
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 10876 18368 10928 18420
rect 11520 18368 11572 18420
rect 12164 18368 12216 18420
rect 13176 18368 13228 18420
rect 10140 18300 10192 18352
rect 10968 18232 11020 18284
rect 8484 18164 8536 18216
rect 13360 18300 13412 18352
rect 13728 18368 13780 18420
rect 14464 18300 14516 18352
rect 15476 18368 15528 18420
rect 12532 18232 12584 18284
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 15568 18096 15620 18148
rect 17316 18368 17368 18420
rect 18052 18368 18104 18420
rect 18328 18368 18380 18420
rect 17500 18232 17552 18284
rect 17776 18275 17828 18284
rect 17776 18241 17785 18275
rect 17785 18241 17819 18275
rect 17819 18241 17828 18275
rect 17776 18232 17828 18241
rect 17224 18207 17276 18216
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 17960 18275 18012 18284
rect 17960 18241 17995 18275
rect 17995 18241 18012 18275
rect 17960 18232 18012 18241
rect 18604 18368 18656 18420
rect 19432 18368 19484 18420
rect 19340 18300 19392 18352
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 20444 18368 20496 18420
rect 22652 18411 22704 18420
rect 22652 18377 22661 18411
rect 22661 18377 22695 18411
rect 22695 18377 22704 18411
rect 22652 18368 22704 18377
rect 23204 18368 23256 18420
rect 20720 18300 20772 18352
rect 20812 18300 20864 18352
rect 28724 18368 28776 18420
rect 29184 18411 29236 18420
rect 29184 18377 29193 18411
rect 29193 18377 29227 18411
rect 29227 18377 29236 18411
rect 29184 18368 29236 18377
rect 30288 18368 30340 18420
rect 36728 18368 36780 18420
rect 37004 18368 37056 18420
rect 25044 18343 25096 18352
rect 25044 18309 25053 18343
rect 25053 18309 25087 18343
rect 25087 18309 25096 18343
rect 25044 18300 25096 18309
rect 34980 18300 35032 18352
rect 18972 18207 19024 18216
rect 18972 18173 18981 18207
rect 18981 18173 19015 18207
rect 19015 18173 19024 18207
rect 18972 18164 19024 18173
rect 19340 18164 19392 18216
rect 20076 18164 20128 18216
rect 9864 18028 9916 18080
rect 11612 18071 11664 18080
rect 11612 18037 11621 18071
rect 11621 18037 11655 18071
rect 11655 18037 11664 18071
rect 11612 18028 11664 18037
rect 11796 18028 11848 18080
rect 13452 18028 13504 18080
rect 15476 18028 15528 18080
rect 16764 18028 16816 18080
rect 19432 18096 19484 18148
rect 18144 18028 18196 18080
rect 21916 18275 21968 18284
rect 21916 18241 21925 18275
rect 21925 18241 21959 18275
rect 21959 18241 21968 18275
rect 21916 18232 21968 18241
rect 20996 18164 21048 18216
rect 21824 18164 21876 18216
rect 22928 18232 22980 18284
rect 24400 18232 24452 18284
rect 25504 18275 25556 18284
rect 25504 18241 25513 18275
rect 25513 18241 25547 18275
rect 25547 18241 25556 18275
rect 25504 18232 25556 18241
rect 25688 18232 25740 18284
rect 25964 18232 26016 18284
rect 27528 18232 27580 18284
rect 31944 18232 31996 18284
rect 20904 18096 20956 18148
rect 26608 18164 26660 18216
rect 27620 18207 27672 18216
rect 27620 18173 27629 18207
rect 27629 18173 27663 18207
rect 27663 18173 27672 18207
rect 27620 18164 27672 18173
rect 31208 18164 31260 18216
rect 35348 18275 35400 18284
rect 35348 18241 35357 18275
rect 35357 18241 35391 18275
rect 35391 18241 35400 18275
rect 35348 18232 35400 18241
rect 36636 18343 36688 18352
rect 36636 18309 36645 18343
rect 36645 18309 36679 18343
rect 36679 18309 36688 18343
rect 36636 18300 36688 18309
rect 36084 18232 36136 18284
rect 36360 18275 36412 18284
rect 36360 18241 36369 18275
rect 36369 18241 36403 18275
rect 36403 18241 36412 18275
rect 36360 18232 36412 18241
rect 36452 18275 36504 18284
rect 36452 18241 36462 18275
rect 36462 18241 36496 18275
rect 36496 18241 36504 18275
rect 36452 18232 36504 18241
rect 25872 18096 25924 18148
rect 23296 18028 23348 18080
rect 25412 18028 25464 18080
rect 25596 18028 25648 18080
rect 31024 18028 31076 18080
rect 34796 18028 34848 18080
rect 36728 18275 36780 18284
rect 36728 18241 36737 18275
rect 36737 18241 36771 18275
rect 36771 18241 36780 18275
rect 36728 18232 36780 18241
rect 36912 18232 36964 18284
rect 37188 18232 37240 18284
rect 37280 18275 37332 18284
rect 37280 18241 37289 18275
rect 37289 18241 37323 18275
rect 37323 18241 37332 18275
rect 37280 18232 37332 18241
rect 38476 18028 38528 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 8484 17824 8536 17876
rect 10600 17824 10652 17876
rect 10876 17824 10928 17876
rect 13084 17824 13136 17876
rect 20720 17867 20772 17876
rect 20720 17833 20729 17867
rect 20729 17833 20763 17867
rect 20763 17833 20772 17867
rect 20720 17824 20772 17833
rect 20352 17756 20404 17808
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 11520 17688 11572 17740
rect 11612 17688 11664 17740
rect 13176 17688 13228 17740
rect 13728 17688 13780 17740
rect 15108 17731 15160 17740
rect 15108 17697 15117 17731
rect 15117 17697 15151 17731
rect 15151 17697 15160 17731
rect 15108 17688 15160 17697
rect 19340 17688 19392 17740
rect 22284 17824 22336 17876
rect 24400 17824 24452 17876
rect 21640 17688 21692 17740
rect 21824 17731 21876 17740
rect 21824 17697 21833 17731
rect 21833 17697 21867 17731
rect 21867 17697 21876 17731
rect 21824 17688 21876 17697
rect 17868 17620 17920 17672
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 23020 17688 23072 17740
rect 23296 17688 23348 17740
rect 12716 17552 12768 17604
rect 15384 17595 15436 17604
rect 15384 17561 15418 17595
rect 15418 17561 15436 17595
rect 15384 17552 15436 17561
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 11796 17484 11848 17536
rect 15568 17484 15620 17536
rect 16580 17527 16632 17536
rect 16580 17493 16589 17527
rect 16589 17493 16623 17527
rect 16623 17493 16632 17527
rect 16580 17484 16632 17493
rect 19340 17595 19392 17604
rect 19340 17561 19349 17595
rect 19349 17561 19383 17595
rect 19383 17561 19392 17595
rect 19340 17552 19392 17561
rect 19524 17552 19576 17604
rect 20628 17552 20680 17604
rect 23940 17688 23992 17740
rect 22376 17552 22428 17604
rect 23204 17552 23256 17604
rect 23756 17620 23808 17672
rect 23848 17552 23900 17604
rect 25136 17663 25188 17672
rect 25136 17629 25145 17663
rect 25145 17629 25179 17663
rect 25179 17629 25188 17663
rect 25136 17620 25188 17629
rect 25412 17663 25464 17672
rect 25412 17629 25446 17663
rect 25446 17629 25464 17663
rect 27620 17824 27672 17876
rect 31208 17824 31260 17876
rect 30288 17688 30340 17740
rect 30656 17688 30708 17740
rect 27988 17663 28040 17672
rect 25412 17620 25464 17629
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 28264 17663 28316 17672
rect 28264 17629 28273 17663
rect 28273 17629 28307 17663
rect 28307 17629 28316 17663
rect 28264 17620 28316 17629
rect 30748 17663 30800 17672
rect 30748 17629 30757 17663
rect 30757 17629 30791 17663
rect 30791 17629 30800 17663
rect 30748 17620 30800 17629
rect 30840 17663 30892 17672
rect 30840 17629 30849 17663
rect 30849 17629 30883 17663
rect 30883 17629 30892 17663
rect 30840 17620 30892 17629
rect 31024 17620 31076 17672
rect 31484 17663 31536 17672
rect 31484 17629 31493 17663
rect 31493 17629 31527 17663
rect 31527 17629 31536 17663
rect 31484 17620 31536 17629
rect 35348 17824 35400 17876
rect 33968 17756 34020 17808
rect 34520 17620 34572 17672
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 21088 17527 21140 17536
rect 21088 17493 21097 17527
rect 21097 17493 21131 17527
rect 21131 17493 21140 17527
rect 21088 17484 21140 17493
rect 22100 17484 22152 17536
rect 22192 17527 22244 17536
rect 22192 17493 22201 17527
rect 22201 17493 22235 17527
rect 22235 17493 22244 17527
rect 22192 17484 22244 17493
rect 22284 17527 22336 17536
rect 22284 17493 22293 17527
rect 22293 17493 22327 17527
rect 22327 17493 22336 17527
rect 22284 17484 22336 17493
rect 26516 17484 26568 17536
rect 29828 17527 29880 17536
rect 29828 17493 29837 17527
rect 29837 17493 29871 17527
rect 29871 17493 29880 17527
rect 29828 17484 29880 17493
rect 35900 17824 35952 17876
rect 36084 17799 36136 17808
rect 36084 17765 36093 17799
rect 36093 17765 36127 17799
rect 36127 17765 36136 17799
rect 36084 17756 36136 17765
rect 38292 17867 38344 17876
rect 38292 17833 38301 17867
rect 38301 17833 38335 17867
rect 38335 17833 38344 17867
rect 38292 17824 38344 17833
rect 36452 17620 36504 17672
rect 36820 17663 36872 17672
rect 36820 17629 36829 17663
rect 36829 17629 36863 17663
rect 36863 17629 36872 17663
rect 36820 17620 36872 17629
rect 36912 17620 36964 17672
rect 36728 17552 36780 17604
rect 33784 17484 33836 17536
rect 34704 17484 34756 17536
rect 37188 17663 37240 17672
rect 37188 17629 37197 17663
rect 37197 17629 37231 17663
rect 37231 17629 37240 17663
rect 37188 17620 37240 17629
rect 37832 17663 37884 17672
rect 37832 17629 37841 17663
rect 37841 17629 37875 17663
rect 37875 17629 37884 17663
rect 37832 17620 37884 17629
rect 37924 17595 37976 17604
rect 37924 17561 37933 17595
rect 37933 17561 37967 17595
rect 37967 17561 37976 17595
rect 37924 17552 37976 17561
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4068 17280 4120 17332
rect 7748 17212 7800 17264
rect 8484 17212 8536 17264
rect 9128 17212 9180 17264
rect 9956 17212 10008 17264
rect 10876 17212 10928 17264
rect 12716 17280 12768 17332
rect 15384 17280 15436 17332
rect 17224 17280 17276 17332
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 19064 17323 19116 17332
rect 19064 17289 19073 17323
rect 19073 17289 19107 17323
rect 19107 17289 19116 17323
rect 19064 17280 19116 17289
rect 18880 17212 18932 17264
rect 19156 17212 19208 17264
rect 24676 17280 24728 17332
rect 25504 17280 25556 17332
rect 8760 17076 8812 17128
rect 9680 17144 9732 17196
rect 13820 17144 13872 17196
rect 15016 17144 15068 17196
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 9864 17076 9916 17128
rect 10692 17076 10744 17128
rect 9312 16940 9364 16992
rect 10140 16940 10192 16992
rect 14924 16940 14976 16992
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15476 17144 15528 17153
rect 15568 17187 15620 17196
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 15660 17076 15712 17128
rect 16028 17076 16080 17128
rect 16580 17144 16632 17196
rect 18144 17144 18196 17196
rect 18972 17144 19024 17196
rect 16764 17076 16816 17128
rect 17592 17119 17644 17128
rect 17592 17085 17601 17119
rect 17601 17085 17635 17119
rect 17635 17085 17644 17119
rect 17592 17076 17644 17085
rect 15844 16983 15896 16992
rect 15844 16949 15853 16983
rect 15853 16949 15887 16983
rect 15887 16949 15896 16983
rect 15844 16940 15896 16949
rect 16396 16940 16448 16992
rect 19064 17076 19116 17128
rect 21640 17144 21692 17196
rect 22284 17144 22336 17196
rect 23112 17255 23164 17264
rect 23112 17221 23121 17255
rect 23121 17221 23155 17255
rect 23155 17221 23164 17255
rect 23112 17212 23164 17221
rect 26332 17280 26384 17332
rect 25964 17212 26016 17264
rect 26700 17280 26752 17332
rect 28264 17280 28316 17332
rect 29736 17323 29788 17332
rect 29736 17289 29745 17323
rect 29745 17289 29779 17323
rect 29779 17289 29788 17323
rect 29736 17280 29788 17289
rect 29828 17280 29880 17332
rect 20444 17076 20496 17128
rect 21272 17119 21324 17128
rect 21272 17085 21281 17119
rect 21281 17085 21315 17119
rect 21315 17085 21324 17119
rect 21272 17076 21324 17085
rect 23204 17076 23256 17128
rect 26608 17187 26660 17196
rect 26608 17153 26617 17187
rect 26617 17153 26651 17187
rect 26651 17153 26660 17187
rect 26608 17144 26660 17153
rect 26700 17144 26752 17196
rect 29644 17187 29696 17196
rect 29644 17153 29653 17187
rect 29653 17153 29687 17187
rect 29687 17153 29696 17187
rect 29644 17144 29696 17153
rect 34612 17280 34664 17332
rect 34704 17323 34756 17332
rect 34704 17289 34713 17323
rect 34713 17289 34747 17323
rect 34747 17289 34756 17323
rect 34704 17280 34756 17289
rect 34796 17280 34848 17332
rect 36820 17280 36872 17332
rect 37832 17280 37884 17332
rect 33784 17212 33836 17264
rect 33968 17212 34020 17264
rect 31852 17144 31904 17196
rect 27712 17076 27764 17128
rect 27896 17119 27948 17128
rect 27896 17085 27905 17119
rect 27905 17085 27939 17119
rect 27939 17085 27948 17119
rect 27896 17076 27948 17085
rect 30748 17076 30800 17128
rect 19524 17008 19576 17060
rect 22652 17008 22704 17060
rect 25228 17051 25280 17060
rect 25228 17017 25237 17051
rect 25237 17017 25271 17051
rect 25271 17017 25280 17051
rect 25228 17008 25280 17017
rect 25688 17008 25740 17060
rect 19432 16940 19484 16992
rect 20812 16940 20864 16992
rect 22376 16940 22428 16992
rect 23112 16940 23164 16992
rect 25872 16940 25924 16992
rect 27620 16983 27672 16992
rect 27620 16949 27629 16983
rect 27629 16949 27663 16983
rect 27663 16949 27672 16983
rect 27620 16940 27672 16949
rect 28264 16940 28316 16992
rect 33416 16940 33468 16992
rect 34520 17076 34572 17128
rect 37096 17212 37148 17264
rect 38292 17280 38344 17332
rect 36820 17119 36872 17128
rect 36820 17085 36829 17119
rect 36829 17085 36863 17119
rect 36863 17085 36872 17119
rect 36820 17076 36872 17085
rect 37188 17076 37240 17128
rect 37924 17119 37976 17128
rect 37924 17085 37933 17119
rect 37933 17085 37967 17119
rect 37967 17085 37976 17119
rect 37924 17076 37976 17085
rect 38108 16983 38160 16992
rect 38108 16949 38117 16983
rect 38117 16949 38151 16983
rect 38151 16949 38160 16983
rect 38108 16940 38160 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 8484 16736 8536 16788
rect 8760 16736 8812 16788
rect 13728 16736 13780 16788
rect 8668 16600 8720 16652
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 10048 16668 10100 16720
rect 11428 16668 11480 16720
rect 11520 16600 11572 16652
rect 9496 16507 9548 16516
rect 9496 16473 9505 16507
rect 9505 16473 9539 16507
rect 9539 16473 9548 16507
rect 9496 16464 9548 16473
rect 9864 16507 9916 16516
rect 9864 16473 9873 16507
rect 9873 16473 9907 16507
rect 9907 16473 9916 16507
rect 9864 16464 9916 16473
rect 9956 16507 10008 16516
rect 9956 16473 9965 16507
rect 9965 16473 9999 16507
rect 9999 16473 10008 16507
rect 9956 16464 10008 16473
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 12624 16600 12676 16652
rect 15016 16736 15068 16788
rect 18144 16736 18196 16788
rect 18972 16736 19024 16788
rect 11888 16575 11940 16584
rect 11888 16541 11890 16575
rect 11890 16541 11924 16575
rect 11924 16541 11940 16575
rect 10416 16507 10468 16516
rect 10416 16473 10425 16507
rect 10425 16473 10459 16507
rect 10459 16473 10468 16507
rect 10416 16464 10468 16473
rect 11060 16464 11112 16516
rect 11888 16532 11940 16541
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 14740 16575 14792 16584
rect 14740 16541 14749 16575
rect 14749 16541 14783 16575
rect 14783 16541 14792 16575
rect 14740 16532 14792 16541
rect 16396 16668 16448 16720
rect 15568 16600 15620 16652
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 19432 16668 19484 16720
rect 19524 16668 19576 16720
rect 19984 16736 20036 16788
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 12440 16396 12492 16405
rect 13084 16396 13136 16448
rect 14188 16439 14240 16448
rect 14188 16405 14197 16439
rect 14197 16405 14231 16439
rect 14231 16405 14240 16439
rect 14188 16396 14240 16405
rect 19340 16532 19392 16584
rect 27896 16736 27948 16788
rect 25044 16600 25096 16652
rect 25228 16668 25280 16720
rect 25412 16600 25464 16652
rect 22100 16532 22152 16584
rect 23112 16575 23164 16584
rect 23112 16541 23146 16575
rect 23146 16541 23164 16575
rect 23112 16532 23164 16541
rect 27988 16643 28040 16652
rect 27988 16609 27997 16643
rect 27997 16609 28031 16643
rect 28031 16609 28040 16643
rect 27988 16600 28040 16609
rect 30656 16736 30708 16788
rect 31484 16736 31536 16788
rect 37924 16736 37976 16788
rect 25780 16575 25832 16584
rect 25780 16541 25789 16575
rect 25789 16541 25823 16575
rect 25823 16541 25832 16575
rect 25780 16532 25832 16541
rect 25872 16575 25924 16584
rect 25872 16541 25881 16575
rect 25881 16541 25915 16575
rect 25915 16541 25924 16575
rect 25872 16532 25924 16541
rect 20536 16464 20588 16516
rect 21824 16464 21876 16516
rect 16028 16439 16080 16448
rect 16028 16405 16037 16439
rect 16037 16405 16071 16439
rect 16071 16405 16080 16439
rect 16028 16396 16080 16405
rect 17684 16396 17736 16448
rect 18972 16396 19024 16448
rect 21180 16439 21232 16448
rect 21180 16405 21189 16439
rect 21189 16405 21223 16439
rect 21223 16405 21232 16439
rect 21180 16396 21232 16405
rect 22744 16439 22796 16448
rect 22744 16405 22753 16439
rect 22753 16405 22787 16439
rect 22787 16405 22796 16439
rect 22744 16396 22796 16405
rect 23756 16396 23808 16448
rect 24952 16439 25004 16448
rect 24952 16405 24961 16439
rect 24961 16405 24995 16439
rect 24995 16405 25004 16439
rect 24952 16396 25004 16405
rect 26516 16532 26568 16584
rect 27620 16532 27672 16584
rect 27804 16575 27856 16584
rect 27804 16541 27813 16575
rect 27813 16541 27847 16575
rect 27847 16541 27856 16575
rect 27804 16532 27856 16541
rect 28540 16464 28592 16516
rect 29920 16575 29972 16584
rect 29920 16541 29929 16575
rect 29929 16541 29963 16575
rect 29963 16541 29972 16575
rect 29920 16532 29972 16541
rect 30104 16532 30156 16584
rect 31852 16600 31904 16652
rect 34520 16600 34572 16652
rect 38108 16532 38160 16584
rect 30748 16464 30800 16516
rect 26148 16396 26200 16448
rect 26424 16439 26476 16448
rect 26424 16405 26433 16439
rect 26433 16405 26467 16439
rect 26467 16405 26476 16439
rect 26424 16396 26476 16405
rect 29828 16396 29880 16448
rect 30840 16396 30892 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 9680 16235 9732 16244
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 10692 16192 10744 16244
rect 12256 16192 12308 16244
rect 12440 16192 12492 16244
rect 9864 16167 9916 16176
rect 9864 16133 9875 16167
rect 9875 16133 9916 16167
rect 9864 16124 9916 16133
rect 10048 16167 10100 16176
rect 10048 16133 10057 16167
rect 10057 16133 10091 16167
rect 10091 16133 10100 16167
rect 10048 16124 10100 16133
rect 9680 15988 9732 16040
rect 11244 16056 11296 16108
rect 11520 16056 11572 16108
rect 9312 15852 9364 15904
rect 12440 16056 12492 16108
rect 13084 16192 13136 16244
rect 15752 16192 15804 16244
rect 15844 16192 15896 16244
rect 18236 16192 18288 16244
rect 18972 16235 19024 16244
rect 18972 16201 18981 16235
rect 18981 16201 19015 16235
rect 19015 16201 19024 16235
rect 18972 16192 19024 16201
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 17684 16124 17736 16176
rect 19800 16192 19852 16244
rect 21272 16192 21324 16244
rect 21824 16235 21876 16244
rect 21824 16201 21833 16235
rect 21833 16201 21867 16235
rect 21867 16201 21876 16235
rect 21824 16192 21876 16201
rect 22744 16192 22796 16244
rect 24952 16192 25004 16244
rect 27804 16192 27856 16244
rect 14556 15988 14608 16040
rect 15292 15988 15344 16040
rect 16580 15988 16632 16040
rect 17776 16031 17828 16040
rect 12532 15920 12584 15972
rect 16028 15920 16080 15972
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 13728 15895 13780 15904
rect 13728 15861 13737 15895
rect 13737 15861 13771 15895
rect 13771 15861 13780 15895
rect 13728 15852 13780 15861
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 15660 15852 15712 15904
rect 17776 15997 17785 16031
rect 17785 15997 17819 16031
rect 17819 15997 17828 16031
rect 17776 15988 17828 15997
rect 16856 15920 16908 15972
rect 17500 15920 17552 15972
rect 18420 16056 18472 16108
rect 20812 16124 20864 16176
rect 18972 16056 19024 16108
rect 19340 16056 19392 16108
rect 19800 16056 19852 16108
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 20996 16056 21048 16108
rect 21180 16056 21232 16108
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 25228 16124 25280 16176
rect 23296 16056 23348 16108
rect 19064 15920 19116 15972
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 23940 16031 23992 16040
rect 23940 15997 23949 16031
rect 23949 15997 23983 16031
rect 23983 15997 23992 16031
rect 23940 15988 23992 15997
rect 26884 16056 26936 16108
rect 27988 16124 28040 16176
rect 28264 16056 28316 16108
rect 28540 16235 28592 16244
rect 28540 16201 28549 16235
rect 28549 16201 28583 16235
rect 28583 16201 28592 16235
rect 28540 16192 28592 16201
rect 29920 16192 29972 16244
rect 34796 16235 34848 16244
rect 30104 16124 30156 16176
rect 34796 16201 34805 16235
rect 34805 16201 34839 16235
rect 34839 16201 34848 16235
rect 34796 16192 34848 16201
rect 35348 16235 35400 16244
rect 35348 16201 35357 16235
rect 35357 16201 35391 16235
rect 35391 16201 35400 16235
rect 35348 16192 35400 16201
rect 20444 15920 20496 15972
rect 29828 15988 29880 16040
rect 30840 15988 30892 16040
rect 31760 16056 31812 16108
rect 33416 16099 33468 16108
rect 31484 15988 31536 16040
rect 33416 16065 33425 16099
rect 33425 16065 33459 16099
rect 33459 16065 33468 16099
rect 33416 16056 33468 16065
rect 34060 16056 34112 16108
rect 34612 16056 34664 16108
rect 20536 15852 20588 15904
rect 20812 15852 20864 15904
rect 21456 15852 21508 15904
rect 22560 15895 22612 15904
rect 22560 15861 22569 15895
rect 22569 15861 22603 15895
rect 22603 15861 22612 15895
rect 22560 15852 22612 15861
rect 23388 15895 23440 15904
rect 23388 15861 23397 15895
rect 23397 15861 23431 15895
rect 23431 15861 23440 15895
rect 23388 15852 23440 15861
rect 25872 15852 25924 15904
rect 26976 15852 27028 15904
rect 27160 15852 27212 15904
rect 34704 15920 34756 15972
rect 30748 15895 30800 15904
rect 30748 15861 30757 15895
rect 30757 15861 30791 15895
rect 30791 15861 30800 15895
rect 30748 15852 30800 15861
rect 32036 15852 32088 15904
rect 32496 15895 32548 15904
rect 32496 15861 32505 15895
rect 32505 15861 32539 15895
rect 32539 15861 32548 15895
rect 32496 15852 32548 15861
rect 33324 15852 33376 15904
rect 34612 15852 34664 15904
rect 37372 15852 37424 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 11060 15648 11112 15700
rect 9496 15580 9548 15632
rect 9588 15555 9640 15564
rect 9588 15521 9597 15555
rect 9597 15521 9631 15555
rect 9631 15521 9640 15555
rect 9588 15512 9640 15521
rect 7012 15487 7064 15496
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 11152 15623 11204 15632
rect 11152 15589 11161 15623
rect 11161 15589 11195 15623
rect 11195 15589 11204 15623
rect 11152 15580 11204 15589
rect 12164 15648 12216 15700
rect 16028 15648 16080 15700
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 7288 15419 7340 15428
rect 7288 15385 7297 15419
rect 7297 15385 7331 15419
rect 7331 15385 7340 15419
rect 7288 15376 7340 15385
rect 8576 15376 8628 15428
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 11520 15444 11572 15496
rect 14188 15512 14240 15564
rect 15200 15487 15252 15496
rect 15200 15453 15218 15487
rect 15218 15453 15252 15487
rect 15200 15444 15252 15453
rect 15384 15444 15436 15496
rect 17592 15555 17644 15564
rect 17592 15521 17601 15555
rect 17601 15521 17635 15555
rect 17635 15521 17644 15555
rect 17592 15512 17644 15521
rect 17684 15512 17736 15564
rect 20260 15648 20312 15700
rect 21732 15648 21784 15700
rect 22560 15648 22612 15700
rect 23204 15691 23256 15700
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 23388 15648 23440 15700
rect 26608 15648 26660 15700
rect 27804 15648 27856 15700
rect 29920 15648 29972 15700
rect 32496 15648 32548 15700
rect 34060 15648 34112 15700
rect 34704 15648 34756 15700
rect 35348 15648 35400 15700
rect 19524 15512 19576 15564
rect 19800 15512 19852 15564
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 30840 15580 30892 15632
rect 18972 15444 19024 15496
rect 19708 15444 19760 15496
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 9588 15308 9640 15360
rect 11520 15308 11572 15360
rect 14188 15376 14240 15428
rect 14556 15376 14608 15428
rect 14096 15351 14148 15360
rect 14096 15317 14105 15351
rect 14105 15317 14139 15351
rect 14139 15317 14148 15351
rect 14096 15308 14148 15317
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 16580 15376 16632 15428
rect 17500 15376 17552 15428
rect 17684 15351 17736 15360
rect 17684 15317 17693 15351
rect 17693 15317 17727 15351
rect 17727 15317 17736 15351
rect 17684 15308 17736 15317
rect 20076 15308 20128 15360
rect 21456 15444 21508 15496
rect 21732 15487 21784 15496
rect 21732 15453 21741 15487
rect 21741 15453 21775 15487
rect 21775 15453 21784 15487
rect 21732 15444 21784 15453
rect 21640 15419 21692 15428
rect 21640 15385 21649 15419
rect 21649 15385 21683 15419
rect 21683 15385 21692 15419
rect 21640 15376 21692 15385
rect 22192 15376 22244 15428
rect 20628 15351 20680 15360
rect 20628 15317 20637 15351
rect 20637 15317 20671 15351
rect 20671 15317 20680 15351
rect 20628 15308 20680 15317
rect 22652 15444 22704 15496
rect 23020 15487 23072 15496
rect 23020 15453 23029 15487
rect 23029 15453 23063 15487
rect 23063 15453 23072 15487
rect 23020 15444 23072 15453
rect 23296 15487 23348 15496
rect 23296 15453 23305 15487
rect 23305 15453 23339 15487
rect 23339 15453 23348 15487
rect 23296 15444 23348 15453
rect 23480 15444 23532 15496
rect 23940 15444 23992 15496
rect 25136 15444 25188 15496
rect 25688 15444 25740 15496
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 27804 15487 27856 15496
rect 27804 15453 27813 15487
rect 27813 15453 27847 15487
rect 27847 15453 27856 15487
rect 27804 15444 27856 15453
rect 30104 15512 30156 15564
rect 30748 15512 30800 15564
rect 29828 15487 29880 15496
rect 29828 15453 29837 15487
rect 29837 15453 29871 15487
rect 29871 15453 29880 15487
rect 29828 15444 29880 15453
rect 30012 15487 30064 15496
rect 30012 15453 30021 15487
rect 30021 15453 30055 15487
rect 30055 15453 30064 15487
rect 30012 15444 30064 15453
rect 24492 15376 24544 15428
rect 24860 15376 24912 15428
rect 25320 15376 25372 15428
rect 26516 15419 26568 15428
rect 26516 15385 26525 15419
rect 26525 15385 26559 15419
rect 26559 15385 26568 15419
rect 26516 15376 26568 15385
rect 31300 15487 31352 15496
rect 31300 15453 31309 15487
rect 31309 15453 31343 15487
rect 31343 15453 31352 15487
rect 31300 15444 31352 15453
rect 31484 15444 31536 15496
rect 32036 15487 32088 15496
rect 32036 15453 32070 15487
rect 32070 15453 32088 15487
rect 32036 15444 32088 15453
rect 33784 15487 33836 15496
rect 33784 15453 33793 15487
rect 33793 15453 33827 15487
rect 33827 15453 33836 15487
rect 33784 15444 33836 15453
rect 33876 15444 33928 15496
rect 22744 15351 22796 15360
rect 22744 15317 22753 15351
rect 22753 15317 22787 15351
rect 22787 15317 22796 15351
rect 22744 15308 22796 15317
rect 23572 15351 23624 15360
rect 23572 15317 23581 15351
rect 23581 15317 23615 15351
rect 23615 15317 23624 15351
rect 23572 15308 23624 15317
rect 26792 15308 26844 15360
rect 27528 15308 27580 15360
rect 28448 15351 28500 15360
rect 28448 15317 28457 15351
rect 28457 15317 28491 15351
rect 28491 15317 28500 15351
rect 28448 15308 28500 15317
rect 29552 15351 29604 15360
rect 29552 15317 29561 15351
rect 29561 15317 29595 15351
rect 29595 15317 29604 15351
rect 29552 15308 29604 15317
rect 29920 15308 29972 15360
rect 30932 15351 30984 15360
rect 30932 15317 30941 15351
rect 30941 15317 30975 15351
rect 30975 15317 30984 15351
rect 30932 15308 30984 15317
rect 33324 15376 33376 15428
rect 34336 15444 34388 15496
rect 34612 15444 34664 15496
rect 34796 15444 34848 15496
rect 37372 15487 37424 15496
rect 37372 15453 37381 15487
rect 37381 15453 37415 15487
rect 37415 15453 37424 15487
rect 37372 15444 37424 15453
rect 68284 15444 68336 15496
rect 33232 15351 33284 15360
rect 33232 15317 33241 15351
rect 33241 15317 33275 15351
rect 33275 15317 33284 15351
rect 33232 15308 33284 15317
rect 33692 15308 33744 15360
rect 35348 15376 35400 15428
rect 36452 15351 36504 15360
rect 36452 15317 36461 15351
rect 36461 15317 36495 15351
rect 36495 15317 36504 15351
rect 36452 15308 36504 15317
rect 37280 15351 37332 15360
rect 37280 15317 37289 15351
rect 37289 15317 37323 15351
rect 37323 15317 37332 15351
rect 37280 15308 37332 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 7288 15104 7340 15156
rect 8576 15147 8628 15156
rect 8576 15113 8585 15147
rect 8585 15113 8619 15147
rect 8619 15113 8628 15147
rect 8576 15104 8628 15113
rect 9036 15104 9088 15156
rect 9680 15147 9732 15156
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 9588 15036 9640 15088
rect 9956 15036 10008 15088
rect 8668 15011 8720 15020
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 11336 15036 11388 15088
rect 11152 14968 11204 15020
rect 12624 15104 12676 15156
rect 12716 15104 12768 15156
rect 14188 15147 14240 15156
rect 14188 15113 14197 15147
rect 14197 15113 14231 15147
rect 14231 15113 14240 15147
rect 14188 15104 14240 15113
rect 11888 15036 11940 15088
rect 12256 15036 12308 15088
rect 12900 14968 12952 15020
rect 12992 14968 13044 15020
rect 14096 15036 14148 15088
rect 12716 14900 12768 14952
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 15936 15104 15988 15156
rect 15752 14968 15804 15020
rect 15844 15011 15896 15020
rect 15844 14977 15853 15011
rect 15853 14977 15887 15011
rect 15887 14977 15896 15011
rect 15844 14968 15896 14977
rect 16580 14968 16632 15020
rect 17500 15104 17552 15156
rect 19248 15104 19300 15156
rect 19432 15104 19484 15156
rect 19524 15104 19576 15156
rect 20076 15104 20128 15156
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 20628 15036 20680 15088
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 23756 15147 23808 15156
rect 23756 15113 23765 15147
rect 23765 15113 23799 15147
rect 23799 15113 23808 15147
rect 23756 15104 23808 15113
rect 24492 15104 24544 15156
rect 30012 15104 30064 15156
rect 30932 15104 30984 15156
rect 33784 15104 33836 15156
rect 35348 15147 35400 15156
rect 35348 15113 35357 15147
rect 35357 15113 35391 15147
rect 35391 15113 35400 15147
rect 35348 15104 35400 15113
rect 36452 15104 36504 15156
rect 37096 15104 37148 15156
rect 20444 15011 20496 15020
rect 20444 14977 20453 15011
rect 20453 14977 20487 15011
rect 20487 14977 20496 15011
rect 20444 14968 20496 14977
rect 20536 15011 20588 15020
rect 20536 14977 20545 15011
rect 20545 14977 20579 15011
rect 20579 14977 20588 15011
rect 20536 14968 20588 14977
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 23572 14968 23624 15020
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 25044 15036 25096 15088
rect 26148 15036 26200 15088
rect 26792 15036 26844 15088
rect 29552 15036 29604 15088
rect 11060 14764 11112 14816
rect 12164 14764 12216 14816
rect 12440 14832 12492 14884
rect 13084 14764 13136 14816
rect 14740 14875 14792 14884
rect 14740 14841 14749 14875
rect 14749 14841 14783 14875
rect 14783 14841 14792 14875
rect 14740 14832 14792 14841
rect 15292 14832 15344 14884
rect 15200 14764 15252 14816
rect 17040 14943 17092 14952
rect 17040 14909 17049 14943
rect 17049 14909 17083 14943
rect 17083 14909 17092 14943
rect 17040 14900 17092 14909
rect 18788 14943 18840 14952
rect 18788 14909 18797 14943
rect 18797 14909 18831 14943
rect 18831 14909 18840 14943
rect 18788 14900 18840 14909
rect 18972 14832 19024 14884
rect 19156 14832 19208 14884
rect 21640 14900 21692 14952
rect 24492 15011 24544 15020
rect 24492 14977 24501 15011
rect 24501 14977 24535 15011
rect 24535 14977 24544 15011
rect 24492 14968 24544 14977
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 25504 14968 25556 15020
rect 27068 14968 27120 15020
rect 27528 15011 27580 15020
rect 27528 14977 27537 15011
rect 27537 14977 27571 15011
rect 27571 14977 27580 15011
rect 27528 14968 27580 14977
rect 27620 14968 27672 15020
rect 27988 14968 28040 15020
rect 28172 14968 28224 15020
rect 25412 14900 25464 14952
rect 18880 14764 18932 14816
rect 24584 14875 24636 14884
rect 24584 14841 24593 14875
rect 24593 14841 24627 14875
rect 24627 14841 24636 14875
rect 24584 14832 24636 14841
rect 25596 14832 25648 14884
rect 19984 14764 20036 14816
rect 20076 14807 20128 14816
rect 20076 14773 20085 14807
rect 20085 14773 20119 14807
rect 20119 14773 20128 14807
rect 20076 14764 20128 14773
rect 25412 14764 25464 14816
rect 26332 14900 26384 14952
rect 31760 15036 31812 15088
rect 33232 15079 33284 15088
rect 33232 15045 33250 15079
rect 33250 15045 33284 15079
rect 34336 15079 34388 15088
rect 33232 15036 33284 15045
rect 30748 14900 30800 14952
rect 31300 14900 31352 14952
rect 25780 14832 25832 14884
rect 25872 14764 25924 14816
rect 26516 14764 26568 14816
rect 27436 14807 27488 14816
rect 27436 14773 27445 14807
rect 27445 14773 27479 14807
rect 27479 14773 27488 14807
rect 27436 14764 27488 14773
rect 27804 14807 27856 14816
rect 27804 14773 27813 14807
rect 27813 14773 27847 14807
rect 27847 14773 27856 14807
rect 27804 14764 27856 14773
rect 30656 14807 30708 14816
rect 30656 14773 30665 14807
rect 30665 14773 30699 14807
rect 30699 14773 30708 14807
rect 30656 14764 30708 14773
rect 30840 14807 30892 14816
rect 30840 14773 30849 14807
rect 30849 14773 30883 14807
rect 30883 14773 30892 14807
rect 30840 14764 30892 14773
rect 33416 14968 33468 15020
rect 34336 15045 34345 15079
rect 34345 15045 34379 15079
rect 34379 15045 34388 15079
rect 34336 15036 34388 15045
rect 33600 15011 33652 15020
rect 33600 14977 33609 15011
rect 33609 14977 33643 15011
rect 33643 14977 33652 15011
rect 33600 14968 33652 14977
rect 32588 14764 32640 14816
rect 35716 14968 35768 15020
rect 67640 14900 67692 14952
rect 37280 14764 37332 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 10876 14560 10928 14612
rect 11428 14560 11480 14612
rect 12072 14560 12124 14612
rect 14740 14560 14792 14612
rect 15660 14560 15712 14612
rect 15844 14560 15896 14612
rect 17040 14560 17092 14612
rect 19156 14560 19208 14612
rect 11060 14492 11112 14544
rect 12164 14492 12216 14544
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 9496 14356 9548 14408
rect 10140 14356 10192 14408
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 12072 14467 12124 14476
rect 12072 14433 12081 14467
rect 12081 14433 12115 14467
rect 12115 14433 12124 14467
rect 12072 14424 12124 14433
rect 11888 14356 11940 14408
rect 18512 14492 18564 14544
rect 20076 14560 20128 14612
rect 19432 14492 19484 14544
rect 21640 14560 21692 14612
rect 24492 14560 24544 14612
rect 25136 14560 25188 14612
rect 25688 14560 25740 14612
rect 26056 14560 26108 14612
rect 16856 14467 16908 14476
rect 16856 14433 16865 14467
rect 16865 14433 16899 14467
rect 16899 14433 16908 14467
rect 16856 14424 16908 14433
rect 17408 14424 17460 14476
rect 18788 14424 18840 14476
rect 11980 14288 12032 14340
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 11336 14220 11388 14272
rect 11428 14220 11480 14272
rect 12900 14288 12952 14340
rect 12992 14331 13044 14340
rect 12992 14297 13001 14331
rect 13001 14297 13035 14331
rect 13035 14297 13044 14331
rect 12992 14288 13044 14297
rect 13084 14288 13136 14340
rect 12808 14220 12860 14272
rect 15108 14356 15160 14408
rect 15384 14356 15436 14408
rect 14924 14288 14976 14340
rect 17316 14356 17368 14408
rect 18144 14399 18196 14408
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 20260 14424 20312 14476
rect 19524 14356 19576 14408
rect 14188 14220 14240 14272
rect 17592 14263 17644 14272
rect 17592 14229 17601 14263
rect 17601 14229 17635 14263
rect 17635 14229 17644 14263
rect 17592 14220 17644 14229
rect 19708 14220 19760 14272
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 20076 14356 20128 14408
rect 24584 14492 24636 14544
rect 20444 14220 20496 14272
rect 22744 14356 22796 14408
rect 23020 14356 23072 14408
rect 24952 14492 25004 14544
rect 24860 14424 24912 14476
rect 26792 14424 26844 14476
rect 22100 14288 22152 14340
rect 24768 14356 24820 14408
rect 27436 14560 27488 14612
rect 27344 14424 27396 14476
rect 27620 14492 27672 14544
rect 28172 14535 28224 14544
rect 28172 14501 28181 14535
rect 28181 14501 28215 14535
rect 28215 14501 28224 14535
rect 28172 14492 28224 14501
rect 25688 14288 25740 14340
rect 24676 14220 24728 14272
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 26700 14263 26752 14272
rect 26700 14229 26709 14263
rect 26709 14229 26743 14263
rect 26743 14229 26752 14263
rect 26700 14220 26752 14229
rect 27620 14288 27672 14340
rect 28448 14356 28500 14408
rect 29552 14220 29604 14272
rect 29644 14220 29696 14272
rect 30380 14356 30432 14408
rect 30840 14560 30892 14612
rect 35716 14560 35768 14612
rect 33600 14492 33652 14544
rect 33784 14356 33836 14408
rect 33508 14288 33560 14340
rect 35348 14288 35400 14340
rect 31944 14220 31996 14272
rect 34336 14220 34388 14272
rect 36084 14220 36136 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 9128 14016 9180 14068
rect 7012 13880 7064 13932
rect 8116 13948 8168 14000
rect 8576 13948 8628 14000
rect 10140 14059 10192 14068
rect 10140 14025 10149 14059
rect 10149 14025 10183 14059
rect 10183 14025 10192 14059
rect 10140 14016 10192 14025
rect 10968 14016 11020 14068
rect 10692 13991 10744 14000
rect 9956 13880 10008 13932
rect 10692 13957 10714 13991
rect 10714 13957 10744 13991
rect 10692 13948 10744 13957
rect 10876 13991 10928 14000
rect 10876 13957 10885 13991
rect 10885 13957 10919 13991
rect 10919 13957 10928 13991
rect 10876 13948 10928 13957
rect 8944 13744 8996 13796
rect 12256 14016 12308 14068
rect 17592 14016 17644 14068
rect 18144 14016 18196 14068
rect 12900 13991 12952 14000
rect 12900 13957 12909 13991
rect 12909 13957 12943 13991
rect 12943 13957 12952 13991
rect 12900 13948 12952 13957
rect 13912 13948 13964 14000
rect 14924 13948 14976 14000
rect 15108 13948 15160 14000
rect 11888 13744 11940 13796
rect 15200 13923 15252 13932
rect 15200 13889 15209 13923
rect 15209 13889 15243 13923
rect 15243 13889 15252 13923
rect 15200 13880 15252 13889
rect 18512 13948 18564 14000
rect 17684 13880 17736 13932
rect 18236 13880 18288 13932
rect 20628 14016 20680 14068
rect 21088 14016 21140 14068
rect 19984 13991 20036 14000
rect 19984 13957 20002 13991
rect 20002 13957 20036 13991
rect 19984 13948 20036 13957
rect 19432 13880 19484 13932
rect 14188 13744 14240 13796
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 20260 13855 20312 13864
rect 20260 13821 20269 13855
rect 20269 13821 20303 13855
rect 20303 13821 20312 13855
rect 20260 13812 20312 13821
rect 20444 13812 20496 13864
rect 23664 14016 23716 14068
rect 24860 14016 24912 14068
rect 25412 14016 25464 14068
rect 26332 14016 26384 14068
rect 23112 13880 23164 13932
rect 24768 13948 24820 14000
rect 29644 14016 29696 14068
rect 17224 13719 17276 13728
rect 17224 13685 17233 13719
rect 17233 13685 17267 13719
rect 17267 13685 17276 13719
rect 17224 13676 17276 13685
rect 17868 13676 17920 13728
rect 23020 13812 23072 13864
rect 23480 13855 23532 13864
rect 23480 13821 23489 13855
rect 23489 13821 23523 13855
rect 23523 13821 23532 13855
rect 23480 13812 23532 13821
rect 22468 13744 22520 13796
rect 25044 13880 25096 13932
rect 25228 13880 25280 13932
rect 25504 13880 25556 13932
rect 25872 13880 25924 13932
rect 25780 13812 25832 13864
rect 26424 13880 26476 13932
rect 26700 13923 26752 13932
rect 26700 13889 26709 13923
rect 26709 13889 26743 13923
rect 26743 13889 26752 13923
rect 26700 13880 26752 13889
rect 26976 13923 27028 13932
rect 26976 13889 26985 13923
rect 26985 13889 27019 13923
rect 27019 13889 27028 13923
rect 26976 13880 27028 13889
rect 27252 13923 27304 13932
rect 27252 13889 27286 13923
rect 27286 13889 27304 13923
rect 27252 13880 27304 13889
rect 29552 13948 29604 14000
rect 33784 14016 33836 14068
rect 32588 13923 32640 13932
rect 32588 13889 32597 13923
rect 32597 13889 32631 13923
rect 32631 13889 32640 13923
rect 32588 13880 32640 13889
rect 34336 13948 34388 14000
rect 35440 13880 35492 13932
rect 36176 13923 36228 13932
rect 36176 13889 36185 13923
rect 36185 13889 36219 13923
rect 36219 13889 36228 13923
rect 36176 13880 36228 13889
rect 25964 13744 26016 13796
rect 30564 13744 30616 13796
rect 31208 13812 31260 13864
rect 32680 13855 32732 13864
rect 32680 13821 32689 13855
rect 32689 13821 32723 13855
rect 32723 13821 32732 13855
rect 32680 13812 32732 13821
rect 34796 13855 34848 13864
rect 34796 13821 34805 13855
rect 34805 13821 34839 13855
rect 34839 13821 34848 13855
rect 34796 13812 34848 13821
rect 26056 13676 26108 13728
rect 28356 13719 28408 13728
rect 28356 13685 28365 13719
rect 28365 13685 28399 13719
rect 28399 13685 28408 13719
rect 28356 13676 28408 13685
rect 31024 13719 31076 13728
rect 31024 13685 31033 13719
rect 31033 13685 31067 13719
rect 31067 13685 31076 13719
rect 31024 13676 31076 13685
rect 33140 13719 33192 13728
rect 33140 13685 33149 13719
rect 33149 13685 33183 13719
rect 33183 13685 33192 13719
rect 33140 13676 33192 13685
rect 34152 13676 34204 13728
rect 35348 13812 35400 13864
rect 36360 13812 36412 13864
rect 36268 13676 36320 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 9956 13472 10008 13524
rect 10692 13472 10744 13524
rect 11060 13404 11112 13456
rect 8668 13268 8720 13320
rect 10416 13268 10468 13320
rect 9588 13200 9640 13252
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 12532 13515 12584 13524
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 13912 13472 13964 13524
rect 17960 13515 18012 13524
rect 17960 13481 17969 13515
rect 17969 13481 18003 13515
rect 18003 13481 18012 13515
rect 17960 13472 18012 13481
rect 18512 13472 18564 13524
rect 22836 13472 22888 13524
rect 30380 13515 30432 13524
rect 30380 13481 30389 13515
rect 30389 13481 30423 13515
rect 30423 13481 30432 13515
rect 30380 13472 30432 13481
rect 30656 13472 30708 13524
rect 31024 13472 31076 13524
rect 34428 13472 34480 13524
rect 34796 13472 34848 13524
rect 35440 13472 35492 13524
rect 12164 13404 12216 13456
rect 11336 13336 11388 13345
rect 12808 13336 12860 13388
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 11060 13311 11112 13320
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 8944 13132 8996 13184
rect 10692 13132 10744 13184
rect 11704 13268 11756 13320
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 13084 13404 13136 13456
rect 29092 13404 29144 13456
rect 13820 13336 13872 13388
rect 13636 13268 13688 13320
rect 15108 13379 15160 13388
rect 15108 13345 15117 13379
rect 15117 13345 15151 13379
rect 15151 13345 15160 13379
rect 15108 13336 15160 13345
rect 20260 13336 20312 13388
rect 22468 13336 22520 13388
rect 23756 13336 23808 13388
rect 26976 13379 27028 13388
rect 26976 13345 26985 13379
rect 26985 13345 27019 13379
rect 27019 13345 27028 13379
rect 26976 13336 27028 13345
rect 28356 13336 28408 13388
rect 33508 13336 33560 13388
rect 17224 13268 17276 13320
rect 17868 13268 17920 13320
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 20444 13311 20496 13320
rect 20444 13277 20453 13311
rect 20453 13277 20487 13311
rect 20487 13277 20496 13311
rect 20444 13268 20496 13277
rect 27620 13268 27672 13320
rect 29920 13268 29972 13320
rect 15384 13243 15436 13252
rect 15384 13209 15418 13243
rect 15418 13209 15436 13243
rect 15384 13200 15436 13209
rect 21456 13200 21508 13252
rect 30564 13268 30616 13320
rect 36176 13404 36228 13456
rect 30932 13311 30984 13320
rect 30932 13277 30941 13311
rect 30941 13277 30975 13311
rect 30975 13277 30984 13311
rect 30932 13268 30984 13277
rect 35532 13268 35584 13320
rect 36360 13336 36412 13388
rect 36268 13268 36320 13320
rect 12164 13132 12216 13184
rect 16948 13132 17000 13184
rect 18236 13132 18288 13184
rect 21824 13132 21876 13184
rect 22836 13175 22888 13184
rect 22836 13141 22845 13175
rect 22845 13141 22879 13175
rect 22879 13141 22888 13175
rect 22836 13132 22888 13141
rect 28172 13175 28224 13184
rect 28172 13141 28181 13175
rect 28181 13141 28215 13175
rect 28215 13141 28224 13175
rect 28172 13132 28224 13141
rect 30104 13132 30156 13184
rect 32496 13243 32548 13252
rect 32496 13209 32505 13243
rect 32505 13209 32539 13243
rect 32539 13209 32548 13243
rect 32496 13200 32548 13209
rect 33140 13200 33192 13252
rect 34152 13243 34204 13252
rect 34152 13209 34161 13243
rect 34161 13209 34195 13243
rect 34195 13209 34204 13243
rect 34152 13200 34204 13209
rect 34612 13200 34664 13252
rect 35808 13243 35860 13252
rect 35808 13209 35817 13243
rect 35817 13209 35851 13243
rect 35851 13209 35860 13243
rect 35808 13200 35860 13209
rect 35992 13200 36044 13252
rect 36176 13243 36228 13252
rect 36176 13209 36185 13243
rect 36185 13209 36219 13243
rect 36219 13209 36228 13243
rect 36176 13200 36228 13209
rect 36728 13175 36780 13184
rect 36728 13141 36737 13175
rect 36737 13141 36771 13175
rect 36771 13141 36780 13175
rect 36728 13132 36780 13141
rect 36820 13132 36872 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 8300 12792 8352 12844
rect 11888 12928 11940 12980
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 8944 12860 8996 12912
rect 9680 12860 9732 12912
rect 11060 12860 11112 12912
rect 17868 12928 17920 12980
rect 15108 12860 15160 12912
rect 11704 12792 11756 12844
rect 10692 12724 10744 12776
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 15476 12792 15528 12844
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 17868 12835 17920 12844
rect 17868 12801 17877 12835
rect 17877 12801 17911 12835
rect 17911 12801 17920 12835
rect 17868 12792 17920 12801
rect 18144 12928 18196 12980
rect 20444 12971 20496 12980
rect 20444 12937 20453 12971
rect 20453 12937 20487 12971
rect 20487 12937 20496 12971
rect 20444 12928 20496 12937
rect 20628 12928 20680 12980
rect 20904 12928 20956 12980
rect 21456 12971 21508 12980
rect 21456 12937 21465 12971
rect 21465 12937 21499 12971
rect 21499 12937 21508 12971
rect 21456 12928 21508 12937
rect 22836 12928 22888 12980
rect 20260 12860 20312 12912
rect 18236 12792 18288 12844
rect 23112 12792 23164 12844
rect 23480 12792 23532 12844
rect 25964 12860 26016 12912
rect 28356 12860 28408 12912
rect 29092 12860 29144 12912
rect 13636 12724 13688 12776
rect 15384 12724 15436 12776
rect 17776 12724 17828 12776
rect 20904 12724 20956 12776
rect 21548 12724 21600 12776
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 22100 12724 22152 12733
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 12348 12631 12400 12640
rect 12348 12597 12357 12631
rect 12357 12597 12391 12631
rect 12391 12597 12400 12631
rect 12348 12588 12400 12597
rect 17592 12631 17644 12640
rect 17592 12597 17601 12631
rect 17601 12597 17635 12631
rect 17635 12597 17644 12631
rect 17592 12588 17644 12597
rect 19616 12631 19668 12640
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 26148 12724 26200 12776
rect 26792 12724 26844 12776
rect 28540 12724 28592 12776
rect 29092 12767 29144 12776
rect 29092 12733 29101 12767
rect 29101 12733 29135 12767
rect 29135 12733 29144 12767
rect 29092 12724 29144 12733
rect 32496 12928 32548 12980
rect 34428 12928 34480 12980
rect 30656 12903 30708 12912
rect 30656 12869 30665 12903
rect 30665 12869 30699 12903
rect 30699 12869 30708 12903
rect 30656 12860 30708 12869
rect 30380 12835 30432 12844
rect 30380 12801 30389 12835
rect 30389 12801 30423 12835
rect 30423 12801 30432 12835
rect 30380 12792 30432 12801
rect 30932 12835 30984 12844
rect 30932 12801 30941 12835
rect 30941 12801 30975 12835
rect 30975 12801 30984 12835
rect 30932 12792 30984 12801
rect 31208 12835 31260 12844
rect 31208 12801 31217 12835
rect 31217 12801 31251 12835
rect 31251 12801 31260 12835
rect 31208 12792 31260 12801
rect 34152 12860 34204 12912
rect 24952 12656 25004 12708
rect 25412 12631 25464 12640
rect 25412 12597 25421 12631
rect 25421 12597 25455 12631
rect 25455 12597 25464 12631
rect 25412 12588 25464 12597
rect 26056 12699 26108 12708
rect 26056 12665 26065 12699
rect 26065 12665 26099 12699
rect 26099 12665 26108 12699
rect 26056 12656 26108 12665
rect 28264 12588 28316 12640
rect 28540 12588 28592 12640
rect 29184 12631 29236 12640
rect 29184 12597 29193 12631
rect 29193 12597 29227 12631
rect 29227 12597 29236 12631
rect 29184 12588 29236 12597
rect 30656 12631 30708 12640
rect 30656 12597 30665 12631
rect 30665 12597 30699 12631
rect 30699 12597 30708 12631
rect 30656 12588 30708 12597
rect 31392 12588 31444 12640
rect 34244 12792 34296 12844
rect 34428 12656 34480 12708
rect 35808 12928 35860 12980
rect 35900 12860 35952 12912
rect 36360 12860 36412 12912
rect 34796 12724 34848 12776
rect 33968 12588 34020 12640
rect 34520 12588 34572 12640
rect 35348 12767 35400 12776
rect 35348 12733 35357 12767
rect 35357 12733 35391 12767
rect 35391 12733 35400 12767
rect 35348 12724 35400 12733
rect 36820 12588 36872 12640
rect 37280 12631 37332 12640
rect 37280 12597 37289 12631
rect 37289 12597 37323 12631
rect 37323 12597 37332 12631
rect 37280 12588 37332 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 9680 12384 9732 12436
rect 13636 12384 13688 12436
rect 15476 12384 15528 12436
rect 20076 12384 20128 12436
rect 17868 12316 17920 12368
rect 20720 12384 20772 12436
rect 22100 12384 22152 12436
rect 11888 12248 11940 12300
rect 12348 12248 12400 12300
rect 11520 12180 11572 12232
rect 17132 12180 17184 12232
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 9588 12112 9640 12164
rect 12992 12112 13044 12164
rect 16488 12112 16540 12164
rect 20628 12316 20680 12368
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 19616 12180 19668 12189
rect 20076 12180 20128 12232
rect 20904 12112 20956 12164
rect 21364 12155 21416 12164
rect 21364 12121 21373 12155
rect 21373 12121 21407 12155
rect 21407 12121 21416 12155
rect 21364 12112 21416 12121
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 18328 12044 18380 12096
rect 18420 12044 18472 12096
rect 19340 12044 19392 12096
rect 19984 12087 20036 12096
rect 19984 12053 19993 12087
rect 19993 12053 20027 12087
rect 20027 12053 20036 12087
rect 19984 12044 20036 12053
rect 21824 12223 21876 12232
rect 21824 12189 21833 12223
rect 21833 12189 21867 12223
rect 21867 12189 21876 12223
rect 21824 12180 21876 12189
rect 21916 12180 21968 12232
rect 22192 12044 22244 12096
rect 23112 12180 23164 12232
rect 25964 12384 26016 12436
rect 26700 12384 26752 12436
rect 30380 12384 30432 12436
rect 33692 12384 33744 12436
rect 34152 12427 34204 12436
rect 34152 12393 34161 12427
rect 34161 12393 34195 12427
rect 34195 12393 34204 12427
rect 34152 12384 34204 12393
rect 34244 12384 34296 12436
rect 35900 12427 35952 12436
rect 35900 12393 35909 12427
rect 35909 12393 35943 12427
rect 35943 12393 35952 12427
rect 35900 12384 35952 12393
rect 36360 12427 36412 12436
rect 36360 12393 36369 12427
rect 36369 12393 36403 12427
rect 36403 12393 36412 12427
rect 36360 12384 36412 12393
rect 25044 12291 25096 12300
rect 25044 12257 25053 12291
rect 25053 12257 25087 12291
rect 25087 12257 25096 12291
rect 25044 12248 25096 12257
rect 27252 12248 27304 12300
rect 29000 12248 29052 12300
rect 24952 12180 25004 12232
rect 27712 12223 27764 12232
rect 27712 12189 27721 12223
rect 27721 12189 27755 12223
rect 27755 12189 27764 12223
rect 27712 12180 27764 12189
rect 28540 12180 28592 12232
rect 25320 12155 25372 12164
rect 25320 12121 25329 12155
rect 25329 12121 25363 12155
rect 25363 12121 25372 12155
rect 25320 12112 25372 12121
rect 25596 12112 25648 12164
rect 29092 12223 29144 12232
rect 29092 12189 29101 12223
rect 29101 12189 29135 12223
rect 29135 12189 29144 12223
rect 29092 12180 29144 12189
rect 30748 12112 30800 12164
rect 30932 12180 30984 12232
rect 31208 12180 31260 12232
rect 32680 12316 32732 12368
rect 33324 12316 33376 12368
rect 33876 12316 33928 12368
rect 33968 12316 34020 12368
rect 32864 12248 32916 12300
rect 34520 12248 34572 12300
rect 24768 12044 24820 12096
rect 25688 12044 25740 12096
rect 31116 12044 31168 12096
rect 31300 12044 31352 12096
rect 32956 12180 33008 12232
rect 33416 12180 33468 12232
rect 31760 12044 31812 12096
rect 31852 12087 31904 12096
rect 31852 12053 31861 12087
rect 31861 12053 31895 12087
rect 31895 12053 31904 12087
rect 31852 12044 31904 12053
rect 32588 12087 32640 12096
rect 32588 12053 32597 12087
rect 32597 12053 32631 12087
rect 32631 12053 32640 12087
rect 32588 12044 32640 12053
rect 33600 12087 33652 12096
rect 33600 12053 33609 12087
rect 33609 12053 33643 12087
rect 33643 12053 33652 12087
rect 33600 12044 33652 12053
rect 33876 12223 33928 12232
rect 33876 12189 33885 12223
rect 33885 12189 33919 12223
rect 33919 12189 33928 12223
rect 33876 12180 33928 12189
rect 34244 12223 34296 12232
rect 34244 12189 34253 12223
rect 34253 12189 34287 12223
rect 34287 12189 34296 12223
rect 34244 12180 34296 12189
rect 35532 12316 35584 12368
rect 35440 12180 35492 12232
rect 37280 12248 37332 12300
rect 35992 12180 36044 12232
rect 36084 12180 36136 12232
rect 36268 12223 36320 12232
rect 36268 12189 36277 12223
rect 36277 12189 36311 12223
rect 36311 12189 36320 12223
rect 36268 12180 36320 12189
rect 36636 12180 36688 12232
rect 35256 12112 35308 12164
rect 34796 12044 34848 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 12992 11840 13044 11892
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 17960 11840 18012 11892
rect 15476 11772 15528 11824
rect 16488 11772 16540 11824
rect 9588 11704 9640 11756
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 17500 11704 17552 11756
rect 21364 11840 21416 11892
rect 22560 11840 22612 11892
rect 24952 11840 25004 11892
rect 25044 11840 25096 11892
rect 25320 11883 25372 11892
rect 25320 11849 25329 11883
rect 25329 11849 25363 11883
rect 25363 11849 25372 11883
rect 25320 11840 25372 11849
rect 19708 11772 19760 11824
rect 21824 11815 21876 11824
rect 21824 11781 21833 11815
rect 21833 11781 21867 11815
rect 21867 11781 21876 11815
rect 21824 11772 21876 11781
rect 22468 11772 22520 11824
rect 23940 11772 23992 11824
rect 14648 11636 14700 11688
rect 17868 11636 17920 11688
rect 21732 11704 21784 11756
rect 21916 11704 21968 11756
rect 21824 11636 21876 11688
rect 13820 11568 13872 11620
rect 18788 11568 18840 11620
rect 22192 11679 22244 11688
rect 22192 11645 22201 11679
rect 22201 11645 22235 11679
rect 22235 11645 22244 11679
rect 22192 11636 22244 11645
rect 22284 11636 22336 11688
rect 25228 11704 25280 11756
rect 25596 11772 25648 11824
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 26792 11883 26844 11892
rect 26792 11849 26801 11883
rect 26801 11849 26835 11883
rect 26835 11849 26844 11883
rect 26792 11840 26844 11849
rect 28172 11840 28224 11892
rect 30748 11883 30800 11892
rect 30748 11849 30757 11883
rect 30757 11849 30791 11883
rect 30791 11849 30800 11883
rect 30748 11840 30800 11849
rect 31300 11840 31352 11892
rect 33140 11883 33192 11892
rect 33140 11849 33149 11883
rect 33149 11849 33183 11883
rect 33183 11849 33192 11883
rect 33140 11840 33192 11849
rect 30012 11772 30064 11824
rect 34612 11840 34664 11892
rect 27160 11747 27212 11756
rect 24860 11636 24912 11688
rect 27160 11713 27169 11747
rect 27169 11713 27203 11747
rect 27203 11713 27212 11747
rect 27160 11704 27212 11713
rect 29000 11747 29052 11756
rect 29000 11713 29009 11747
rect 29009 11713 29043 11747
rect 29043 11713 29052 11747
rect 29000 11704 29052 11713
rect 11612 11543 11664 11552
rect 11612 11509 11621 11543
rect 11621 11509 11655 11543
rect 11655 11509 11664 11543
rect 11612 11500 11664 11509
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 18052 11500 18104 11552
rect 18144 11543 18196 11552
rect 18144 11509 18153 11543
rect 18153 11509 18187 11543
rect 18187 11509 18196 11543
rect 18144 11500 18196 11509
rect 18696 11500 18748 11552
rect 22376 11568 22428 11620
rect 20904 11543 20956 11552
rect 20904 11509 20913 11543
rect 20913 11509 20947 11543
rect 20947 11509 20956 11543
rect 20904 11500 20956 11509
rect 25228 11500 25280 11552
rect 25964 11568 26016 11620
rect 28080 11679 28132 11688
rect 28080 11645 28089 11679
rect 28089 11645 28123 11679
rect 28123 11645 28132 11679
rect 28816 11679 28868 11688
rect 28080 11636 28132 11645
rect 28816 11645 28825 11679
rect 28825 11645 28859 11679
rect 28859 11645 28868 11679
rect 28816 11636 28868 11645
rect 30656 11636 30708 11688
rect 30288 11500 30340 11552
rect 31024 11543 31076 11552
rect 31024 11509 31033 11543
rect 31033 11509 31067 11543
rect 31067 11509 31076 11543
rect 31024 11500 31076 11509
rect 31300 11747 31352 11756
rect 31300 11713 31309 11747
rect 31309 11713 31343 11747
rect 31343 11713 31352 11747
rect 31300 11704 31352 11713
rect 33416 11772 33468 11824
rect 35256 11883 35308 11892
rect 35256 11849 35265 11883
rect 35265 11849 35299 11883
rect 35299 11849 35308 11883
rect 35256 11840 35308 11849
rect 35440 11840 35492 11892
rect 32772 11747 32824 11756
rect 32772 11713 32781 11747
rect 32781 11713 32815 11747
rect 32815 11713 32824 11747
rect 32772 11704 32824 11713
rect 32864 11704 32916 11756
rect 33140 11747 33192 11756
rect 33140 11713 33178 11747
rect 33178 11713 33192 11747
rect 33140 11704 33192 11713
rect 33692 11704 33744 11756
rect 34796 11704 34848 11756
rect 31392 11636 31444 11688
rect 31668 11679 31720 11688
rect 31668 11645 31677 11679
rect 31677 11645 31711 11679
rect 31711 11645 31720 11679
rect 31668 11636 31720 11645
rect 33232 11568 33284 11620
rect 31760 11500 31812 11552
rect 32496 11543 32548 11552
rect 32496 11509 32505 11543
rect 32505 11509 32539 11543
rect 32539 11509 32548 11543
rect 32496 11500 32548 11509
rect 32772 11500 32824 11552
rect 32864 11543 32916 11552
rect 32864 11509 32873 11543
rect 32873 11509 32907 11543
rect 32907 11509 32916 11543
rect 32864 11500 32916 11509
rect 34428 11636 34480 11688
rect 33600 11543 33652 11552
rect 33600 11509 33609 11543
rect 33609 11509 33643 11543
rect 33643 11509 33652 11543
rect 33600 11500 33652 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 10692 11296 10744 11348
rect 18144 11296 18196 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19340 11296 19392 11348
rect 19708 11339 19760 11348
rect 19708 11305 19717 11339
rect 19717 11305 19751 11339
rect 19751 11305 19760 11339
rect 19708 11296 19760 11305
rect 20628 11296 20680 11348
rect 21732 11296 21784 11348
rect 23940 11339 23992 11348
rect 23940 11305 23949 11339
rect 23949 11305 23983 11339
rect 23983 11305 23992 11339
rect 23940 11296 23992 11305
rect 24860 11296 24912 11348
rect 25964 11296 26016 11348
rect 18052 11228 18104 11280
rect 11612 11092 11664 11144
rect 12164 11092 12216 11144
rect 14648 11092 14700 11144
rect 17132 11092 17184 11144
rect 16396 11024 16448 11076
rect 18144 11135 18196 11144
rect 18144 11101 18153 11135
rect 18153 11101 18187 11135
rect 18187 11101 18196 11135
rect 18144 11092 18196 11101
rect 18696 11160 18748 11212
rect 19708 11160 19760 11212
rect 18788 11092 18840 11144
rect 26792 11228 26844 11280
rect 19984 11160 20036 11212
rect 20904 11160 20956 11212
rect 19248 11024 19300 11076
rect 19708 11024 19760 11076
rect 20812 11135 20864 11144
rect 20812 11101 20821 11135
rect 20821 11101 20855 11135
rect 20855 11101 20864 11135
rect 20812 11092 20864 11101
rect 22192 11160 22244 11212
rect 27252 11203 27304 11212
rect 27252 11169 27261 11203
rect 27261 11169 27295 11203
rect 27295 11169 27304 11203
rect 27252 11160 27304 11169
rect 28816 11296 28868 11348
rect 30012 11296 30064 11348
rect 31300 11296 31352 11348
rect 31760 11339 31812 11348
rect 31760 11305 31769 11339
rect 31769 11305 31803 11339
rect 31803 11305 31812 11339
rect 31760 11296 31812 11305
rect 31852 11296 31904 11348
rect 31944 11228 31996 11280
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 21824 11092 21876 11144
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 25504 11135 25556 11144
rect 25504 11101 25513 11135
rect 25513 11101 25547 11135
rect 25547 11101 25556 11135
rect 25504 11092 25556 11101
rect 25780 11092 25832 11144
rect 30288 11160 30340 11212
rect 20720 11024 20772 11076
rect 25136 11024 25188 11076
rect 31208 11092 31260 11144
rect 31484 11092 31536 11144
rect 31668 11135 31720 11144
rect 31668 11101 31677 11135
rect 31677 11101 31711 11135
rect 31711 11101 31720 11135
rect 31668 11092 31720 11101
rect 31576 11067 31628 11076
rect 31576 11033 31585 11067
rect 31585 11033 31619 11067
rect 31619 11033 31628 11067
rect 31576 11024 31628 11033
rect 20168 10956 20220 11008
rect 20260 10956 20312 11008
rect 25320 10956 25372 11008
rect 25964 10999 26016 11008
rect 25964 10965 25973 10999
rect 25973 10965 26007 10999
rect 26007 10965 26016 10999
rect 25964 10956 26016 10965
rect 28264 10956 28316 11008
rect 29276 10956 29328 11008
rect 31852 11135 31904 11144
rect 31852 11101 31861 11135
rect 31861 11101 31895 11135
rect 31895 11101 31904 11135
rect 31852 11092 31904 11101
rect 34336 11296 34388 11348
rect 32772 11228 32824 11280
rect 32588 11203 32640 11212
rect 32588 11169 32597 11203
rect 32597 11169 32631 11203
rect 32631 11169 32640 11203
rect 32588 11160 32640 11169
rect 32496 11092 32548 11144
rect 32312 11024 32364 11076
rect 33324 11135 33376 11144
rect 33324 11101 33333 11135
rect 33333 11101 33367 11135
rect 33367 11101 33376 11135
rect 33324 11092 33376 11101
rect 33140 11024 33192 11076
rect 33692 11160 33744 11212
rect 34336 11160 34388 11212
rect 35256 11203 35308 11212
rect 34244 11135 34296 11144
rect 34244 11101 34253 11135
rect 34253 11101 34287 11135
rect 34287 11101 34296 11135
rect 34244 11092 34296 11101
rect 35256 11169 35265 11203
rect 35265 11169 35299 11203
rect 35299 11169 35308 11203
rect 35256 11160 35308 11169
rect 36176 11160 36228 11212
rect 34520 11135 34572 11144
rect 34520 11101 34529 11135
rect 34529 11101 34563 11135
rect 34563 11101 34572 11135
rect 34520 11092 34572 11101
rect 34612 11092 34664 11144
rect 35072 11092 35124 11144
rect 33600 10956 33652 11008
rect 34704 10956 34756 11008
rect 36820 11024 36872 11076
rect 35900 10956 35952 11008
rect 36544 10956 36596 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 18052 10795 18104 10804
rect 18052 10761 18061 10795
rect 18061 10761 18095 10795
rect 18095 10761 18104 10795
rect 18052 10752 18104 10761
rect 17592 10684 17644 10736
rect 18236 10684 18288 10736
rect 18328 10727 18380 10736
rect 18328 10693 18337 10727
rect 18337 10693 18371 10727
rect 18371 10693 18380 10727
rect 18328 10684 18380 10693
rect 18420 10727 18472 10736
rect 18420 10693 18429 10727
rect 18429 10693 18463 10727
rect 18463 10693 18472 10727
rect 18420 10684 18472 10693
rect 18696 10684 18748 10736
rect 16488 10659 16540 10668
rect 16488 10625 16505 10659
rect 16505 10625 16539 10659
rect 16539 10625 16540 10659
rect 16488 10616 16540 10625
rect 17132 10616 17184 10668
rect 17684 10616 17736 10668
rect 19064 10752 19116 10804
rect 20720 10752 20772 10804
rect 22284 10752 22336 10804
rect 28356 10795 28408 10804
rect 28356 10761 28365 10795
rect 28365 10761 28399 10795
rect 28399 10761 28408 10795
rect 28356 10752 28408 10761
rect 32956 10795 33008 10804
rect 32956 10761 32965 10795
rect 32965 10761 32999 10795
rect 32999 10761 33008 10795
rect 32956 10752 33008 10761
rect 34520 10752 34572 10804
rect 17132 10480 17184 10532
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 17224 10455 17276 10464
rect 17224 10421 17233 10455
rect 17233 10421 17267 10455
rect 17267 10421 17276 10455
rect 17224 10412 17276 10421
rect 19340 10684 19392 10736
rect 22468 10727 22520 10736
rect 22468 10693 22477 10727
rect 22477 10693 22511 10727
rect 22511 10693 22520 10727
rect 22468 10684 22520 10693
rect 23664 10684 23716 10736
rect 26700 10684 26752 10736
rect 19156 10548 19208 10600
rect 19432 10616 19484 10668
rect 19984 10616 20036 10668
rect 22560 10616 22612 10668
rect 25320 10616 25372 10668
rect 25872 10659 25924 10668
rect 25872 10625 25881 10659
rect 25881 10625 25915 10659
rect 25915 10625 25924 10659
rect 25872 10616 25924 10625
rect 25964 10616 26016 10668
rect 26516 10616 26568 10668
rect 19432 10480 19484 10532
rect 24492 10548 24544 10600
rect 25504 10591 25556 10600
rect 25504 10557 25513 10591
rect 25513 10557 25547 10591
rect 25547 10557 25556 10591
rect 25504 10548 25556 10557
rect 26700 10548 26752 10600
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 28172 10684 28224 10736
rect 28264 10684 28316 10736
rect 28080 10659 28132 10668
rect 28080 10625 28089 10659
rect 28089 10625 28123 10659
rect 28123 10625 28132 10659
rect 28080 10616 28132 10625
rect 30472 10684 30524 10736
rect 31024 10684 31076 10736
rect 31484 10727 31536 10736
rect 31484 10693 31493 10727
rect 31493 10693 31527 10727
rect 31527 10693 31536 10727
rect 31484 10684 31536 10693
rect 32680 10684 32732 10736
rect 33416 10727 33468 10736
rect 33416 10693 33425 10727
rect 33425 10693 33459 10727
rect 33459 10693 33468 10727
rect 33416 10684 33468 10693
rect 34704 10684 34756 10736
rect 35164 10795 35216 10804
rect 35164 10761 35173 10795
rect 35173 10761 35207 10795
rect 35207 10761 35216 10795
rect 35164 10752 35216 10761
rect 35440 10752 35492 10804
rect 35900 10752 35952 10804
rect 36820 10795 36872 10804
rect 36820 10761 36829 10795
rect 36829 10761 36863 10795
rect 36863 10761 36872 10795
rect 36820 10752 36872 10761
rect 29000 10616 29052 10668
rect 36268 10616 36320 10668
rect 35992 10548 36044 10600
rect 36544 10591 36596 10600
rect 36544 10557 36553 10591
rect 36553 10557 36587 10591
rect 36587 10557 36596 10591
rect 36544 10548 36596 10557
rect 18972 10455 19024 10464
rect 18972 10421 18981 10455
rect 18981 10421 19015 10455
rect 19015 10421 19024 10455
rect 18972 10412 19024 10421
rect 20076 10455 20128 10464
rect 20076 10421 20085 10455
rect 20085 10421 20119 10455
rect 20119 10421 20128 10455
rect 20076 10412 20128 10421
rect 23020 10412 23072 10464
rect 32864 10480 32916 10532
rect 34428 10480 34480 10532
rect 24860 10455 24912 10464
rect 24860 10421 24869 10455
rect 24869 10421 24903 10455
rect 24903 10421 24912 10455
rect 24860 10412 24912 10421
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 25596 10412 25648 10421
rect 26332 10412 26384 10464
rect 26424 10455 26476 10464
rect 26424 10421 26433 10455
rect 26433 10421 26467 10455
rect 26467 10421 26476 10455
rect 26424 10412 26476 10421
rect 27804 10455 27856 10464
rect 27804 10421 27813 10455
rect 27813 10421 27847 10455
rect 27847 10421 27856 10455
rect 27804 10412 27856 10421
rect 34796 10412 34848 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 17224 10208 17276 10260
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 16396 10004 16448 10056
rect 16764 10004 16816 10056
rect 17500 10004 17552 10056
rect 17684 10004 17736 10056
rect 18696 10004 18748 10056
rect 20168 10208 20220 10260
rect 20812 10208 20864 10260
rect 23664 10251 23716 10260
rect 23664 10217 23673 10251
rect 23673 10217 23707 10251
rect 23707 10217 23716 10251
rect 23664 10208 23716 10217
rect 24492 10251 24544 10260
rect 24492 10217 24501 10251
rect 24501 10217 24535 10251
rect 24535 10217 24544 10251
rect 24492 10208 24544 10217
rect 24860 10208 24912 10260
rect 25228 10251 25280 10260
rect 25228 10217 25237 10251
rect 25237 10217 25271 10251
rect 25271 10217 25280 10251
rect 25228 10208 25280 10217
rect 25596 10208 25648 10260
rect 26516 10251 26568 10260
rect 26516 10217 26525 10251
rect 26525 10217 26559 10251
rect 26559 10217 26568 10251
rect 26516 10208 26568 10217
rect 30472 10251 30524 10260
rect 30472 10217 30481 10251
rect 30481 10217 30515 10251
rect 30515 10217 30524 10251
rect 30472 10208 30524 10217
rect 31392 10208 31444 10260
rect 32680 10208 32732 10260
rect 33784 10208 33836 10260
rect 34244 10208 34296 10260
rect 19340 10140 19392 10192
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 19984 10072 20036 10124
rect 20076 10072 20128 10124
rect 23020 10072 23072 10124
rect 25320 10004 25372 10056
rect 23848 9936 23900 9988
rect 17408 9911 17460 9920
rect 17408 9877 17417 9911
rect 17417 9877 17451 9911
rect 17451 9877 17460 9911
rect 17408 9868 17460 9877
rect 19340 9868 19392 9920
rect 24860 9979 24912 9988
rect 24860 9945 24869 9979
rect 24869 9945 24903 9979
rect 24903 9945 24912 9979
rect 24860 9936 24912 9945
rect 24952 9979 25004 9988
rect 24952 9945 24987 9979
rect 24987 9945 25004 9979
rect 24952 9936 25004 9945
rect 25136 9936 25188 9988
rect 25596 10047 25648 10056
rect 25596 10013 25605 10047
rect 25605 10013 25639 10047
rect 25639 10013 25648 10047
rect 25596 10004 25648 10013
rect 25688 10047 25740 10056
rect 25688 10013 25697 10047
rect 25697 10013 25731 10047
rect 25731 10013 25740 10047
rect 25688 10004 25740 10013
rect 25780 10004 25832 10056
rect 26056 10004 26108 10056
rect 31576 10115 31628 10124
rect 31576 10081 31585 10115
rect 31585 10081 31619 10115
rect 31619 10081 31628 10115
rect 31576 10072 31628 10081
rect 31944 10072 31996 10124
rect 33140 10140 33192 10192
rect 33416 10140 33468 10192
rect 26700 10047 26752 10056
rect 26700 10013 26709 10047
rect 26709 10013 26743 10047
rect 26743 10013 26752 10047
rect 26700 10004 26752 10013
rect 29276 10004 29328 10056
rect 30288 10004 30340 10056
rect 31116 10004 31168 10056
rect 32404 10072 32456 10124
rect 33324 10072 33376 10124
rect 35256 10115 35308 10124
rect 35256 10081 35265 10115
rect 35265 10081 35299 10115
rect 35299 10081 35308 10115
rect 35256 10072 35308 10081
rect 32864 10047 32916 10056
rect 32864 10013 32873 10047
rect 32873 10013 32907 10047
rect 32907 10013 32916 10047
rect 32864 10004 32916 10013
rect 33140 10047 33192 10056
rect 33140 10013 33149 10047
rect 33149 10013 33183 10047
rect 33183 10013 33192 10047
rect 33140 10004 33192 10013
rect 33692 10047 33744 10056
rect 33692 10013 33701 10047
rect 33701 10013 33735 10047
rect 33735 10013 33744 10047
rect 33692 10004 33744 10013
rect 34796 10004 34848 10056
rect 25504 9936 25556 9988
rect 68468 10047 68520 10056
rect 68468 10013 68477 10047
rect 68477 10013 68511 10047
rect 68511 10013 68520 10047
rect 68468 10004 68520 10013
rect 26332 9911 26384 9920
rect 26332 9877 26341 9911
rect 26341 9877 26375 9911
rect 26375 9877 26384 9911
rect 26332 9868 26384 9877
rect 28816 9868 28868 9920
rect 30932 9911 30984 9920
rect 30932 9877 30941 9911
rect 30941 9877 30975 9911
rect 30975 9877 30984 9911
rect 30932 9868 30984 9877
rect 32588 9911 32640 9920
rect 32588 9877 32597 9911
rect 32597 9877 32631 9911
rect 32631 9877 32640 9911
rect 32588 9868 32640 9877
rect 33416 9911 33468 9920
rect 33416 9877 33425 9911
rect 33425 9877 33459 9911
rect 33459 9877 33468 9911
rect 33416 9868 33468 9877
rect 34704 9911 34756 9920
rect 34704 9877 34713 9911
rect 34713 9877 34747 9911
rect 34747 9877 34756 9911
rect 34704 9868 34756 9877
rect 35532 9911 35584 9920
rect 35532 9877 35541 9911
rect 35541 9877 35575 9911
rect 35575 9877 35584 9911
rect 35532 9868 35584 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 17132 9664 17184 9716
rect 17500 9664 17552 9716
rect 15936 9596 15988 9648
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 16764 9460 16816 9512
rect 16948 9571 17000 9580
rect 16948 9537 16957 9571
rect 16957 9537 16991 9571
rect 16991 9537 17000 9571
rect 16948 9528 17000 9537
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 17132 9571 17184 9580
rect 17132 9537 17167 9571
rect 17167 9537 17184 9571
rect 17132 9528 17184 9537
rect 17408 9528 17460 9580
rect 15568 9324 15620 9376
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 18144 9639 18196 9648
rect 18144 9605 18153 9639
rect 18153 9605 18187 9639
rect 18187 9605 18196 9639
rect 18144 9596 18196 9605
rect 18880 9639 18932 9648
rect 17960 9528 18012 9580
rect 18880 9605 18891 9639
rect 18891 9605 18932 9639
rect 18880 9596 18932 9605
rect 23020 9707 23072 9716
rect 23020 9673 23029 9707
rect 23029 9673 23063 9707
rect 23063 9673 23072 9707
rect 23020 9664 23072 9673
rect 24952 9664 25004 9716
rect 25228 9664 25280 9716
rect 25688 9664 25740 9716
rect 26700 9664 26752 9716
rect 27804 9664 27856 9716
rect 19432 9596 19484 9648
rect 20260 9596 20312 9648
rect 21272 9639 21324 9648
rect 21272 9605 21281 9639
rect 21281 9605 21315 9639
rect 21315 9605 21324 9639
rect 21272 9596 21324 9605
rect 26240 9596 26292 9648
rect 26424 9596 26476 9648
rect 28816 9596 28868 9648
rect 31116 9664 31168 9716
rect 18972 9528 19024 9580
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 17684 9503 17736 9512
rect 17684 9469 17693 9503
rect 17693 9469 17727 9503
rect 17727 9469 17736 9503
rect 17684 9460 17736 9469
rect 18604 9503 18656 9512
rect 18604 9469 18619 9503
rect 18619 9469 18653 9503
rect 18653 9469 18656 9503
rect 18604 9460 18656 9469
rect 18512 9435 18564 9444
rect 18512 9401 18521 9435
rect 18521 9401 18555 9435
rect 18555 9401 18564 9435
rect 18512 9392 18564 9401
rect 21088 9460 21140 9512
rect 21548 9571 21600 9580
rect 21548 9537 21557 9571
rect 21557 9537 21591 9571
rect 21591 9537 21600 9571
rect 21548 9528 21600 9537
rect 21916 9460 21968 9512
rect 20904 9392 20956 9444
rect 24768 9571 24820 9580
rect 24768 9537 24777 9571
rect 24777 9537 24811 9571
rect 24811 9537 24820 9571
rect 24768 9528 24820 9537
rect 24952 9571 25004 9580
rect 24952 9537 24961 9571
rect 24961 9537 24995 9571
rect 24995 9537 25004 9571
rect 24952 9528 25004 9537
rect 25780 9528 25832 9580
rect 25872 9528 25924 9580
rect 27160 9528 27212 9580
rect 31208 9596 31260 9648
rect 31944 9639 31996 9648
rect 31944 9605 31953 9639
rect 31953 9605 31987 9639
rect 31987 9605 31996 9639
rect 31944 9596 31996 9605
rect 29552 9571 29604 9580
rect 29552 9537 29561 9571
rect 29561 9537 29595 9571
rect 29595 9537 29604 9571
rect 29552 9528 29604 9537
rect 24400 9503 24452 9512
rect 24400 9469 24409 9503
rect 24409 9469 24443 9503
rect 24443 9469 24452 9503
rect 24400 9460 24452 9469
rect 25964 9460 26016 9512
rect 26424 9503 26476 9512
rect 26424 9469 26433 9503
rect 26433 9469 26467 9503
rect 26467 9469 26476 9503
rect 26424 9460 26476 9469
rect 18604 9324 18656 9376
rect 19340 9324 19392 9376
rect 20720 9367 20772 9376
rect 20720 9333 20729 9367
rect 20729 9333 20763 9367
rect 20763 9333 20772 9367
rect 20720 9324 20772 9333
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 20996 9324 21048 9333
rect 22284 9324 22336 9376
rect 23112 9367 23164 9376
rect 23112 9333 23121 9367
rect 23121 9333 23155 9367
rect 23155 9333 23164 9367
rect 23112 9324 23164 9333
rect 24676 9324 24728 9376
rect 25044 9367 25096 9376
rect 25044 9333 25053 9367
rect 25053 9333 25087 9367
rect 25087 9333 25096 9367
rect 25044 9324 25096 9333
rect 26332 9367 26384 9376
rect 26332 9333 26341 9367
rect 26341 9333 26375 9367
rect 26375 9333 26384 9367
rect 26332 9324 26384 9333
rect 26516 9324 26568 9376
rect 27436 9324 27488 9376
rect 27804 9503 27856 9512
rect 27804 9469 27813 9503
rect 27813 9469 27847 9503
rect 27847 9469 27856 9503
rect 27804 9460 27856 9469
rect 29000 9460 29052 9512
rect 30748 9460 30800 9512
rect 32404 9664 32456 9716
rect 32588 9664 32640 9716
rect 32864 9664 32916 9716
rect 32680 9639 32732 9648
rect 32680 9605 32715 9639
rect 32715 9605 32732 9639
rect 32680 9596 32732 9605
rect 32588 9571 32640 9580
rect 32588 9537 32597 9571
rect 32597 9537 32631 9571
rect 32631 9537 32640 9571
rect 32588 9528 32640 9537
rect 33416 9664 33468 9716
rect 35256 9664 35308 9716
rect 33600 9639 33652 9648
rect 33600 9605 33622 9639
rect 33622 9605 33652 9639
rect 33600 9596 33652 9605
rect 34244 9639 34296 9648
rect 34244 9605 34253 9639
rect 34253 9605 34287 9639
rect 34287 9605 34296 9639
rect 34244 9596 34296 9605
rect 29736 9367 29788 9376
rect 29736 9333 29745 9367
rect 29745 9333 29779 9367
rect 29779 9333 29788 9367
rect 29736 9324 29788 9333
rect 29828 9324 29880 9376
rect 32220 9367 32272 9376
rect 32220 9333 32229 9367
rect 32229 9333 32263 9367
rect 32263 9333 32272 9367
rect 32220 9324 32272 9333
rect 33416 9324 33468 9376
rect 33968 9571 34020 9580
rect 33968 9537 33977 9571
rect 33977 9537 34011 9571
rect 34011 9537 34020 9571
rect 33968 9528 34020 9537
rect 35992 9571 36044 9580
rect 35992 9537 36001 9571
rect 36001 9537 36035 9571
rect 36035 9537 36044 9571
rect 35992 9528 36044 9537
rect 34704 9460 34756 9512
rect 33784 9392 33836 9444
rect 35532 9324 35584 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 15936 9163 15988 9172
rect 15936 9129 15945 9163
rect 15945 9129 15979 9163
rect 15979 9129 15988 9163
rect 15936 9120 15988 9129
rect 16948 9120 17000 9172
rect 20076 9120 20128 9172
rect 20536 9120 20588 9172
rect 20996 9120 21048 9172
rect 17960 9052 18012 9104
rect 18328 9052 18380 9104
rect 19064 9052 19116 9104
rect 17684 8984 17736 9036
rect 18972 8984 19024 9036
rect 19248 8984 19300 9036
rect 16488 8916 16540 8968
rect 16764 8916 16816 8968
rect 17592 8916 17644 8968
rect 22468 9120 22520 9172
rect 24400 9120 24452 9172
rect 24768 9120 24820 9172
rect 25596 9120 25648 9172
rect 25872 9120 25924 9172
rect 26424 9163 26476 9172
rect 26424 9129 26433 9163
rect 26433 9129 26467 9163
rect 26467 9129 26476 9163
rect 26424 9120 26476 9129
rect 26516 9120 26568 9172
rect 22284 9095 22336 9104
rect 22284 9061 22293 9095
rect 22293 9061 22327 9095
rect 22327 9061 22336 9095
rect 22284 9052 22336 9061
rect 22008 8984 22060 9036
rect 23112 8984 23164 9036
rect 25320 9027 25372 9036
rect 25320 8993 25329 9027
rect 25329 8993 25363 9027
rect 25363 8993 25372 9027
rect 25320 8984 25372 8993
rect 17132 8780 17184 8832
rect 18696 8780 18748 8832
rect 19340 8780 19392 8832
rect 19984 8780 20036 8832
rect 20904 8848 20956 8900
rect 22652 8848 22704 8900
rect 23664 8848 23716 8900
rect 25964 8916 26016 8968
rect 26516 8916 26568 8968
rect 27160 9120 27212 9172
rect 27804 9163 27856 9172
rect 27804 9129 27813 9163
rect 27813 9129 27847 9163
rect 27847 9129 27856 9163
rect 27804 9120 27856 9129
rect 29736 9120 29788 9172
rect 31208 9120 31260 9172
rect 29552 9052 29604 9104
rect 29644 9052 29696 9104
rect 27344 8891 27396 8900
rect 27344 8857 27353 8891
rect 27353 8857 27387 8891
rect 27387 8857 27396 8891
rect 27344 8848 27396 8857
rect 27528 8891 27580 8900
rect 27528 8857 27569 8891
rect 27569 8857 27580 8891
rect 27528 8848 27580 8857
rect 28908 8891 28960 8900
rect 28908 8857 28917 8891
rect 28917 8857 28951 8891
rect 28951 8857 28960 8891
rect 28908 8848 28960 8857
rect 29276 8848 29328 8900
rect 29828 8984 29880 9036
rect 33876 9120 33928 9172
rect 34796 9120 34848 9172
rect 33508 9052 33560 9104
rect 34612 9052 34664 9104
rect 32220 8984 32272 9036
rect 33324 9027 33376 9036
rect 33324 8993 33333 9027
rect 33333 8993 33367 9027
rect 33367 8993 33376 9027
rect 33324 8984 33376 8993
rect 30656 8916 30708 8968
rect 33692 8959 33744 8968
rect 33692 8925 33701 8959
rect 33701 8925 33735 8959
rect 33735 8925 33744 8959
rect 33692 8916 33744 8925
rect 32036 8848 32088 8900
rect 33232 8848 33284 8900
rect 21548 8780 21600 8832
rect 27252 8780 27304 8832
rect 28264 8780 28316 8832
rect 28540 8780 28592 8832
rect 31208 8780 31260 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 18696 8619 18748 8628
rect 17040 8576 17092 8585
rect 18696 8585 18705 8619
rect 18705 8585 18739 8619
rect 18739 8585 18748 8619
rect 18696 8576 18748 8585
rect 19064 8576 19116 8628
rect 19984 8576 20036 8628
rect 20076 8576 20128 8628
rect 17132 8551 17184 8560
rect 17132 8517 17141 8551
rect 17141 8517 17175 8551
rect 17175 8517 17184 8551
rect 17132 8508 17184 8517
rect 18328 8483 18380 8492
rect 18328 8449 18337 8483
rect 18337 8449 18371 8483
rect 18371 8449 18380 8483
rect 18328 8440 18380 8449
rect 19156 8508 19208 8560
rect 17592 8372 17644 8424
rect 18512 8347 18564 8356
rect 18512 8313 18521 8347
rect 18521 8313 18555 8347
rect 18555 8313 18564 8347
rect 18512 8304 18564 8313
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 19064 8440 19116 8492
rect 20812 8576 20864 8628
rect 21088 8576 21140 8628
rect 21272 8576 21324 8628
rect 22652 8619 22704 8628
rect 22652 8585 22661 8619
rect 22661 8585 22695 8619
rect 22695 8585 22704 8619
rect 22652 8576 22704 8585
rect 23664 8576 23716 8628
rect 23848 8576 23900 8628
rect 25044 8576 25096 8628
rect 30656 8619 30708 8628
rect 20720 8508 20772 8560
rect 21916 8440 21968 8492
rect 22744 8483 22796 8492
rect 22744 8449 22753 8483
rect 22753 8449 22787 8483
rect 22787 8449 22796 8483
rect 22744 8440 22796 8449
rect 24952 8508 25004 8560
rect 25320 8440 25372 8492
rect 27252 8508 27304 8560
rect 30656 8585 30665 8619
rect 30665 8585 30699 8619
rect 30699 8585 30708 8619
rect 30656 8576 30708 8585
rect 30748 8619 30800 8628
rect 30748 8585 30757 8619
rect 30757 8585 30791 8619
rect 30791 8585 30800 8619
rect 30748 8576 30800 8585
rect 30932 8576 30984 8628
rect 32036 8576 32088 8628
rect 24124 8372 24176 8424
rect 24676 8415 24728 8424
rect 24676 8381 24685 8415
rect 24685 8381 24719 8415
rect 24719 8381 24728 8415
rect 24676 8372 24728 8381
rect 19248 8304 19300 8356
rect 19616 8304 19668 8356
rect 20536 8304 20588 8356
rect 24952 8415 25004 8424
rect 24952 8381 24961 8415
rect 24961 8381 24995 8415
rect 24995 8381 25004 8415
rect 24952 8372 25004 8381
rect 27160 8372 27212 8424
rect 28172 8483 28224 8492
rect 28172 8449 28181 8483
rect 28181 8449 28215 8483
rect 28215 8449 28224 8483
rect 28172 8440 28224 8449
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 28540 8483 28592 8492
rect 28540 8449 28549 8483
rect 28549 8449 28583 8483
rect 28583 8449 28592 8483
rect 28540 8440 28592 8449
rect 29276 8508 29328 8560
rect 30196 8508 30248 8560
rect 28816 8440 28868 8492
rect 28908 8483 28960 8492
rect 28908 8449 28917 8483
rect 28917 8449 28951 8483
rect 28951 8449 28960 8483
rect 28908 8440 28960 8449
rect 25872 8304 25924 8356
rect 28264 8304 28316 8356
rect 16672 8279 16724 8288
rect 16672 8245 16681 8279
rect 16681 8245 16715 8279
rect 16715 8245 16724 8279
rect 16672 8236 16724 8245
rect 19064 8279 19116 8288
rect 19064 8245 19073 8279
rect 19073 8245 19107 8279
rect 19107 8245 19116 8279
rect 19064 8236 19116 8245
rect 19156 8279 19208 8288
rect 19156 8245 19165 8279
rect 19165 8245 19199 8279
rect 19199 8245 19208 8279
rect 19156 8236 19208 8245
rect 19340 8279 19392 8288
rect 19340 8245 19349 8279
rect 19349 8245 19383 8279
rect 19383 8245 19392 8279
rect 19340 8236 19392 8245
rect 20168 8279 20220 8288
rect 20168 8245 20177 8279
rect 20177 8245 20211 8279
rect 20211 8245 20220 8279
rect 20168 8236 20220 8245
rect 25136 8279 25188 8288
rect 25136 8245 25145 8279
rect 25145 8245 25179 8279
rect 25179 8245 25188 8279
rect 25136 8236 25188 8245
rect 25228 8279 25280 8288
rect 25228 8245 25237 8279
rect 25237 8245 25271 8279
rect 25271 8245 25280 8279
rect 25228 8236 25280 8245
rect 25964 8279 26016 8288
rect 25964 8245 25973 8279
rect 25973 8245 26007 8279
rect 26007 8245 26016 8279
rect 25964 8236 26016 8245
rect 27344 8279 27396 8288
rect 27344 8245 27353 8279
rect 27353 8245 27387 8279
rect 27387 8245 27396 8279
rect 27344 8236 27396 8245
rect 31208 8372 31260 8424
rect 29184 8236 29236 8288
rect 30288 8236 30340 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 17592 8032 17644 8084
rect 18512 8032 18564 8084
rect 19248 8032 19300 8084
rect 28172 8032 28224 8084
rect 29552 8032 29604 8084
rect 30196 8075 30248 8084
rect 30196 8041 30205 8075
rect 30205 8041 30239 8075
rect 30239 8041 30248 8075
rect 30196 8032 30248 8041
rect 24768 7964 24820 8016
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 15844 7896 15896 7948
rect 19064 7896 19116 7948
rect 20076 7896 20128 7948
rect 15936 7760 15988 7812
rect 16856 7760 16908 7812
rect 18972 7871 19024 7880
rect 18972 7837 18981 7871
rect 18981 7837 19015 7871
rect 19015 7837 19024 7871
rect 18972 7828 19024 7837
rect 19156 7828 19208 7880
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 21824 7828 21876 7880
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 24124 7828 24176 7880
rect 25136 7828 25188 7880
rect 26056 7871 26108 7880
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 26148 7828 26200 7880
rect 26608 7828 26660 7880
rect 27528 7828 27580 7880
rect 27896 7828 27948 7880
rect 29184 7871 29236 7880
rect 29184 7837 29193 7871
rect 29193 7837 29227 7871
rect 29227 7837 29236 7871
rect 29184 7828 29236 7837
rect 30288 7871 30340 7880
rect 30288 7837 30297 7871
rect 30297 7837 30331 7871
rect 30331 7837 30340 7871
rect 30288 7828 30340 7837
rect 17868 7735 17920 7744
rect 17868 7701 17877 7735
rect 17877 7701 17911 7735
rect 17911 7701 17920 7735
rect 17868 7692 17920 7701
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 21180 7735 21232 7744
rect 21180 7701 21189 7735
rect 21189 7701 21223 7735
rect 21223 7701 21232 7735
rect 21180 7692 21232 7701
rect 22836 7735 22888 7744
rect 22836 7701 22845 7735
rect 22845 7701 22879 7735
rect 22879 7701 22888 7735
rect 22836 7692 22888 7701
rect 23664 7692 23716 7744
rect 25596 7760 25648 7812
rect 29736 7760 29788 7812
rect 27804 7692 27856 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 15936 7488 15988 7540
rect 16672 7488 16724 7540
rect 16856 7488 16908 7540
rect 17868 7488 17920 7540
rect 18972 7488 19024 7540
rect 19248 7488 19300 7540
rect 18328 7420 18380 7472
rect 16764 7352 16816 7404
rect 19800 7352 19852 7404
rect 22008 7488 22060 7540
rect 20168 7463 20220 7472
rect 20168 7429 20177 7463
rect 20177 7429 20211 7463
rect 20211 7429 20220 7463
rect 20168 7420 20220 7429
rect 21180 7420 21232 7472
rect 23664 7488 23716 7540
rect 24124 7488 24176 7540
rect 22192 7420 22244 7472
rect 22836 7420 22888 7472
rect 15844 7284 15896 7336
rect 24768 7463 24820 7472
rect 24768 7429 24777 7463
rect 24777 7429 24811 7463
rect 24811 7429 24820 7463
rect 24768 7420 24820 7429
rect 26056 7488 26108 7540
rect 25964 7463 26016 7472
rect 24952 7352 25004 7404
rect 25228 7352 25280 7404
rect 21916 7216 21968 7268
rect 24124 7216 24176 7268
rect 24216 7216 24268 7268
rect 25964 7429 25973 7463
rect 25973 7429 26007 7463
rect 26007 7429 26016 7463
rect 25964 7420 26016 7429
rect 19524 7191 19576 7200
rect 19524 7157 19533 7191
rect 19533 7157 19567 7191
rect 19567 7157 19576 7191
rect 19524 7148 19576 7157
rect 24400 7191 24452 7200
rect 24400 7157 24409 7191
rect 24409 7157 24443 7191
rect 24443 7157 24452 7191
rect 24400 7148 24452 7157
rect 25872 7352 25924 7404
rect 27160 7488 27212 7540
rect 27528 7488 27580 7540
rect 27804 7420 27856 7472
rect 28080 7420 28132 7472
rect 26516 7284 26568 7336
rect 27344 7395 27396 7404
rect 27344 7361 27353 7395
rect 27353 7361 27387 7395
rect 27387 7361 27396 7395
rect 27344 7352 27396 7361
rect 27896 7352 27948 7404
rect 27068 7327 27120 7336
rect 27068 7293 27077 7327
rect 27077 7293 27111 7327
rect 27111 7293 27120 7327
rect 27068 7284 27120 7293
rect 27804 7327 27856 7336
rect 27804 7293 27813 7327
rect 27813 7293 27847 7327
rect 27847 7293 27856 7327
rect 27804 7284 27856 7293
rect 27988 7216 28040 7268
rect 28172 7148 28224 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 16764 6944 16816 6996
rect 18328 6944 18380 6996
rect 19524 6944 19576 6996
rect 24400 6944 24452 6996
rect 27344 6987 27396 6996
rect 27344 6953 27353 6987
rect 27353 6953 27387 6987
rect 27387 6953 27396 6987
rect 27344 6944 27396 6953
rect 20076 6808 20128 6860
rect 22192 6851 22244 6860
rect 22192 6817 22201 6851
rect 22201 6817 22235 6851
rect 22235 6817 22244 6851
rect 22192 6808 22244 6817
rect 24216 6851 24268 6860
rect 24216 6817 24225 6851
rect 24225 6817 24259 6851
rect 24259 6817 24268 6851
rect 24216 6808 24268 6817
rect 27436 6851 27488 6860
rect 27436 6817 27445 6851
rect 27445 6817 27479 6851
rect 27479 6817 27488 6851
rect 27436 6808 27488 6817
rect 28816 6876 28868 6928
rect 28264 6808 28316 6860
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 21824 6783 21876 6792
rect 21824 6749 21833 6783
rect 21833 6749 21867 6783
rect 21867 6749 21876 6783
rect 21824 6740 21876 6749
rect 23572 6740 23624 6792
rect 26056 6672 26108 6724
rect 26516 6672 26568 6724
rect 26608 6672 26660 6724
rect 27160 6783 27212 6792
rect 27160 6749 27169 6783
rect 27169 6749 27203 6783
rect 27203 6749 27212 6783
rect 27160 6740 27212 6749
rect 29736 6783 29788 6792
rect 29736 6749 29745 6783
rect 29745 6749 29779 6783
rect 29779 6749 29788 6783
rect 29736 6740 29788 6749
rect 27712 6715 27764 6724
rect 27712 6681 27721 6715
rect 27721 6681 27755 6715
rect 27755 6681 27764 6715
rect 27712 6672 27764 6681
rect 29460 6604 29512 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 23572 6443 23624 6452
rect 23572 6409 23581 6443
rect 23581 6409 23615 6443
rect 23615 6409 23624 6443
rect 23572 6400 23624 6409
rect 23848 6400 23900 6452
rect 26056 6400 26108 6452
rect 27712 6400 27764 6452
rect 27804 6332 27856 6384
rect 27988 6375 28040 6384
rect 27988 6341 27997 6375
rect 27997 6341 28031 6375
rect 28031 6341 28040 6375
rect 27988 6332 28040 6341
rect 28172 6332 28224 6384
rect 26516 6264 26568 6316
rect 28080 6307 28132 6316
rect 28080 6273 28089 6307
rect 28089 6273 28123 6307
rect 28123 6273 28132 6307
rect 28080 6264 28132 6273
rect 29460 6196 29512 6248
rect 28264 6171 28316 6180
rect 28264 6137 28273 6171
rect 28273 6137 28307 6171
rect 28307 6137 28316 6171
rect 28264 6128 28316 6137
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 8392 3476 8444 3528
rect 13728 3476 13780 3528
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 20352 3000 20404 3052
rect 43260 2839 43312 2848
rect 43260 2805 43269 2839
rect 43269 2805 43303 2839
rect 43303 2805 43312 2839
rect 43260 2796 43312 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 26516 2431 26568 2440
rect 26516 2397 26525 2431
rect 26525 2397 26559 2431
rect 26559 2397 26568 2431
rect 26516 2388 26568 2397
rect 43260 2388 43312 2440
rect 67640 2431 67692 2440
rect 67640 2397 67649 2431
rect 67649 2397 67683 2431
rect 67683 2397 67692 2431
rect 67640 2388 67692 2397
rect 43812 2252 43864 2304
rect 68008 2252 68060 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 3882 69200 3938 70000
rect 12898 69306 12954 70000
rect 12898 69278 13032 69306
rect 12898 69200 12954 69278
rect 13004 67250 13032 69278
rect 21270 69200 21326 70000
rect 30286 69200 30342 70000
rect 39302 69306 39358 70000
rect 39302 69278 39436 69306
rect 39302 69200 39358 69278
rect 30300 67538 30328 69200
rect 30300 67510 30420 67538
rect 19574 67484 19882 67493
rect 19574 67482 19580 67484
rect 19636 67482 19660 67484
rect 19716 67482 19740 67484
rect 19796 67482 19820 67484
rect 19876 67482 19882 67484
rect 19636 67430 19638 67482
rect 19818 67430 19820 67482
rect 19574 67428 19580 67430
rect 19636 67428 19660 67430
rect 19716 67428 19740 67430
rect 19796 67428 19820 67430
rect 19876 67428 19882 67430
rect 19574 67419 19882 67428
rect 30392 67250 30420 67510
rect 39408 67250 39436 69278
rect 47674 69200 47730 70000
rect 56690 69200 56746 70000
rect 65706 69200 65762 70000
rect 50294 67484 50602 67493
rect 50294 67482 50300 67484
rect 50356 67482 50380 67484
rect 50436 67482 50460 67484
rect 50516 67482 50540 67484
rect 50596 67482 50602 67484
rect 50356 67430 50358 67482
rect 50538 67430 50540 67482
rect 50294 67428 50300 67430
rect 50356 67428 50380 67430
rect 50436 67428 50460 67430
rect 50516 67428 50540 67430
rect 50596 67428 50602 67430
rect 50294 67419 50602 67428
rect 12992 67244 13044 67250
rect 12992 67186 13044 67192
rect 30380 67244 30432 67250
rect 30380 67186 30432 67192
rect 39396 67244 39448 67250
rect 39396 67186 39448 67192
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 19574 66396 19882 66405
rect 19574 66394 19580 66396
rect 19636 66394 19660 66396
rect 19716 66394 19740 66396
rect 19796 66394 19820 66396
rect 19876 66394 19882 66396
rect 19636 66342 19638 66394
rect 19818 66342 19820 66394
rect 19574 66340 19580 66342
rect 19636 66340 19660 66342
rect 19716 66340 19740 66342
rect 19796 66340 19820 66342
rect 19876 66340 19882 66342
rect 19574 66331 19882 66340
rect 50294 66396 50602 66405
rect 50294 66394 50300 66396
rect 50356 66394 50380 66396
rect 50436 66394 50460 66396
rect 50516 66394 50540 66396
rect 50596 66394 50602 66396
rect 50356 66342 50358 66394
rect 50538 66342 50540 66394
rect 50294 66340 50300 66342
rect 50356 66340 50380 66342
rect 50436 66340 50460 66342
rect 50516 66340 50540 66342
rect 50596 66340 50602 66342
rect 50294 66331 50602 66340
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 19574 65308 19882 65317
rect 19574 65306 19580 65308
rect 19636 65306 19660 65308
rect 19716 65306 19740 65308
rect 19796 65306 19820 65308
rect 19876 65306 19882 65308
rect 19636 65254 19638 65306
rect 19818 65254 19820 65306
rect 19574 65252 19580 65254
rect 19636 65252 19660 65254
rect 19716 65252 19740 65254
rect 19796 65252 19820 65254
rect 19876 65252 19882 65254
rect 19574 65243 19882 65252
rect 50294 65308 50602 65317
rect 50294 65306 50300 65308
rect 50356 65306 50380 65308
rect 50436 65306 50460 65308
rect 50516 65306 50540 65308
rect 50596 65306 50602 65308
rect 50356 65254 50358 65306
rect 50538 65254 50540 65306
rect 50294 65252 50300 65254
rect 50356 65252 50380 65254
rect 50436 65252 50460 65254
rect 50516 65252 50540 65254
rect 50596 65252 50602 65254
rect 50294 65243 50602 65252
rect 1400 65000 1452 65006
rect 1400 64942 1452 64948
rect 1412 64841 1440 64942
rect 1398 64832 1454 64841
rect 1398 64767 1454 64776
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 34934 64764 35242 64773
rect 34934 64762 34940 64764
rect 34996 64762 35020 64764
rect 35076 64762 35100 64764
rect 35156 64762 35180 64764
rect 35236 64762 35242 64764
rect 34996 64710 34998 64762
rect 35178 64710 35180 64762
rect 34934 64708 34940 64710
rect 34996 64708 35020 64710
rect 35076 64708 35100 64710
rect 35156 64708 35180 64710
rect 35236 64708 35242 64710
rect 34934 64699 35242 64708
rect 65654 64764 65962 64773
rect 65654 64762 65660 64764
rect 65716 64762 65740 64764
rect 65796 64762 65820 64764
rect 65876 64762 65900 64764
rect 65956 64762 65962 64764
rect 65716 64710 65718 64762
rect 65898 64710 65900 64762
rect 65654 64708 65660 64710
rect 65716 64708 65740 64710
rect 65796 64708 65820 64710
rect 65876 64708 65900 64710
rect 65956 64708 65962 64710
rect 65654 64699 65962 64708
rect 19574 64220 19882 64229
rect 19574 64218 19580 64220
rect 19636 64218 19660 64220
rect 19716 64218 19740 64220
rect 19796 64218 19820 64220
rect 19876 64218 19882 64220
rect 19636 64166 19638 64218
rect 19818 64166 19820 64218
rect 19574 64164 19580 64166
rect 19636 64164 19660 64166
rect 19716 64164 19740 64166
rect 19796 64164 19820 64166
rect 19876 64164 19882 64166
rect 19574 64155 19882 64164
rect 50294 64220 50602 64229
rect 50294 64218 50300 64220
rect 50356 64218 50380 64220
rect 50436 64218 50460 64220
rect 50516 64218 50540 64220
rect 50596 64218 50602 64220
rect 50356 64166 50358 64218
rect 50538 64166 50540 64218
rect 50294 64164 50300 64166
rect 50356 64164 50380 64166
rect 50436 64164 50460 64166
rect 50516 64164 50540 64166
rect 50596 64164 50602 64166
rect 50294 64155 50602 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 34934 63676 35242 63685
rect 34934 63674 34940 63676
rect 34996 63674 35020 63676
rect 35076 63674 35100 63676
rect 35156 63674 35180 63676
rect 35236 63674 35242 63676
rect 34996 63622 34998 63674
rect 35178 63622 35180 63674
rect 34934 63620 34940 63622
rect 34996 63620 35020 63622
rect 35076 63620 35100 63622
rect 35156 63620 35180 63622
rect 35236 63620 35242 63622
rect 34934 63611 35242 63620
rect 65654 63676 65962 63685
rect 65654 63674 65660 63676
rect 65716 63674 65740 63676
rect 65796 63674 65820 63676
rect 65876 63674 65900 63676
rect 65956 63674 65962 63676
rect 65716 63622 65718 63674
rect 65898 63622 65900 63674
rect 65654 63620 65660 63622
rect 65716 63620 65740 63622
rect 65796 63620 65820 63622
rect 65876 63620 65900 63622
rect 65956 63620 65962 63622
rect 65654 63611 65962 63620
rect 19574 63132 19882 63141
rect 19574 63130 19580 63132
rect 19636 63130 19660 63132
rect 19716 63130 19740 63132
rect 19796 63130 19820 63132
rect 19876 63130 19882 63132
rect 19636 63078 19638 63130
rect 19818 63078 19820 63130
rect 19574 63076 19580 63078
rect 19636 63076 19660 63078
rect 19716 63076 19740 63078
rect 19796 63076 19820 63078
rect 19876 63076 19882 63078
rect 19574 63067 19882 63076
rect 50294 63132 50602 63141
rect 50294 63130 50300 63132
rect 50356 63130 50380 63132
rect 50436 63130 50460 63132
rect 50516 63130 50540 63132
rect 50596 63130 50602 63132
rect 50356 63078 50358 63130
rect 50538 63078 50540 63130
rect 50294 63076 50300 63078
rect 50356 63076 50380 63078
rect 50436 63076 50460 63078
rect 50516 63076 50540 63078
rect 50596 63076 50602 63078
rect 50294 63067 50602 63076
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 34934 62588 35242 62597
rect 34934 62586 34940 62588
rect 34996 62586 35020 62588
rect 35076 62586 35100 62588
rect 35156 62586 35180 62588
rect 35236 62586 35242 62588
rect 34996 62534 34998 62586
rect 35178 62534 35180 62586
rect 34934 62532 34940 62534
rect 34996 62532 35020 62534
rect 35076 62532 35100 62534
rect 35156 62532 35180 62534
rect 35236 62532 35242 62534
rect 34934 62523 35242 62532
rect 65654 62588 65962 62597
rect 65654 62586 65660 62588
rect 65716 62586 65740 62588
rect 65796 62586 65820 62588
rect 65876 62586 65900 62588
rect 65956 62586 65962 62588
rect 65716 62534 65718 62586
rect 65898 62534 65900 62586
rect 65654 62532 65660 62534
rect 65716 62532 65740 62534
rect 65796 62532 65820 62534
rect 65876 62532 65900 62534
rect 65956 62532 65962 62534
rect 65654 62523 65962 62532
rect 19574 62044 19882 62053
rect 19574 62042 19580 62044
rect 19636 62042 19660 62044
rect 19716 62042 19740 62044
rect 19796 62042 19820 62044
rect 19876 62042 19882 62044
rect 19636 61990 19638 62042
rect 19818 61990 19820 62042
rect 19574 61988 19580 61990
rect 19636 61988 19660 61990
rect 19716 61988 19740 61990
rect 19796 61988 19820 61990
rect 19876 61988 19882 61990
rect 19574 61979 19882 61988
rect 50294 62044 50602 62053
rect 50294 62042 50300 62044
rect 50356 62042 50380 62044
rect 50436 62042 50460 62044
rect 50516 62042 50540 62044
rect 50596 62042 50602 62044
rect 50356 61990 50358 62042
rect 50538 61990 50540 62042
rect 50294 61988 50300 61990
rect 50356 61988 50380 61990
rect 50436 61988 50460 61990
rect 50516 61988 50540 61990
rect 50596 61988 50602 61990
rect 50294 61979 50602 61988
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 65654 61500 65962 61509
rect 65654 61498 65660 61500
rect 65716 61498 65740 61500
rect 65796 61498 65820 61500
rect 65876 61498 65900 61500
rect 65956 61498 65962 61500
rect 65716 61446 65718 61498
rect 65898 61446 65900 61498
rect 65654 61444 65660 61446
rect 65716 61444 65740 61446
rect 65796 61444 65820 61446
rect 65876 61444 65900 61446
rect 65956 61444 65962 61446
rect 65654 61435 65962 61444
rect 19574 60956 19882 60965
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60891 19882 60900
rect 50294 60956 50602 60965
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60891 50602 60900
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 65654 60412 65962 60421
rect 65654 60410 65660 60412
rect 65716 60410 65740 60412
rect 65796 60410 65820 60412
rect 65876 60410 65900 60412
rect 65956 60410 65962 60412
rect 65716 60358 65718 60410
rect 65898 60358 65900 60410
rect 65654 60356 65660 60358
rect 65716 60356 65740 60358
rect 65796 60356 65820 60358
rect 65876 60356 65900 60358
rect 65956 60356 65962 60358
rect 65654 60347 65962 60356
rect 19574 59868 19882 59877
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59803 19882 59812
rect 50294 59868 50602 59877
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59803 50602 59812
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 34934 59324 35242 59333
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59259 35242 59268
rect 65654 59324 65962 59333
rect 65654 59322 65660 59324
rect 65716 59322 65740 59324
rect 65796 59322 65820 59324
rect 65876 59322 65900 59324
rect 65956 59322 65962 59324
rect 65716 59270 65718 59322
rect 65898 59270 65900 59322
rect 65654 59268 65660 59270
rect 65716 59268 65740 59270
rect 65796 59268 65820 59270
rect 65876 59268 65900 59270
rect 65956 59268 65962 59270
rect 65654 59259 65962 59268
rect 19574 58780 19882 58789
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58715 19882 58724
rect 50294 58780 50602 58789
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58715 50602 58724
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 34934 58236 35242 58245
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58171 35242 58180
rect 65654 58236 65962 58245
rect 65654 58234 65660 58236
rect 65716 58234 65740 58236
rect 65796 58234 65820 58236
rect 65876 58234 65900 58236
rect 65956 58234 65962 58236
rect 65716 58182 65718 58234
rect 65898 58182 65900 58234
rect 65654 58180 65660 58182
rect 65716 58180 65740 58182
rect 65796 58180 65820 58182
rect 65876 58180 65900 58182
rect 65956 58180 65962 58182
rect 65654 58171 65962 58180
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 68468 56160 68520 56166
rect 68468 56102 68520 56108
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 65654 56060 65962 56069
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 68480 55865 68508 56102
rect 68466 55856 68522 55865
rect 68466 55791 68522 55800
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 1768 46572 1820 46578
rect 1768 46514 1820 46520
rect 940 46368 992 46374
rect 938 46336 940 46345
rect 992 46336 994 46345
rect 938 46271 994 46280
rect 940 37188 992 37194
rect 940 37130 992 37136
rect 952 36825 980 37130
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 1780 19718 1808 46514
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 65654 46268 65962 46277
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 65654 44092 65962 44101
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 65654 40828 65962 40837
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 18236 37324 18288 37330
rect 18236 37266 18288 37272
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 17972 27010 18000 28358
rect 17880 26994 18000 27010
rect 17868 26988 18000 26994
rect 17920 26982 18000 26988
rect 17868 26930 17920 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 10416 26308 10468 26314
rect 10416 26250 10468 26256
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 10428 25362 10456 26250
rect 12452 25770 12480 26250
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13912 26240 13964 26246
rect 13912 26182 13964 26188
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 13832 25906 13860 26182
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 12440 25764 12492 25770
rect 12440 25706 12492 25712
rect 12728 25498 12756 25842
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12716 25492 12768 25498
rect 12716 25434 12768 25440
rect 12624 25424 12676 25430
rect 12624 25366 12676 25372
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 9312 24880 9364 24886
rect 9312 24822 9364 24828
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 7944 23662 7972 24550
rect 9324 24410 9352 24822
rect 9784 24698 9812 25298
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 9600 24682 9812 24698
rect 9864 24744 9916 24750
rect 10152 24698 10180 24754
rect 9864 24686 9916 24692
rect 9588 24676 9812 24682
rect 9640 24670 9812 24676
rect 9588 24618 9640 24624
rect 9876 24410 9904 24686
rect 10060 24670 10180 24698
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 7944 22642 7972 23598
rect 8864 23050 8892 24006
rect 9968 23866 9996 24142
rect 10060 23866 10088 24670
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10324 24336 10376 24342
rect 10324 24278 10376 24284
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 8944 23792 8996 23798
rect 8944 23734 8996 23740
rect 8956 23322 8984 23734
rect 9968 23594 9996 23802
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 8944 23316 8996 23322
rect 8944 23258 8996 23264
rect 8852 23044 8904 23050
rect 8852 22986 8904 22992
rect 7932 22636 7984 22642
rect 7932 22578 7984 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 8864 22030 8892 22986
rect 10060 22778 10088 23802
rect 10336 23730 10364 24278
rect 10508 24200 10560 24206
rect 10508 24142 10560 24148
rect 10520 23866 10548 24142
rect 10796 24138 10824 24550
rect 10784 24132 10836 24138
rect 10784 24074 10836 24080
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10612 23866 10640 24006
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10600 23860 10652 23866
rect 10600 23802 10652 23808
rect 10520 23730 10548 23802
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 8944 22704 8996 22710
rect 8944 22646 8996 22652
rect 8956 22234 8984 22646
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 8496 20534 8524 21286
rect 8864 20874 8892 21966
rect 9876 21554 9904 22578
rect 9968 22234 9996 22578
rect 10152 22506 10180 23054
rect 10336 22710 10364 23666
rect 10600 23044 10652 23050
rect 10600 22986 10652 22992
rect 10324 22704 10376 22710
rect 10324 22646 10376 22652
rect 10140 22500 10192 22506
rect 10140 22442 10192 22448
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 10336 21690 10364 22646
rect 10612 22642 10640 22986
rect 10692 22976 10744 22982
rect 10692 22918 10744 22924
rect 10704 22778 10732 22918
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10612 22030 10640 22578
rect 10888 22030 10916 22578
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10520 21894 10548 21966
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 10612 21010 10640 21966
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 8852 20868 8904 20874
rect 8852 20810 8904 20816
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8680 20534 8708 20742
rect 8484 20528 8536 20534
rect 8484 20470 8536 20476
rect 8668 20528 8720 20534
rect 8668 20470 8720 20476
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4066 18456 4122 18465
rect 7944 18426 7972 20334
rect 9416 19836 9444 20810
rect 9600 20058 9628 20878
rect 10336 20466 10364 20946
rect 10796 20874 10824 21626
rect 10888 21554 10916 21966
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10888 21418 10916 21490
rect 10876 21412 10928 21418
rect 10876 21354 10928 21360
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10324 20460 10376 20466
rect 10888 20448 10916 21354
rect 10980 21010 11008 25298
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 11164 24954 11192 25162
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 11992 24954 12020 25094
rect 12176 24954 12204 25094
rect 11152 24948 11204 24954
rect 11152 24890 11204 24896
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 11244 24880 11296 24886
rect 11244 24822 11296 24828
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 11164 24070 11192 24754
rect 11256 24206 11284 24822
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11532 24206 11560 24686
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11256 24070 11284 24142
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11348 23866 11376 24142
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11532 23798 11560 24142
rect 11992 23866 12020 24550
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 11520 23792 11572 23798
rect 11520 23734 11572 23740
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 11072 23322 11100 23666
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11348 23050 11376 23666
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11348 22778 11376 22986
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11532 22658 11560 23734
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11624 23254 11652 23462
rect 11612 23248 11664 23254
rect 11612 23190 11664 23196
rect 11624 22778 11652 23190
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11900 23050 11928 23122
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 11152 22636 11204 22642
rect 11532 22630 11652 22658
rect 11152 22578 11204 22584
rect 11164 21894 11192 22578
rect 11624 22574 11652 22630
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11624 22094 11652 22510
rect 11624 22066 11744 22094
rect 11716 21962 11744 22066
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11164 21554 11192 21830
rect 11900 21622 11928 22986
rect 12452 22642 12480 25094
rect 12636 24614 12664 25366
rect 12820 24886 12848 25774
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12636 24274 12664 24550
rect 12820 24410 12848 24822
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 12912 24410 12940 24550
rect 12808 24404 12860 24410
rect 12808 24346 12860 24352
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12900 24132 12952 24138
rect 12900 24074 12952 24080
rect 12912 23866 12940 24074
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 13096 23730 13124 24142
rect 13176 24064 13228 24070
rect 13176 24006 13228 24012
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 13004 23610 13032 23666
rect 13188 23610 13216 24006
rect 13372 23798 13400 25230
rect 13832 24818 13860 25842
rect 13924 25838 13952 26182
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 13924 25294 13952 25774
rect 14292 25498 14320 25774
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 14280 25492 14332 25498
rect 14280 25434 14332 25440
rect 15764 25362 15792 25638
rect 14004 25356 14056 25362
rect 14004 25298 14056 25304
rect 15752 25356 15804 25362
rect 15752 25298 15804 25304
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 14016 24954 14044 25298
rect 14004 24948 14056 24954
rect 14004 24890 14056 24896
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13360 23792 13412 23798
rect 13360 23734 13412 23740
rect 12544 23186 12572 23598
rect 13004 23582 13216 23610
rect 13268 23656 13320 23662
rect 13268 23598 13320 23604
rect 13188 23322 13216 23582
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 12532 23180 12584 23186
rect 12532 23122 12584 23128
rect 12808 23112 12860 23118
rect 13176 23112 13228 23118
rect 12860 23072 13124 23100
rect 12808 23054 12860 23060
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12176 22234 12204 22510
rect 12452 22386 12480 22578
rect 12544 22522 12572 22918
rect 12544 22494 12664 22522
rect 12452 22358 12572 22386
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 12440 22160 12492 22166
rect 12440 22102 12492 22108
rect 12452 21894 12480 22102
rect 12544 22030 12572 22358
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 11992 21690 12020 21830
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11164 21434 11192 21490
rect 11336 21480 11388 21486
rect 11164 21406 11284 21434
rect 11336 21422 11388 21428
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20602 11100 20878
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11060 20460 11112 20466
rect 10888 20420 11060 20448
rect 10324 20402 10376 20408
rect 11060 20402 11112 20408
rect 11072 20330 11100 20402
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 9496 19848 9548 19854
rect 9416 19808 9496 19836
rect 9496 19790 9548 19796
rect 9508 18766 9536 19790
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 4066 18391 4122 18400
rect 7932 18420 7984 18426
rect 4080 17338 4108 18391
rect 7932 18362 7984 18368
rect 9508 18358 9536 18566
rect 10152 18358 10180 18566
rect 9496 18352 9548 18358
rect 9496 18294 9548 18300
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 7760 17270 7788 18226
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8496 17882 8524 18158
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9140 17270 9168 17614
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 8496 16794 8524 17206
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8772 16794 8800 17070
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 7024 13938 7052 15438
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 7300 15162 7328 15370
rect 8588 15162 8616 15370
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8680 15026 8708 16594
rect 9324 16454 9352 16934
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 15910 9352 16390
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9508 15638 9536 16458
rect 9692 16250 9720 17138
rect 9876 17134 9904 18022
rect 10612 17882 10640 18702
rect 10888 18426 10916 19858
rect 11164 19786 11192 21286
rect 11256 20534 11284 21406
rect 11348 20942 11376 21422
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11440 20602 11468 20810
rect 11716 20602 11744 21490
rect 11900 21418 11928 21558
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 11888 21412 11940 21418
rect 11888 21354 11940 21360
rect 12268 20942 12296 21490
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 12256 20936 12308 20942
rect 12256 20878 12308 20884
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11704 20460 11756 20466
rect 11808 20448 11836 20742
rect 11756 20420 11836 20448
rect 11704 20402 11756 20408
rect 11900 20398 11928 20878
rect 12084 20602 12112 20878
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 12268 20262 12296 20878
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12268 19854 12296 20198
rect 12544 19922 12572 20810
rect 12636 20534 12664 22494
rect 12728 21554 12756 22918
rect 12912 22642 12940 22918
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12912 22234 12940 22374
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 13096 22166 13124 23072
rect 13176 23054 13228 23060
rect 13188 22778 13216 23054
rect 13280 22778 13308 23598
rect 13832 23186 13860 24754
rect 14016 24410 14044 24890
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14292 24410 14320 24754
rect 15764 24682 15792 25298
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 16040 24954 16068 25230
rect 16224 25226 16252 26182
rect 16304 25968 16356 25974
rect 16304 25910 16356 25916
rect 16316 25498 16344 25910
rect 17972 25906 18000 26982
rect 18248 26382 18276 37266
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 21088 28960 21140 28966
rect 21088 28902 21140 28908
rect 21100 28490 21128 28902
rect 20352 28484 20404 28490
rect 20352 28426 20404 28432
rect 21088 28484 21140 28490
rect 21088 28426 21140 28432
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 20364 28218 20392 28426
rect 20352 28212 20404 28218
rect 20352 28154 20404 28160
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 20996 27464 21048 27470
rect 20996 27406 21048 27412
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20640 27130 20668 27270
rect 21008 27130 21036 27406
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 20996 27124 21048 27130
rect 20996 27066 21048 27072
rect 18788 27056 18840 27062
rect 18788 26998 18840 27004
rect 18800 26586 18828 26998
rect 19800 26920 19852 26926
rect 19800 26862 19852 26868
rect 20352 26920 20404 26926
rect 20352 26862 20404 26868
rect 19708 26784 19760 26790
rect 19708 26726 19760 26732
rect 19720 26586 19748 26726
rect 19812 26586 19840 26862
rect 20260 26784 20312 26790
rect 20260 26726 20312 26732
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18788 26580 18840 26586
rect 18788 26522 18840 26528
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19800 26580 19852 26586
rect 19800 26522 19852 26528
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 16304 25492 16356 25498
rect 16304 25434 16356 25440
rect 17972 25362 18000 25842
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16212 25220 16264 25226
rect 16212 25162 16264 25168
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 15752 24676 15804 24682
rect 15752 24618 15804 24624
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 15764 24274 15792 24618
rect 15752 24268 15804 24274
rect 15752 24210 15804 24216
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 15384 24064 15436 24070
rect 15384 24006 15436 24012
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 14096 23180 14148 23186
rect 14096 23122 14148 23128
rect 13176 22772 13228 22778
rect 13176 22714 13228 22720
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 13280 22030 13308 22714
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13372 21672 13400 22034
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13280 21644 13400 21672
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 13280 20942 13308 21644
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13372 20942 13400 21490
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 13280 20466 13308 20878
rect 13556 20466 13584 21830
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13924 21554 13952 21626
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 13910 20496 13966 20505
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13544 20460 13596 20466
rect 13910 20431 13912 20440
rect 13544 20402 13596 20408
rect 13964 20431 13966 20440
rect 13912 20402 13964 20408
rect 13268 20256 13320 20262
rect 14016 20244 14044 21830
rect 14108 21486 14136 23122
rect 14384 23118 14412 23462
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14292 22778 14320 22918
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14568 22642 14596 23122
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14752 21554 14780 24006
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14844 22778 14872 22986
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14936 21690 14964 23258
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15028 22778 15056 22918
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 15212 22098 15240 22918
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 14924 21684 14976 21690
rect 14924 21626 14976 21632
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 14108 21010 14136 21422
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14292 21010 14320 21286
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14844 20602 14872 20810
rect 14936 20602 14964 21626
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 14096 20256 14148 20262
rect 14016 20216 14096 20244
rect 13268 20198 13320 20204
rect 14096 20198 14148 20204
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11624 19514 11652 19722
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11072 18766 11100 19246
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10888 17882 10916 18362
rect 10980 18290 11008 18566
rect 11532 18426 11560 18702
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12176 18426 12204 18566
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 11532 17746 11560 18362
rect 12544 18290 12572 19858
rect 12992 19780 13044 19786
rect 12992 19722 13044 19728
rect 13004 19514 13032 19722
rect 12992 19508 13044 19514
rect 12992 19450 13044 19456
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11624 17746 11652 18022
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10888 17270 10916 17478
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9968 16522 9996 17206
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9876 16182 9904 16458
rect 10060 16182 10088 16662
rect 10152 16590 10180 16934
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10416 16516 10468 16522
rect 10416 16458 10468 16464
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15366 9628 15506
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9048 15162 9076 15302
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 8128 13818 8156 13942
rect 8128 13790 8340 13818
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 8312 12850 8340 13790
rect 8588 13530 8616 13942
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8680 13326 8708 14962
rect 9508 14414 9536 15302
rect 9600 15094 9628 15302
rect 9692 15162 9720 15982
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 13802 8984 14214
rect 9140 14074 9168 14350
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9968 13938 9996 15030
rect 10152 14414 10180 15438
rect 10428 14414 10456 16458
rect 10704 16250 10732 17070
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 11072 15706 11100 16458
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 14822 11100 15438
rect 11164 15026 11192 15574
rect 11256 15502 11284 16050
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10152 14074 10180 14350
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 9968 13530 9996 13874
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 10428 13326 10456 14350
rect 10888 14006 10916 14554
rect 11072 14550 11100 14758
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 11072 14090 11100 14486
rect 10980 14074 11100 14090
rect 10968 14068 11100 14074
rect 11020 14062 11100 14068
rect 10968 14010 11020 14016
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10704 13530 10732 13942
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11072 13326 11100 13398
rect 11256 13326 11284 15438
rect 11348 15094 11376 15846
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11440 14618 11468 16662
rect 11532 16658 11560 17682
rect 11808 17542 11836 18022
rect 11796 17536 11848 17542
rect 11848 17496 11928 17524
rect 11796 17478 11848 17484
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11900 16590 11928 17496
rect 12636 16658 12664 18770
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13096 17882 13124 18566
rect 13188 18426 13216 18566
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13188 17746 13216 18226
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 17338 12756 17546
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11532 15502 11560 16050
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11532 15366 11560 15438
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11900 15094 11928 16526
rect 12268 16250 12296 16526
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12452 16250 12480 16390
rect 13096 16250 13124 16390
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13280 16114 13308 20198
rect 14108 19786 14136 20198
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14660 19446 14688 20198
rect 15212 20058 15240 20198
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13372 18358 13400 18702
rect 13464 18698 13492 19314
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14108 18902 14136 19246
rect 14292 18970 14320 19314
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13740 18426 13768 18566
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 13372 18170 13400 18294
rect 13372 18142 13492 18170
rect 13464 18086 13492 18142
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 14108 17954 14136 18838
rect 14476 18358 14504 19110
rect 15304 18766 15332 20334
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 15396 17954 15424 24006
rect 15948 23526 15976 24142
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15948 23118 15976 23462
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16132 22982 16160 23054
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15488 22234 15516 22578
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15948 20466 15976 20742
rect 16040 20466 16068 21354
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16040 20058 16068 20402
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15580 18834 15608 19722
rect 16224 19718 16252 25162
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16500 24834 16528 25094
rect 16592 24954 16620 25162
rect 16684 24954 16712 25230
rect 17960 25220 18012 25226
rect 17960 25162 18012 25168
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16672 24948 16724 24954
rect 16672 24890 16724 24896
rect 16304 24812 16356 24818
rect 16500 24806 16620 24834
rect 16304 24754 16356 24760
rect 16316 23866 16344 24754
rect 16592 24206 16620 24806
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16592 23322 16620 24142
rect 16684 24070 16712 24550
rect 16776 24410 16804 24754
rect 16764 24404 16816 24410
rect 16764 24346 16816 24352
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16684 23254 16712 24006
rect 17236 23662 17264 24006
rect 17512 23730 17540 24074
rect 17972 23866 18000 25162
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18064 24818 18092 25094
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18156 24410 18184 24550
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 16948 23588 17000 23594
rect 16948 23530 17000 23536
rect 16672 23248 16724 23254
rect 16672 23190 16724 23196
rect 16684 22710 16712 23190
rect 16672 22704 16724 22710
rect 16672 22646 16724 22652
rect 16960 22438 16988 23530
rect 17132 23248 17184 23254
rect 17132 23190 17184 23196
rect 17144 22778 17172 23190
rect 17236 23118 17264 23598
rect 17512 23186 17540 23666
rect 18064 23322 18092 23666
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17500 23180 17552 23186
rect 17500 23122 17552 23128
rect 17224 23112 17276 23118
rect 17224 23054 17276 23060
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17604 22642 17632 23054
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16684 22094 16712 22374
rect 16960 22234 16988 22374
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 17788 22094 17816 22918
rect 16592 22066 16712 22094
rect 17604 22066 17816 22094
rect 18248 22094 18276 26318
rect 18340 23594 18368 26522
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19352 26042 19380 26454
rect 20272 26382 20300 26726
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 20076 26308 20128 26314
rect 20128 26268 20208 26296
rect 20076 26250 20128 26256
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19444 25974 19472 26182
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18708 24682 18736 25230
rect 18696 24676 18748 24682
rect 18696 24618 18748 24624
rect 19076 24274 19104 25298
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19984 25220 20036 25226
rect 19984 25162 20036 25168
rect 19444 24954 19472 25162
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19996 24954 20024 25162
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19260 24410 19288 24754
rect 20180 24750 20208 26268
rect 20364 25974 20392 26862
rect 20444 26852 20496 26858
rect 20444 26794 20496 26800
rect 20456 26586 20484 26794
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20548 26586 20576 26726
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20536 26580 20588 26586
rect 20536 26522 20588 26528
rect 20352 25968 20404 25974
rect 20352 25910 20404 25916
rect 20640 25906 20668 27066
rect 20812 26988 20864 26994
rect 20812 26930 20864 26936
rect 20824 26586 20852 26930
rect 20812 26580 20864 26586
rect 20812 26522 20864 26528
rect 21192 26450 21220 28018
rect 21272 27328 21324 27334
rect 21272 27270 21324 27276
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21284 27130 21312 27270
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21284 26450 21312 27066
rect 21652 27062 21680 27270
rect 21640 27056 21692 27062
rect 21640 26998 21692 27004
rect 21652 26586 21680 26998
rect 21640 26580 21692 26586
rect 21640 26522 21692 26528
rect 21180 26444 21232 26450
rect 21180 26386 21232 26392
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21192 26042 21220 26386
rect 21652 26382 21680 26522
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21640 26376 21692 26382
rect 21640 26318 21692 26324
rect 21560 26042 21588 26318
rect 21180 26036 21232 26042
rect 21180 25978 21232 25984
rect 21548 26036 21600 26042
rect 21548 25978 21600 25984
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 21456 25220 21508 25226
rect 21456 25162 21508 25168
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 20824 24818 20852 25094
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20168 24744 20220 24750
rect 20168 24686 20220 24692
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 19892 24608 19944 24614
rect 19892 24550 19944 24556
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18524 23866 18552 24074
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 19076 23730 19104 24210
rect 19904 24138 19932 24550
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18328 23588 18380 23594
rect 18328 23530 18380 23536
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18432 23118 18460 23462
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18248 22066 18368 22094
rect 16592 22030 16620 22066
rect 17604 22030 17632 22066
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 18052 22024 18104 22030
rect 18104 21984 18184 22012
rect 18052 21966 18104 21972
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17328 20942 17356 21286
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17328 20534 17356 20742
rect 17316 20528 17368 20534
rect 17316 20470 17368 20476
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16224 19514 16252 19654
rect 16316 19514 16344 19722
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16302 19408 16358 19417
rect 16302 19343 16304 19352
rect 16356 19343 16358 19352
rect 17316 19372 17368 19378
rect 16304 19314 16356 19320
rect 17316 19314 17368 19320
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15488 18086 15516 18362
rect 15580 18154 15608 18770
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15568 18148 15620 18154
rect 15568 18090 15620 18096
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 14108 17926 14228 17954
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13740 16794 13768 17682
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15706 12204 15846
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11440 14278 11468 14554
rect 11900 14414 11928 15030
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12084 14482 12112 14554
rect 12176 14550 12204 14758
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11348 13394 11376 14214
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8956 12918 8984 13126
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 9600 12170 9628 13194
rect 10704 13190 10732 13262
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9692 12442 9720 12854
rect 10704 12782 10732 13126
rect 11072 12918 11100 13262
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11716 12850 11744 13262
rect 11900 12986 11928 13738
rect 11992 12986 12020 14282
rect 12268 14074 12296 15030
rect 12452 14890 12480 16050
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12544 13530 12572 15914
rect 12728 15162 12756 16050
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12912 15116 13124 15144
rect 12636 14940 12664 15098
rect 12912 15026 12940 15116
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12716 14952 12768 14958
rect 12636 14912 12716 14940
rect 12716 14894 12768 14900
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12176 13190 12204 13398
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 11532 12238 11560 12582
rect 11900 12306 11928 12922
rect 12176 12782 12204 13126
rect 12544 12850 12572 13466
rect 12728 13326 12756 14894
rect 13004 14346 13032 14962
rect 13096 14822 13124 15116
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14346 13124 14758
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 13394 12848 14214
rect 12912 14006 12940 14282
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 13096 13462 13124 14282
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 13648 12782 13676 13262
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9600 11762 9628 12106
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 10704 11354 10732 12038
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 11624 11150 11652 11494
rect 12176 11150 12204 12718
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12360 12306 12388 12582
rect 13648 12442 13676 12718
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 13004 11898 13032 12106
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 13740 3534 13768 15846
rect 13832 13394 13860 17138
rect 14200 16454 14228 17926
rect 15212 17926 15424 17954
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 17202 15148 17682
rect 15212 17202 15240 17926
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15396 17338 15424 17546
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15488 17202 15516 18022
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17202 15608 17478
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14740 16584 14792 16590
rect 14936 16572 14964 16934
rect 15028 16794 15056 17138
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 15580 16658 15608 17138
rect 16040 17134 16068 18566
rect 17328 18426 17356 19314
rect 17420 19174 17448 20742
rect 17604 20602 17632 21966
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17696 21554 17724 21830
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17972 21146 18000 21830
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 17592 20596 17644 20602
rect 17592 20538 17644 20544
rect 17972 20466 18000 21082
rect 18064 20602 18092 21422
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17420 18766 17448 19110
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 17202 16620 17478
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16776 17134 16804 18022
rect 17236 17338 17264 18158
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15016 16584 15068 16590
rect 14792 16544 15016 16572
rect 14740 16526 14792 16532
rect 15016 16526 15068 16532
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14200 15570 14228 16390
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14568 15434 14596 15982
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 15502 15240 15846
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 14188 15428 14240 15434
rect 14188 15370 14240 15376
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14108 15094 14136 15302
rect 14200 15162 14228 15370
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14568 15026 14596 15370
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 15304 14890 15332 15982
rect 15672 15910 15700 17070
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 15856 16250 15884 16934
rect 16408 16726 16436 16934
rect 16396 16720 16448 16726
rect 16396 16662 16448 16668
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15764 16130 15792 16186
rect 15948 16130 15976 16526
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 15764 16102 15976 16130
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 14752 14618 14780 14826
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 14924 14340 14976 14346
rect 14924 14282 14976 14288
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13924 13530 13952 13942
rect 14200 13802 14228 14214
rect 14936 14006 14964 14282
rect 15120 14006 15148 14350
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 15120 13394 15148 13942
rect 15212 13938 15240 14758
rect 15396 14414 15424 15438
rect 15672 14618 15700 15846
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 15026 15792 15302
rect 15948 15162 15976 16102
rect 16040 15978 16068 16390
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 16040 15706 16068 15914
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 16592 15434 16620 15982
rect 17512 15978 17540 18226
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 16592 15026 16620 15370
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 15856 14618 15884 14962
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 16868 14482 16896 15914
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17052 14618 17080 14894
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 17328 14414 17356 15846
rect 17420 14482 17448 15846
rect 17604 15570 17632 17070
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 16182 17724 16390
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17788 16046 17816 18226
rect 17880 17678 17908 18702
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18290 18000 18566
rect 18064 18426 18092 18702
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18156 18086 18184 21984
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18248 20874 18276 21286
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 18340 18714 18368 22066
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18432 21690 18460 21966
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18616 20466 18644 23598
rect 19076 22710 19104 23666
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 19076 22234 19104 22646
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19260 22386 19288 22578
rect 19168 22358 19288 22386
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 18788 22160 18840 22166
rect 18708 22108 18788 22114
rect 18708 22102 18840 22108
rect 18708 22086 18828 22102
rect 18708 21894 18736 22086
rect 19168 21962 19196 22358
rect 19248 22228 19300 22234
rect 19248 22170 19300 22176
rect 19260 22098 19288 22170
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18524 19514 18552 20198
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18432 18834 18460 19110
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18524 18766 18552 19450
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18512 18760 18564 18766
rect 18340 18686 18460 18714
rect 18512 18702 18564 18708
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18426 18368 18566
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18156 16794 18184 17138
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18248 16250 18276 17614
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18432 16114 18460 18686
rect 18616 18426 18644 18906
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18708 18290 18736 21830
rect 19076 21434 19104 21830
rect 19168 21622 19196 21898
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19076 21406 19196 21434
rect 19168 20942 19196 21406
rect 19260 21298 19288 22034
rect 19352 21690 19380 22918
rect 19444 22642 19472 23530
rect 19984 23520 20036 23526
rect 20088 23474 20116 24006
rect 20036 23468 20116 23474
rect 19984 23462 20116 23468
rect 19996 23446 20116 23462
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20088 22642 20116 23446
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 19720 22234 19748 22510
rect 19708 22228 19760 22234
rect 19708 22170 19760 22176
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19340 21344 19392 21350
rect 19260 21292 19340 21298
rect 19260 21286 19392 21292
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19260 21270 19380 21286
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 20088 20874 20116 21286
rect 20076 20868 20128 20874
rect 20076 20810 20128 20816
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20466 19380 20742
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19378 20024 19722
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19812 18970 19840 19314
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 18358 19380 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18420 19484 18426
rect 19484 18380 19564 18408
rect 19432 18362 19484 18368
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 18984 17338 19012 18158
rect 19352 17746 19380 18158
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18880 17264 18932 17270
rect 18878 17232 18880 17241
rect 18932 17232 18934 17241
rect 19076 17218 19104 17274
rect 18984 17202 19104 17218
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 18878 17167 18934 17176
rect 18972 17196 19104 17202
rect 19024 17190 19104 17196
rect 18972 17138 19024 17144
rect 19064 17128 19116 17134
rect 18970 17096 19026 17105
rect 19064 17070 19116 17076
rect 18970 17031 19026 17040
rect 18984 16794 19012 17031
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 16250 19012 16390
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17512 15162 17540 15370
rect 17696 15366 17724 15506
rect 18984 15502 19012 16050
rect 19076 15978 19104 17070
rect 19168 16674 19196 17206
rect 19352 17184 19380 17546
rect 19444 17542 19472 18090
rect 19536 17610 19564 18380
rect 20088 18222 20116 19994
rect 20180 19417 20208 24686
rect 20548 23866 20576 24686
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20272 23322 20300 23666
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 20732 22642 20760 24550
rect 20824 24410 20852 24754
rect 20812 24404 20864 24410
rect 20812 24346 20864 24352
rect 21468 24274 21496 25162
rect 21560 24818 21588 25842
rect 21744 24818 21772 29106
rect 23940 29096 23992 29102
rect 23940 29038 23992 29044
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 22100 28484 22152 28490
rect 22100 28426 22152 28432
rect 22468 28484 22520 28490
rect 22468 28426 22520 28432
rect 22112 28014 22140 28426
rect 22480 28218 22508 28426
rect 22468 28212 22520 28218
rect 22468 28154 22520 28160
rect 23308 28082 23336 28902
rect 23492 28490 23520 28902
rect 23480 28484 23532 28490
rect 23480 28426 23532 28432
rect 23952 28422 23980 29038
rect 24860 28960 24912 28966
rect 24860 28902 24912 28908
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 24676 28484 24728 28490
rect 24676 28426 24728 28432
rect 23940 28416 23992 28422
rect 23940 28358 23992 28364
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 23296 28076 23348 28082
rect 23296 28018 23348 28024
rect 22100 28008 22152 28014
rect 22100 27950 22152 27956
rect 22112 27538 22140 27950
rect 22388 27674 22416 28018
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22480 27130 22508 28018
rect 22572 27334 22600 28018
rect 22652 28008 22704 28014
rect 22652 27950 22704 27956
rect 22664 27606 22692 27950
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23756 27872 23808 27878
rect 23756 27814 23808 27820
rect 22652 27600 22704 27606
rect 22652 27542 22704 27548
rect 22928 27532 22980 27538
rect 22928 27474 22980 27480
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22940 27130 22968 27474
rect 23584 27470 23612 27814
rect 23768 27538 23796 27814
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23296 27396 23348 27402
rect 23296 27338 23348 27344
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 21824 26240 21876 26246
rect 21824 26182 21876 26188
rect 21836 25906 21864 26182
rect 22020 26042 22048 26318
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 21916 25900 21968 25906
rect 22020 25888 22048 25978
rect 21968 25860 22048 25888
rect 22100 25900 22152 25906
rect 21916 25842 21968 25848
rect 22100 25842 22152 25848
rect 22112 24818 22140 25842
rect 22204 25702 22232 26318
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21744 24070 21772 24754
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21928 24342 21956 24550
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 22112 24154 22140 24754
rect 22204 24342 22232 25638
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 22296 24800 22324 25298
rect 22376 24812 22428 24818
rect 22296 24772 22376 24800
rect 22376 24754 22428 24760
rect 22192 24336 22244 24342
rect 22192 24278 22244 24284
rect 22192 24200 22244 24206
rect 22112 24148 22192 24154
rect 22112 24142 22244 24148
rect 22112 24126 22232 24142
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21744 22642 21772 24006
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 22030 20760 22374
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20272 20942 20300 21898
rect 20916 21622 20944 22510
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20732 20602 20760 21422
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21008 21146 21036 21286
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20916 20466 20944 20742
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20272 19854 20300 20402
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20166 19408 20222 19417
rect 20166 19343 20222 19352
rect 20272 18766 20300 19790
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20640 18986 20668 19314
rect 20732 19242 20760 19790
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20810 19408 20866 19417
rect 20916 19378 20944 19654
rect 21008 19514 21036 21082
rect 21100 19854 21128 22578
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21376 22094 21404 22374
rect 21284 22066 21404 22094
rect 21284 21962 21312 22066
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21180 20392 21232 20398
rect 21180 20334 21232 20340
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21192 19378 21220 20334
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21376 20058 21404 20266
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21560 19446 21588 20878
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 20810 19343 20866 19352
rect 20904 19372 20956 19378
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20456 18958 20668 18986
rect 20456 18834 20484 18958
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20352 18760 20404 18766
rect 20720 18760 20772 18766
rect 20352 18702 20404 18708
rect 20640 18708 20720 18714
rect 20640 18702 20772 18708
rect 20168 18624 20220 18630
rect 20364 18612 20392 18702
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20640 18686 20760 18702
rect 20220 18584 20392 18612
rect 20168 18566 20220 18572
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19524 17604 19576 17610
rect 19524 17546 19576 17552
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19352 17156 19472 17184
rect 19444 16998 19472 17156
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19536 16810 19564 17002
rect 19352 16782 19564 16810
rect 19984 16788 20036 16794
rect 19246 16688 19302 16697
rect 19168 16646 19246 16674
rect 19246 16623 19302 16632
rect 19352 16590 19380 16782
rect 19984 16730 20036 16736
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 19352 15586 19380 16050
rect 19260 15558 19380 15586
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17604 14074 17632 14214
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17696 13938 17724 15302
rect 19260 15162 19288 15558
rect 19444 15162 19472 16662
rect 19536 16436 19564 16662
rect 19516 16408 19564 16436
rect 19516 16232 19544 16408
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19800 16244 19852 16250
rect 19516 16204 19564 16232
rect 19536 15570 19564 16204
rect 19800 16186 19852 16192
rect 19812 16114 19840 16186
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19812 15570 19840 16050
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19800 15564 19852 15570
rect 19996 15552 20024 16730
rect 20272 15706 20300 18584
rect 20456 18426 20484 18634
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20352 17808 20404 17814
rect 20352 17750 20404 17756
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 19800 15506 19852 15512
rect 19904 15524 20024 15552
rect 19536 15348 19564 15506
rect 19708 15496 19760 15502
rect 19904 15450 19932 15524
rect 20272 15502 20300 15642
rect 20260 15496 20312 15502
rect 19760 15444 19932 15450
rect 19708 15438 19932 15444
rect 19720 15422 19932 15438
rect 19996 15456 20260 15484
rect 19516 15320 19564 15348
rect 19516 15162 19544 15320
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19432 15156 19484 15162
rect 19516 15156 19576 15162
rect 19516 15116 19524 15156
rect 19432 15098 19484 15104
rect 19996 15144 20024 15456
rect 20260 15438 20312 15444
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 20088 15162 20116 15302
rect 19524 15098 19576 15104
rect 19904 15116 20024 15144
rect 20076 15156 20128 15162
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18878 14920 18934 14929
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18156 14074 18184 14350
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18524 14006 18552 14486
rect 18800 14482 18828 14894
rect 18984 14890 19012 14962
rect 18878 14855 18934 14864
rect 18972 14884 19024 14890
rect 18892 14822 18920 14855
rect 18972 14826 19024 14832
rect 19156 14884 19208 14890
rect 19156 14826 19208 14832
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 19168 14618 19196 14826
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 19444 13938 19472 14486
rect 19536 14414 19564 15098
rect 19904 14414 19932 15116
rect 20076 15098 20128 15104
rect 20364 14872 20392 17750
rect 20456 17134 20484 18362
rect 20640 17610 20668 18686
rect 20824 18358 20852 19343
rect 20904 19314 20956 19320
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21192 19242 21220 19314
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21284 19174 21312 19314
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 20916 18766 20944 19110
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20720 18352 20772 18358
rect 20720 18294 20772 18300
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20732 17882 20760 18294
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20824 17082 20852 18294
rect 20916 18154 20944 18702
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20824 17054 20944 17082
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20456 15026 20484 15914
rect 20548 15910 20576 16458
rect 20824 16182 20852 16934
rect 20812 16176 20864 16182
rect 20812 16118 20864 16124
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20732 15892 20760 16050
rect 20812 15904 20864 15910
rect 20732 15864 20812 15892
rect 20548 15026 20576 15846
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20640 15094 20668 15302
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20180 14844 20392 14872
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19708 14272 19760 14278
rect 19904 14260 19932 14350
rect 19760 14232 19932 14260
rect 19708 14214 19760 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14006 20024 14758
rect 20088 14618 20116 14758
rect 20180 14634 20208 14844
rect 20076 14612 20128 14618
rect 20180 14606 20392 14634
rect 20076 14554 20128 14560
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 13832 11626 13860 13330
rect 15120 12918 15148 13330
rect 17236 13326 17264 13670
rect 17880 13326 17908 13670
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15396 12782 15424 13194
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 12850 16988 13126
rect 17880 12986 17908 13262
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15488 12442 15516 12786
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 15476 12436 15528 12442
rect 17604 12434 17632 12582
rect 15476 12378 15528 12384
rect 17420 12406 17632 12434
rect 15488 11830 15516 12378
rect 17420 12238 17448 12406
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11830 16528 12106
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 14660 11150 14688 11630
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14660 10062 14688 11086
rect 16408 11082 16436 11494
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16500 10674 16528 11766
rect 17144 11762 17172 12174
rect 17512 11762 17540 12174
rect 17788 11898 17816 12718
rect 17880 12374 17908 12786
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17972 11898 18000 13466
rect 18248 13326 18276 13874
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18524 13530 18552 13806
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18236 13320 18288 13326
rect 18156 13268 18236 13274
rect 18156 13262 18288 13268
rect 18156 13246 18276 13262
rect 18156 12986 18184 13246
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18248 12850 18276 13126
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17144 11150 17172 11698
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17144 10674 17172 11086
rect 17880 10962 17908 11630
rect 18064 11614 18276 11642
rect 18064 11558 18092 11614
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18156 11354 18184 11494
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 17880 10934 18000 10962
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10062 16436 10406
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 14660 9518 14688 9998
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 7954 15608 9318
rect 15948 9178 15976 9590
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16500 8974 16528 10610
rect 17144 10538 17172 10610
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9518 16804 9998
rect 17144 9722 17172 10474
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 10266 17264 10406
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17038 9616 17094 9625
rect 16948 9580 17000 9586
rect 17420 9586 17448 9862
rect 17512 9722 17540 9998
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17604 9586 17632 10678
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17696 10062 17724 10610
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17038 9551 17040 9560
rect 16948 9522 17000 9528
rect 17092 9551 17094 9560
rect 17132 9580 17184 9586
rect 17040 9522 17092 9528
rect 17132 9522 17184 9528
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16960 9178 16988 9522
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15856 7342 15884 7890
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15948 7546 15976 7754
rect 16684 7546 16712 8230
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16776 7410 16804 8910
rect 17052 8634 17080 9522
rect 17144 8838 17172 9522
rect 17604 8974 17632 9522
rect 17696 9518 17724 9998
rect 17972 9586 18000 10934
rect 18064 10810 18092 11222
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18156 9654 18184 11086
rect 18248 10742 18276 11614
rect 18340 10742 18368 12038
rect 18432 10742 18460 12038
rect 19352 11801 19380 12038
rect 19338 11792 19394 11801
rect 19338 11727 19394 11736
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 11354 18736 11494
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18708 10742 18736 11154
rect 18800 11150 18828 11562
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18420 10736 18472 10742
rect 18696 10736 18748 10742
rect 18472 10696 18552 10724
rect 18420 10678 18472 10684
rect 18144 9648 18196 9654
rect 18524 9625 18552 10696
rect 18696 10678 18748 10684
rect 18708 10062 18736 10678
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18144 9590 18196 9596
rect 18510 9616 18566 9625
rect 17960 9580 18012 9586
rect 18510 9551 18566 9560
rect 17960 9522 18012 9528
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17696 9042 17724 9454
rect 17972 9110 18000 9522
rect 18604 9512 18656 9518
rect 18510 9480 18566 9489
rect 18604 9454 18656 9460
rect 18510 9415 18512 9424
rect 18564 9415 18566 9424
rect 18512 9386 18564 9392
rect 18616 9382 18644 9454
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 18328 9104 18380 9110
rect 18328 9046 18380 9052
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17144 8566 17172 8774
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17604 8430 17632 8910
rect 18340 8498 18368 9046
rect 18708 8838 18736 9998
rect 18892 9654 18920 9998
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18984 9586 19012 10406
rect 19076 10062 19104 10746
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 19076 9110 19104 9998
rect 19168 9489 19196 10542
rect 19260 10010 19288 11018
rect 19352 10742 19380 11290
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19352 10198 19380 10678
rect 19444 10674 19472 13874
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19628 12238 19656 12582
rect 20088 12442 20116 14350
rect 20272 13870 20300 14418
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20272 13394 20300 13806
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20272 12918 20300 13330
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 20088 12238 20116 12378
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19720 11354 19748 11766
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19996 11218 20024 12038
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19720 11082 19748 11154
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19432 10532 19484 10538
rect 19432 10474 19484 10480
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19260 9982 19380 10010
rect 19154 9480 19210 9489
rect 19154 9415 19210 9424
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 19260 9042 19288 9982
rect 19352 9926 19380 9982
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19444 9654 19472 10474
rect 19996 10130 20024 10610
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20088 10130 20116 10406
rect 20180 10266 20208 10950
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 18696 8832 18748 8838
rect 18748 8792 18920 8820
rect 18696 8774 18748 8780
rect 18694 8664 18750 8673
rect 18694 8599 18696 8608
rect 18748 8599 18750 8608
rect 18696 8570 18748 8576
rect 18892 8498 18920 8792
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17604 8090 17632 8366
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18524 8090 18552 8298
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18984 7886 19012 8978
rect 19352 8838 19380 9318
rect 19996 9160 20024 10066
rect 20272 9654 20300 10950
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20076 9172 20128 9178
rect 19996 9132 20076 9160
rect 20076 9114 20128 9120
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19154 8664 19210 8673
rect 19064 8628 19116 8634
rect 19154 8599 19210 8608
rect 19064 8570 19116 8576
rect 19076 8498 19104 8570
rect 19168 8566 19196 8599
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19076 7954 19104 8230
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 19168 7886 19196 8230
rect 19260 8090 19288 8298
rect 19352 8294 19380 8774
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8634 20024 8774
rect 20088 8634 20116 9114
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19628 7886 19656 8298
rect 20088 7954 20116 8570
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16868 7546 16896 7754
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17880 7546 17908 7686
rect 18984 7546 19012 7822
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7546 19288 7686
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 16776 7002 16804 7346
rect 18340 7002 18368 7414
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19536 7002 19564 7142
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19812 6798 19840 7346
rect 20088 6866 20116 7890
rect 20180 7478 20208 8230
rect 20168 7472 20220 7478
rect 20168 7414 20220 7420
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8404 800 8432 3470
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20364 3058 20392 14606
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20456 13870 20484 14214
rect 20640 14074 20668 15030
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20456 12986 20484 13262
rect 20732 13138 20760 15864
rect 20812 15846 20864 15852
rect 20640 13110 20760 13138
rect 20640 12986 20668 13110
rect 20916 12986 20944 17054
rect 21008 16114 21036 18158
rect 21652 17746 21680 19314
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21928 18290 21956 18906
rect 22112 18834 22140 21830
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22204 19854 22232 20198
rect 22296 19990 22324 24074
rect 22480 23662 22508 26250
rect 22664 26042 22692 26862
rect 22756 26586 22784 27066
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22848 26790 22876 26930
rect 22928 26852 22980 26858
rect 22928 26794 22980 26800
rect 22836 26784 22888 26790
rect 22836 26726 22888 26732
rect 22744 26580 22796 26586
rect 22744 26522 22796 26528
rect 22756 26314 22784 26522
rect 22744 26308 22796 26314
rect 22744 26250 22796 26256
rect 22652 26036 22704 26042
rect 22652 25978 22704 25984
rect 22744 25900 22796 25906
rect 22744 25842 22796 25848
rect 22756 25430 22784 25842
rect 22848 25498 22876 26726
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22744 25424 22796 25430
rect 22744 25366 22796 25372
rect 22560 25220 22612 25226
rect 22560 25162 22612 25168
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22572 24954 22600 25162
rect 22664 24954 22692 25162
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22652 24948 22704 24954
rect 22652 24890 22704 24896
rect 22940 24834 22968 26794
rect 23032 25158 23060 27270
rect 23308 27130 23336 27338
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 23308 26518 23336 27066
rect 23400 26858 23428 27406
rect 23584 27062 23612 27406
rect 23952 27402 23980 28358
rect 24216 27600 24268 27606
rect 24216 27542 24268 27548
rect 23940 27396 23992 27402
rect 23940 27338 23992 27344
rect 24228 27062 24256 27542
rect 24688 27130 24716 28426
rect 24872 28150 24900 28902
rect 25148 28490 25176 28902
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 25412 28620 25464 28626
rect 25412 28562 25464 28568
rect 25136 28484 25188 28490
rect 25136 28426 25188 28432
rect 25424 28150 25452 28562
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 24860 28144 24912 28150
rect 24860 28086 24912 28092
rect 25412 28144 25464 28150
rect 25412 28086 25464 28092
rect 25044 28008 25096 28014
rect 25044 27950 25096 27956
rect 25056 27674 25084 27950
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 25424 27606 25452 28086
rect 25412 27600 25464 27606
rect 25412 27542 25464 27548
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 24768 27396 24820 27402
rect 24768 27338 24820 27344
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 24780 27130 24808 27338
rect 24676 27124 24728 27130
rect 24676 27066 24728 27072
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 24216 27056 24268 27062
rect 24216 26998 24268 27004
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23388 26852 23440 26858
rect 23388 26794 23440 26800
rect 23492 26586 23520 26930
rect 23664 26920 23716 26926
rect 23664 26862 23716 26868
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 23296 26512 23348 26518
rect 23296 26454 23348 26460
rect 23676 26450 23704 26862
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23664 26444 23716 26450
rect 23664 26386 23716 26392
rect 23112 26240 23164 26246
rect 23112 26182 23164 26188
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 23124 24954 23152 26182
rect 23860 25906 23888 26726
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23204 25696 23256 25702
rect 23204 25638 23256 25644
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 23112 24948 23164 24954
rect 23112 24890 23164 24896
rect 22664 24806 22968 24834
rect 22664 24206 22692 24806
rect 23216 24596 23244 25638
rect 23296 25492 23348 25498
rect 23296 25434 23348 25440
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23308 25294 23336 25434
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23584 24886 23612 25434
rect 23664 25220 23716 25226
rect 23664 25162 23716 25168
rect 23572 24880 23624 24886
rect 23572 24822 23624 24828
rect 23676 24698 23704 25162
rect 23584 24682 23704 24698
rect 23572 24676 23704 24682
rect 23624 24670 23704 24676
rect 23572 24618 23624 24624
rect 23296 24608 23348 24614
rect 23216 24568 23296 24596
rect 23296 24550 23348 24556
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22664 23662 22692 24142
rect 22928 24064 22980 24070
rect 22928 24006 22980 24012
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22756 22778 22784 23666
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22848 23118 22876 23598
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22848 22166 22876 23054
rect 22836 22160 22888 22166
rect 22836 22102 22888 22108
rect 22940 22094 22968 24006
rect 23308 23526 23336 24550
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23020 23044 23072 23050
rect 23020 22986 23072 22992
rect 23032 22710 23060 22986
rect 23020 22704 23072 22710
rect 23020 22646 23072 22652
rect 22940 22066 23060 22094
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 22848 21486 22876 21898
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22388 20602 22416 20742
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22376 20324 22428 20330
rect 22376 20266 22428 20272
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22296 19446 22324 19926
rect 22388 19854 22416 20266
rect 22480 20058 22508 20810
rect 22558 20496 22614 20505
rect 22558 20431 22614 20440
rect 22572 20058 22600 20431
rect 22848 20262 22876 21422
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22940 20534 22968 20878
rect 22928 20528 22980 20534
rect 22928 20470 22980 20476
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22296 18834 22324 19382
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21824 18216 21876 18222
rect 21824 18158 21876 18164
rect 21836 17746 21864 18158
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21824 17740 21876 17746
rect 21824 17682 21876 17688
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21100 14074 21128 17478
rect 21652 17202 21680 17682
rect 22112 17542 22140 18566
rect 22296 17882 22324 18770
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22296 17762 22324 17818
rect 22296 17734 22416 17762
rect 22388 17610 22416 17734
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16114 21220 16390
rect 21284 16250 21312 17070
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21836 16250 21864 16458
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21192 15570 21220 16050
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21468 15502 21496 15846
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 21744 15502 21772 15642
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21652 14958 21680 15370
rect 22112 15026 22140 16526
rect 22204 15434 22232 17478
rect 22296 17202 22324 17478
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16114 22416 16934
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22480 15314 22508 19790
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22664 18698 22692 19722
rect 22940 19378 22968 20470
rect 23032 20058 23060 22066
rect 23124 22030 23152 23054
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23308 22778 23336 22918
rect 23400 22778 23428 23666
rect 23296 22772 23348 22778
rect 23296 22714 23348 22720
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23216 22094 23244 22578
rect 23664 22500 23716 22506
rect 23664 22442 23716 22448
rect 23216 22066 23336 22094
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21690 23152 21966
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23124 20602 23152 20810
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23308 20466 23336 22066
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23400 21418 23428 21898
rect 23676 21486 23704 22442
rect 23860 22098 23888 22714
rect 23848 22092 23900 22098
rect 23848 22034 23900 22040
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23388 21412 23440 21418
rect 23388 21354 23440 21360
rect 23400 20466 23428 21354
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23492 20466 23520 21286
rect 23952 21010 23980 21490
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 23308 19854 23336 20402
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22664 18426 22692 18634
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22572 15706 22600 15846
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22664 15502 22692 17002
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22756 16250 22784 16390
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22296 15286 22508 15314
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21652 14618 21680 14894
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 22112 14346 22140 14962
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21456 13252 21508 13258
rect 21456 13194 21508 13200
rect 21468 12986 21496 13194
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20628 12980 20680 12986
rect 20904 12980 20956 12986
rect 20628 12922 20680 12928
rect 20732 12940 20904 12968
rect 20640 12374 20668 12922
rect 20732 12442 20760 12940
rect 20904 12922 20956 12928
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20640 11354 20668 12310
rect 20916 12170 20944 12718
rect 21560 12434 21588 12718
rect 21376 12406 21588 12434
rect 21376 12170 21404 12406
rect 21836 12238 21864 13126
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22112 12442 22140 12718
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 20916 11558 20944 12106
rect 21376 11898 21404 12106
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21824 11824 21876 11830
rect 21822 11792 21824 11801
rect 21876 11792 21878 11801
rect 21732 11756 21784 11762
rect 21928 11762 21956 12174
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 21822 11727 21878 11736
rect 21916 11756 21968 11762
rect 21732 11698 21784 11704
rect 21916 11698 21968 11704
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20916 11218 20944 11494
rect 21744 11354 21772 11698
rect 22204 11694 22232 12038
rect 22296 11778 22324 15286
rect 22756 14414 22784 15302
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22468 13796 22520 13802
rect 22468 13738 22520 13744
rect 22480 13394 22508 13738
rect 22848 13530 22876 18702
rect 22940 18290 22968 19314
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23216 18426 23244 18702
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 23308 18086 23336 19314
rect 23400 18766 23428 20198
rect 23768 19854 23796 20198
rect 23952 20058 23980 20946
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23952 19854 23980 19994
rect 24044 19990 24072 25638
rect 24228 25294 24256 26998
rect 25056 26994 25084 27338
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 25044 26988 25096 26994
rect 25044 26930 25096 26936
rect 24216 25288 24268 25294
rect 24216 25230 24268 25236
rect 24320 23866 24348 26930
rect 25332 26926 25360 27406
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25424 26450 25452 27406
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 25504 27056 25556 27062
rect 25504 26998 25556 27004
rect 25516 26858 25544 26998
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25504 26852 25556 26858
rect 25504 26794 25556 26800
rect 25516 26586 25544 26794
rect 25504 26580 25556 26586
rect 25504 26522 25556 26528
rect 25412 26444 25464 26450
rect 25412 26386 25464 26392
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 24952 26240 25004 26246
rect 24952 26182 25004 26188
rect 24964 25906 24992 26182
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 24780 25498 24808 25842
rect 25044 25832 25096 25838
rect 25044 25774 25096 25780
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24584 24880 24636 24886
rect 24584 24822 24636 24828
rect 24596 24410 24624 24822
rect 24676 24608 24728 24614
rect 24872 24596 24900 25298
rect 25056 25294 25084 25774
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 24952 24948 25004 24954
rect 25004 24908 25084 24936
rect 24952 24890 25004 24896
rect 24728 24568 24900 24596
rect 24676 24550 24728 24556
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 24308 23860 24360 23866
rect 24308 23802 24360 23808
rect 24584 23520 24636 23526
rect 24584 23462 24636 23468
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 24136 22778 24164 23054
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 24228 21962 24256 22578
rect 24320 22030 24348 22714
rect 24596 22522 24624 23462
rect 24688 23118 24716 24550
rect 25056 23662 25084 24908
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24688 22642 24716 23054
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 24412 22494 24624 22522
rect 24412 22030 24440 22494
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24216 21956 24268 21962
rect 24216 21898 24268 21904
rect 24228 21418 24256 21898
rect 24216 21412 24268 21418
rect 24216 21354 24268 21360
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 24228 20398 24256 21082
rect 24412 20890 24440 21966
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24504 21486 24532 21830
rect 24688 21554 24716 21898
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24320 20862 24440 20890
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24320 20262 24348 20862
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 24412 20466 24440 20742
rect 24688 20602 24716 20878
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24032 19984 24084 19990
rect 24032 19926 24084 19932
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23492 18850 23520 19110
rect 23584 18970 23612 19790
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24596 19378 24624 19654
rect 24584 19372 24636 19378
rect 24780 19334 24808 22646
rect 24584 19314 24636 19320
rect 24688 19306 24808 19334
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23676 18850 23704 18906
rect 23492 18822 23704 18850
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23296 18080 23348 18086
rect 23296 18022 23348 18028
rect 23308 17746 23336 18022
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 23296 17740 23348 17746
rect 23296 17682 23348 17688
rect 23032 15502 23060 17682
rect 23204 17604 23256 17610
rect 23204 17546 23256 17552
rect 23112 17264 23164 17270
rect 23110 17232 23112 17241
rect 23164 17232 23166 17241
rect 23110 17167 23166 17176
rect 23216 17134 23244 17546
rect 23204 17128 23256 17134
rect 23492 17105 23520 18822
rect 23952 17746 23980 19110
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24412 17882 24440 18226
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23204 17070 23256 17076
rect 23478 17096 23534 17105
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23124 16590 23152 16934
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23216 15706 23244 17070
rect 23478 17031 23534 17040
rect 23768 16454 23796 17614
rect 23848 17604 23900 17610
rect 23848 17546 23900 17552
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23296 16108 23348 16114
rect 23296 16050 23348 16056
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23308 15502 23336 16050
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23400 15706 23428 15846
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23032 14414 23060 15438
rect 23492 15162 23520 15438
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23584 15026 23612 15302
rect 23768 15162 23796 16390
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 23032 13870 23060 14350
rect 23662 14104 23718 14113
rect 23662 14039 23664 14048
rect 23716 14039 23718 14048
rect 23664 14010 23716 14016
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22480 11830 22508 13330
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22848 12986 22876 13126
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 23124 12850 23152 13874
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23492 12850 23520 13806
rect 23768 13394 23796 15098
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23124 12238 23152 12786
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 22560 11892 22612 11898
rect 22560 11834 22612 11840
rect 22468 11824 22520 11830
rect 22296 11750 22416 11778
rect 22468 11766 22520 11772
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 21744 11150 21772 11290
rect 21836 11150 21864 11630
rect 22204 11218 22232 11630
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20732 10810 20760 11018
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20548 9178 20576 9522
rect 20732 9466 20760 10746
rect 20824 10266 20852 11086
rect 22296 10810 22324 11630
rect 22388 11626 22416 11750
rect 22376 11620 22428 11626
rect 22376 11562 22428 11568
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22480 10742 22508 11766
rect 22468 10736 22520 10742
rect 22468 10678 22520 10684
rect 22572 10674 22600 11834
rect 23860 11150 23888 17546
rect 24688 17338 24716 19306
rect 25056 18834 25084 23598
rect 25148 22778 25176 25842
rect 25332 25838 25360 26318
rect 25516 26042 25544 26522
rect 25608 26382 25636 26930
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25504 26036 25556 26042
rect 25504 25978 25556 25984
rect 25320 25832 25372 25838
rect 25320 25774 25372 25780
rect 25596 25764 25648 25770
rect 25596 25706 25648 25712
rect 25320 25696 25372 25702
rect 25320 25638 25372 25644
rect 25332 25294 25360 25638
rect 25608 25294 25636 25706
rect 25792 25294 25820 27270
rect 25976 27062 26004 28426
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 68836 28076 68888 28082
rect 68836 28018 68888 28024
rect 68848 27985 68876 28018
rect 68834 27976 68890 27985
rect 68834 27911 68890 27920
rect 68284 27872 68336 27878
rect 68284 27814 68336 27820
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 30564 27464 30616 27470
rect 30564 27406 30616 27412
rect 25964 27056 26016 27062
rect 25964 26998 26016 27004
rect 26068 25362 26096 27406
rect 26608 27396 26660 27402
rect 26608 27338 26660 27344
rect 28632 27396 28684 27402
rect 28632 27338 28684 27344
rect 26620 27130 26648 27338
rect 27712 27328 27764 27334
rect 27712 27270 27764 27276
rect 26608 27124 26660 27130
rect 26608 27066 26660 27072
rect 27724 26994 27752 27270
rect 28644 27130 28672 27338
rect 29368 27328 29420 27334
rect 29368 27270 29420 27276
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 30288 27328 30340 27334
rect 30288 27270 30340 27276
rect 28632 27124 28684 27130
rect 28632 27066 28684 27072
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 27080 25974 27108 26318
rect 27068 25968 27120 25974
rect 27068 25910 27120 25916
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 26056 25356 26108 25362
rect 26056 25298 26108 25304
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25780 25288 25832 25294
rect 25780 25230 25832 25236
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25504 25220 25556 25226
rect 25504 25162 25556 25168
rect 25424 24954 25452 25162
rect 25516 24954 25544 25162
rect 25412 24948 25464 24954
rect 25412 24890 25464 24896
rect 25504 24948 25556 24954
rect 25504 24890 25556 24896
rect 25780 24812 25832 24818
rect 25780 24754 25832 24760
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 25320 24064 25372 24070
rect 25320 24006 25372 24012
rect 25332 23866 25360 24006
rect 25700 23866 25728 24142
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25792 23730 25820 24754
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 25228 23656 25280 23662
rect 25228 23598 25280 23604
rect 25240 23322 25268 23598
rect 25596 23520 25648 23526
rect 25596 23462 25648 23468
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 25608 23050 25636 23462
rect 25792 23322 25820 23666
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 25596 23044 25648 23050
rect 25596 22986 25648 22992
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 26068 22710 26096 23054
rect 26056 22704 26108 22710
rect 26056 22646 26108 22652
rect 25504 22432 25556 22438
rect 25504 22374 25556 22380
rect 25516 22234 25544 22374
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25240 20806 25268 21422
rect 25424 21146 25452 21490
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 25240 19922 25268 20742
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25516 18850 25544 22170
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25700 21554 25728 21830
rect 26252 21622 26280 25842
rect 27172 25770 27200 26862
rect 27448 26586 27476 26862
rect 27724 26586 27752 26930
rect 28828 26586 28856 26930
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 28540 26580 28592 26586
rect 28540 26522 28592 26528
rect 28816 26580 28868 26586
rect 28816 26522 28868 26528
rect 27448 25906 27476 26522
rect 27804 26376 27856 26382
rect 27804 26318 27856 26324
rect 27712 26240 27764 26246
rect 27712 26182 27764 26188
rect 27724 25906 27752 26182
rect 27436 25900 27488 25906
rect 27436 25842 27488 25848
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 27712 25900 27764 25906
rect 27712 25842 27764 25848
rect 27160 25764 27212 25770
rect 27160 25706 27212 25712
rect 26700 25696 26752 25702
rect 26700 25638 26752 25644
rect 26712 25294 26740 25638
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26976 24064 27028 24070
rect 26976 24006 27028 24012
rect 26988 23866 27016 24006
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 26516 23724 26568 23730
rect 26516 23666 26568 23672
rect 26332 22568 26384 22574
rect 26332 22510 26384 22516
rect 26344 21690 26372 22510
rect 26424 22500 26476 22506
rect 26424 22442 26476 22448
rect 26436 22234 26464 22442
rect 26424 22228 26476 22234
rect 26424 22170 26476 22176
rect 26528 21706 26556 23666
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26712 23118 26740 23462
rect 26700 23112 26752 23118
rect 26700 23054 26752 23060
rect 26896 22166 26924 23598
rect 27172 23594 27200 25706
rect 27632 25498 27660 25842
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 27724 25362 27752 25842
rect 27816 25702 27844 26318
rect 28080 26308 28132 26314
rect 28080 26250 28132 26256
rect 27896 26240 27948 26246
rect 27896 26182 27948 26188
rect 27908 25906 27936 26182
rect 27896 25900 27948 25906
rect 27896 25842 27948 25848
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 27712 25356 27764 25362
rect 27712 25298 27764 25304
rect 27724 25242 27752 25298
rect 27816 25294 27844 25638
rect 27908 25430 27936 25842
rect 27896 25424 27948 25430
rect 27896 25366 27948 25372
rect 28092 25362 28120 26250
rect 28552 26042 28580 26522
rect 29380 26314 29408 27270
rect 29564 27130 29592 27270
rect 30300 27130 30328 27270
rect 29552 27124 29604 27130
rect 29552 27066 29604 27072
rect 30288 27124 30340 27130
rect 30288 27066 30340 27072
rect 29736 26784 29788 26790
rect 29736 26726 29788 26732
rect 30288 26784 30340 26790
rect 30288 26726 30340 26732
rect 29748 26382 29776 26726
rect 29736 26376 29788 26382
rect 29736 26318 29788 26324
rect 29368 26308 29420 26314
rect 29368 26250 29420 26256
rect 28724 26240 28776 26246
rect 28724 26182 28776 26188
rect 29276 26240 29328 26246
rect 30300 26228 30328 26726
rect 30470 26480 30526 26489
rect 30470 26415 30472 26424
rect 30524 26415 30526 26424
rect 30472 26386 30524 26392
rect 30472 26240 30524 26246
rect 30300 26200 30420 26228
rect 29276 26182 29328 26188
rect 28540 26036 28592 26042
rect 28540 25978 28592 25984
rect 28736 25362 28764 26182
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 28816 25764 28868 25770
rect 28816 25706 28868 25712
rect 28080 25356 28132 25362
rect 28080 25298 28132 25304
rect 28724 25356 28776 25362
rect 28724 25298 28776 25304
rect 27632 25214 27752 25242
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27632 24818 27660 25214
rect 27712 25152 27764 25158
rect 27712 25094 27764 25100
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 27356 23866 27384 24142
rect 27344 23860 27396 23866
rect 27344 23802 27396 23808
rect 27160 23588 27212 23594
rect 27160 23530 27212 23536
rect 27528 23588 27580 23594
rect 27528 23530 27580 23536
rect 26884 22160 26936 22166
rect 26884 22102 26936 22108
rect 26700 21888 26752 21894
rect 26700 21830 26752 21836
rect 26332 21684 26384 21690
rect 26528 21678 26648 21706
rect 26332 21626 26384 21632
rect 26240 21616 26292 21622
rect 26292 21564 26556 21570
rect 26240 21558 26556 21564
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25688 21548 25740 21554
rect 26252 21542 26556 21558
rect 25688 21490 25740 21496
rect 25608 21418 25636 21490
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 26424 21480 26476 21486
rect 26424 21422 26476 21428
rect 25596 21412 25648 21418
rect 25596 21354 25648 21360
rect 25608 18970 25636 21354
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25792 20942 25820 21286
rect 26252 20942 26280 21422
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26252 20534 26280 20878
rect 26436 20602 26464 21422
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26240 20528 26292 20534
rect 26240 20470 26292 20476
rect 26252 19922 26280 20470
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 26528 19446 26556 21542
rect 26620 21418 26648 21678
rect 26608 21412 26660 21418
rect 26608 21354 26660 21360
rect 26712 20942 26740 21830
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 26516 19440 26568 19446
rect 26516 19382 26568 19388
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25700 18970 25728 19314
rect 26896 19174 26924 22102
rect 27540 22094 27568 23530
rect 27632 23254 27660 24210
rect 27724 23662 27752 25094
rect 28092 24818 28120 25298
rect 28736 24818 28764 25298
rect 28828 25294 28856 25706
rect 28816 25288 28868 25294
rect 28816 25230 28868 25236
rect 29092 25152 29144 25158
rect 29092 25094 29144 25100
rect 29104 24954 29132 25094
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 28080 24812 28132 24818
rect 28000 24772 28080 24800
rect 28000 24206 28028 24772
rect 28080 24754 28132 24760
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28172 24744 28224 24750
rect 28172 24686 28224 24692
rect 28080 24608 28132 24614
rect 28080 24550 28132 24556
rect 28092 24274 28120 24550
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 28184 24206 28212 24686
rect 29196 24682 29224 25842
rect 29288 25702 29316 26182
rect 29920 25832 29972 25838
rect 29920 25774 29972 25780
rect 29276 25696 29328 25702
rect 29276 25638 29328 25644
rect 29368 25696 29420 25702
rect 29368 25638 29420 25644
rect 29288 25498 29316 25638
rect 29380 25498 29408 25638
rect 29276 25492 29328 25498
rect 29276 25434 29328 25440
rect 29368 25492 29420 25498
rect 29368 25434 29420 25440
rect 29184 24676 29236 24682
rect 29184 24618 29236 24624
rect 29288 24274 29316 25434
rect 29552 24608 29604 24614
rect 29552 24550 29604 24556
rect 29276 24268 29328 24274
rect 29276 24210 29328 24216
rect 27988 24200 28040 24206
rect 27988 24142 28040 24148
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 27896 24064 27948 24070
rect 27896 24006 27948 24012
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27724 23322 27752 23598
rect 27908 23322 27936 24006
rect 28184 23866 28212 24142
rect 28172 23860 28224 23866
rect 28172 23802 28224 23808
rect 28368 23322 28396 24142
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28552 23866 28580 24006
rect 28540 23860 28592 23866
rect 28540 23802 28592 23808
rect 29092 23656 29144 23662
rect 29092 23598 29144 23604
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 28356 23316 28408 23322
rect 28356 23258 28408 23264
rect 27620 23248 27672 23254
rect 27620 23190 27672 23196
rect 29104 23186 29132 23598
rect 29092 23180 29144 23186
rect 29092 23122 29144 23128
rect 28080 23044 28132 23050
rect 28080 22986 28132 22992
rect 28264 23044 28316 23050
rect 28264 22986 28316 22992
rect 27540 22066 27660 22094
rect 27160 21888 27212 21894
rect 27212 21836 27292 21842
rect 27160 21830 27292 21836
rect 27172 21814 27292 21830
rect 27264 19334 27292 21814
rect 27528 19916 27580 19922
rect 27528 19858 27580 19864
rect 27080 19306 27292 19334
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 26884 19168 26936 19174
rect 26884 19110 26936 19116
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25044 18828 25096 18834
rect 25516 18822 25820 18850
rect 25044 18770 25096 18776
rect 25056 18358 25084 18770
rect 25596 18760 25648 18766
rect 25596 18702 25648 18708
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 25424 17678 25452 18022
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23952 15502 23980 15982
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24504 15162 24532 15370
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 24122 15056 24178 15065
rect 24122 14991 24124 15000
rect 24176 14991 24178 15000
rect 24492 15020 24544 15026
rect 24124 14962 24176 14968
rect 24492 14962 24544 14968
rect 24504 14618 24532 14962
rect 24584 14884 24636 14890
rect 24584 14826 24636 14832
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24596 14550 24624 14826
rect 24584 14544 24636 14550
rect 24584 14486 24636 14492
rect 24688 14362 24716 17274
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 24964 16250 24992 16390
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24780 14929 24808 14962
rect 24766 14920 24822 14929
rect 24766 14855 24822 14864
rect 24872 14482 24900 15370
rect 25056 15314 25084 16594
rect 25148 16130 25176 17614
rect 25516 17338 25544 18226
rect 25608 18086 25636 18702
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25596 18080 25648 18086
rect 25596 18022 25648 18028
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25700 17066 25728 18226
rect 25228 17060 25280 17066
rect 25228 17002 25280 17008
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25240 16726 25268 17002
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25228 16176 25280 16182
rect 25148 16124 25228 16130
rect 25148 16118 25280 16124
rect 25148 16102 25268 16118
rect 25148 15502 25176 16102
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25056 15286 25176 15314
rect 25044 15088 25096 15094
rect 25044 15030 25096 15036
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24768 14408 24820 14414
rect 24688 14356 24768 14362
rect 24688 14350 24820 14356
rect 24688 14334 24808 14350
rect 24688 14278 24716 14334
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24872 14074 24900 14418
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24768 14000 24820 14006
rect 24964 13954 24992 14486
rect 24820 13948 24992 13954
rect 24768 13942 24992 13948
rect 24780 13926 24992 13942
rect 25056 13938 25084 15030
rect 25148 14618 25176 15286
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25240 13938 25268 14214
rect 24964 13818 24992 13926
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 24964 13790 25176 13818
rect 24952 12708 25004 12714
rect 24952 12650 25004 12656
rect 24964 12238 24992 12650
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23952 11354 23980 11766
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21088 9512 21140 9518
rect 20732 9438 20852 9466
rect 21088 9454 21140 9460
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20548 8362 20576 9114
rect 20732 8566 20760 9318
rect 20824 8634 20852 9438
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20916 8906 20944 9386
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 21008 9178 21036 9318
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20904 8900 20956 8906
rect 20904 8842 20956 8848
rect 21100 8634 21128 9454
rect 21284 8634 21312 9590
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21560 8838 21588 9522
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 21928 8498 21956 9454
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22296 9110 22324 9318
rect 22572 9194 22600 10610
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23032 10130 23060 10406
rect 23676 10266 23704 10678
rect 23664 10260 23716 10266
rect 23664 10202 23716 10208
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 23032 9722 23060 10066
rect 23860 9994 23888 11086
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24504 10266 24532 10542
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24780 10146 24808 12038
rect 24964 11898 24992 12174
rect 25056 11898 25084 12242
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24872 11354 24900 11630
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 25148 11082 25176 13790
rect 25332 12288 25360 15370
rect 25424 14958 25452 16594
rect 25700 15502 25728 17002
rect 25792 16590 25820 18822
rect 25872 18692 25924 18698
rect 25872 18634 25924 18640
rect 25884 18154 25912 18634
rect 25964 18284 26016 18290
rect 26068 18272 26096 19110
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26016 18244 26096 18272
rect 25964 18226 26016 18232
rect 25872 18148 25924 18154
rect 25872 18090 25924 18096
rect 25884 16998 25912 18090
rect 25976 17270 26004 18226
rect 26620 18222 26648 18702
rect 26608 18216 26660 18222
rect 26608 18158 26660 18164
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26332 17332 26384 17338
rect 26528 17320 26556 17478
rect 26384 17292 26556 17320
rect 26332 17274 26384 17280
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 25884 15910 25912 16526
rect 25872 15904 25924 15910
rect 25872 15846 25924 15852
rect 25688 15496 25740 15502
rect 25688 15438 25740 15444
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25424 14074 25452 14758
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25516 13938 25544 14962
rect 25596 14884 25648 14890
rect 25780 14884 25832 14890
rect 25648 14844 25780 14872
rect 25596 14826 25648 14832
rect 25780 14826 25832 14832
rect 25872 14816 25924 14822
rect 25792 14764 25872 14770
rect 25792 14758 25924 14764
rect 25792 14742 25912 14758
rect 25688 14612 25740 14618
rect 25688 14554 25740 14560
rect 25700 14346 25728 14554
rect 25688 14340 25740 14346
rect 25688 14282 25740 14288
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25240 12260 25360 12288
rect 25240 11762 25268 12260
rect 25320 12164 25372 12170
rect 25320 12106 25372 12112
rect 25332 11898 25360 12106
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25424 11812 25452 12582
rect 25516 12152 25544 13874
rect 25792 13870 25820 14742
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25596 12164 25648 12170
rect 25516 12124 25596 12152
rect 25596 12106 25648 12112
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25596 11824 25648 11830
rect 25424 11784 25596 11812
rect 25596 11766 25648 11772
rect 25700 11762 25728 12038
rect 25228 11756 25280 11762
rect 25228 11698 25280 11704
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24872 10266 24900 10406
rect 25240 10266 25268 11494
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25332 10674 25360 10950
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 24780 10118 24900 10146
rect 24872 9994 24900 10118
rect 25332 10062 25360 10610
rect 25516 10606 25544 11086
rect 25504 10600 25556 10606
rect 25504 10542 25556 10548
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25516 9994 25544 10542
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25608 10266 25636 10406
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 25792 10062 25820 11086
rect 25884 10674 25912 13874
rect 25976 13802 26004 17206
rect 26528 16590 26556 17292
rect 26700 17332 26752 17338
rect 26700 17274 26752 17280
rect 26712 17202 26740 17274
rect 26608 17196 26660 17202
rect 26608 17138 26660 17144
rect 26700 17196 26752 17202
rect 26700 17138 26752 17144
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26160 15094 26188 16390
rect 26148 15088 26200 15094
rect 26148 15030 26200 15036
rect 26160 14770 26188 15030
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26068 14742 26188 14770
rect 26068 14618 26096 14742
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 26344 14074 26372 14894
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26436 13938 26464 16390
rect 26528 15434 26556 16526
rect 26620 15706 26648 17138
rect 26896 16114 26924 19110
rect 27080 18630 27108 19306
rect 27264 19242 27292 19306
rect 27252 19236 27304 19242
rect 27252 19178 27304 19184
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26884 16108 26936 16114
rect 26884 16050 26936 16056
rect 26608 15700 26660 15706
rect 26608 15642 26660 15648
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26528 14822 26556 15370
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26804 15094 26832 15302
rect 26792 15088 26844 15094
rect 26792 15030 26844 15036
rect 26516 14816 26568 14822
rect 26516 14758 26568 14764
rect 26804 14482 26832 15030
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26712 13938 26740 14214
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 25964 13796 26016 13802
rect 25964 13738 26016 13744
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 25976 12442 26004 12854
rect 26068 12714 26096 13670
rect 26804 12782 26832 14418
rect 26896 14113 26924 16050
rect 26976 15904 27028 15910
rect 26976 15846 27028 15852
rect 26988 15502 27016 15846
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 27080 15026 27108 18566
rect 27540 18290 27568 19858
rect 27632 19258 27660 22066
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27712 21616 27764 21622
rect 27712 21558 27764 21564
rect 27724 20602 27752 21558
rect 27816 21146 27844 21966
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 28000 21690 28028 21830
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27908 20466 27936 20742
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 28092 19446 28120 22986
rect 28276 22094 28304 22986
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 28368 22778 28396 22918
rect 28356 22772 28408 22778
rect 28356 22714 28408 22720
rect 29104 22642 29132 23122
rect 29184 22976 29236 22982
rect 29184 22918 29236 22924
rect 29092 22636 29144 22642
rect 29092 22578 29144 22584
rect 28816 22568 28868 22574
rect 28816 22510 28868 22516
rect 28184 22066 28304 22094
rect 28184 22030 28212 22066
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28448 21888 28500 21894
rect 28448 21830 28500 21836
rect 28460 20874 28488 21830
rect 28828 21690 28856 22510
rect 28816 21684 28868 21690
rect 28816 21626 28868 21632
rect 28724 21344 28776 21350
rect 28724 21286 28776 21292
rect 28736 21146 28764 21286
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 28828 20942 28856 21626
rect 29196 21554 29224 22918
rect 29288 22642 29316 24210
rect 29564 23322 29592 24550
rect 29932 24342 29960 25774
rect 30392 25294 30420 26200
rect 30472 26182 30524 26188
rect 30484 26042 30512 26182
rect 30472 26036 30524 26042
rect 30472 25978 30524 25984
rect 30576 25838 30604 27406
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 32956 27056 33008 27062
rect 32956 26998 33008 27004
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 31484 26784 31536 26790
rect 31484 26726 31536 26732
rect 31496 26382 31524 26726
rect 32416 26450 32444 26930
rect 32968 26450 32996 26998
rect 33784 26784 33836 26790
rect 33784 26726 33836 26732
rect 34060 26784 34112 26790
rect 34060 26726 34112 26732
rect 33046 26480 33102 26489
rect 32404 26444 32456 26450
rect 32404 26386 32456 26392
rect 32956 26444 33008 26450
rect 33046 26415 33048 26424
rect 32956 26386 33008 26392
rect 33100 26415 33102 26424
rect 33048 26386 33100 26392
rect 31484 26376 31536 26382
rect 31484 26318 31536 26324
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 32680 26376 32732 26382
rect 32864 26376 32916 26382
rect 32680 26318 32732 26324
rect 32784 26324 32864 26330
rect 32916 26324 33364 26330
rect 30748 26308 30800 26314
rect 30748 26250 30800 26256
rect 30932 26308 30984 26314
rect 30932 26250 30984 26256
rect 30564 25832 30616 25838
rect 30564 25774 30616 25780
rect 30656 25696 30708 25702
rect 30656 25638 30708 25644
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 29920 24336 29972 24342
rect 29920 24278 29972 24284
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 30208 23594 30236 24142
rect 30196 23588 30248 23594
rect 30196 23530 30248 23536
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 29368 23044 29420 23050
rect 29368 22986 29420 22992
rect 29380 22778 29408 22986
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 29276 22636 29328 22642
rect 29328 22596 29408 22624
rect 29276 22578 29328 22584
rect 29380 22234 29408 22596
rect 29368 22228 29420 22234
rect 29368 22170 29420 22176
rect 29460 21956 29512 21962
rect 29460 21898 29512 21904
rect 29472 21690 29500 21898
rect 29460 21684 29512 21690
rect 29460 21626 29512 21632
rect 29184 21548 29236 21554
rect 29184 21490 29236 21496
rect 29276 21480 29328 21486
rect 29276 21422 29328 21428
rect 29368 21480 29420 21486
rect 29368 21422 29420 21428
rect 29288 21146 29316 21422
rect 29380 21146 29408 21422
rect 29564 21146 29592 23258
rect 30392 22574 30420 25230
rect 30668 24818 30696 25638
rect 30760 25158 30788 26250
rect 30944 25430 30972 26250
rect 31208 26240 31260 26246
rect 31208 26182 31260 26188
rect 31220 25906 31248 26182
rect 31496 25906 31524 26318
rect 31772 26246 31800 26318
rect 32692 26246 32720 26318
rect 32784 26314 33364 26324
rect 32784 26308 33376 26314
rect 32784 26302 33324 26308
rect 31760 26240 31812 26246
rect 31760 26182 31812 26188
rect 32220 26240 32272 26246
rect 32220 26182 32272 26188
rect 32680 26240 32732 26246
rect 32680 26182 32732 26188
rect 31208 25900 31260 25906
rect 31208 25842 31260 25848
rect 31484 25900 31536 25906
rect 31484 25842 31536 25848
rect 31116 25832 31168 25838
rect 31116 25774 31168 25780
rect 30932 25424 30984 25430
rect 30932 25366 30984 25372
rect 30748 25152 30800 25158
rect 30748 25094 30800 25100
rect 30760 24954 30788 25094
rect 30748 24948 30800 24954
rect 30748 24890 30800 24896
rect 30944 24818 30972 25366
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30576 23662 30604 24346
rect 30564 23656 30616 23662
rect 30564 23598 30616 23604
rect 30472 23520 30524 23526
rect 30472 23462 30524 23468
rect 30484 22642 30512 23462
rect 30668 22778 30696 24754
rect 30944 24410 30972 24754
rect 31128 24750 31156 25774
rect 31208 25288 31260 25294
rect 31208 25230 31260 25236
rect 31220 24954 31248 25230
rect 31484 25220 31536 25226
rect 31484 25162 31536 25168
rect 31852 25220 31904 25226
rect 31852 25162 31904 25168
rect 31208 24948 31260 24954
rect 31208 24890 31260 24896
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 30932 24404 30984 24410
rect 30932 24346 30984 24352
rect 30932 23656 30984 23662
rect 30932 23598 30984 23604
rect 30944 23322 30972 23598
rect 31496 23322 31524 25162
rect 31760 25152 31812 25158
rect 31760 25094 31812 25100
rect 31772 24614 31800 25094
rect 31864 24886 31892 25162
rect 32128 25152 32180 25158
rect 32128 25094 32180 25100
rect 31852 24880 31904 24886
rect 31852 24822 31904 24828
rect 31864 24750 31892 24822
rect 31852 24744 31904 24750
rect 31852 24686 31904 24692
rect 31760 24608 31812 24614
rect 31760 24550 31812 24556
rect 31864 24274 31892 24686
rect 32140 24410 32168 25094
rect 32232 24954 32260 26182
rect 32312 25152 32364 25158
rect 32312 25094 32364 25100
rect 32324 24954 32352 25094
rect 32220 24948 32272 24954
rect 32220 24890 32272 24896
rect 32312 24948 32364 24954
rect 32312 24890 32364 24896
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32588 24812 32640 24818
rect 32588 24754 32640 24760
rect 32128 24404 32180 24410
rect 32128 24346 32180 24352
rect 31852 24268 31904 24274
rect 31852 24210 31904 24216
rect 32232 24206 32260 24754
rect 32508 24614 32536 24754
rect 32600 24682 32628 24754
rect 32588 24676 32640 24682
rect 32588 24618 32640 24624
rect 32496 24608 32548 24614
rect 32496 24550 32548 24556
rect 32508 24274 32536 24550
rect 32496 24268 32548 24274
rect 32496 24210 32548 24216
rect 32220 24200 32272 24206
rect 32220 24142 32272 24148
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 30932 23316 30984 23322
rect 30932 23258 30984 23264
rect 31484 23316 31536 23322
rect 31484 23258 31536 23264
rect 32232 23186 32260 24142
rect 32220 23180 32272 23186
rect 32220 23122 32272 23128
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 30656 22772 30708 22778
rect 30656 22714 30708 22720
rect 31036 22642 31064 22918
rect 30472 22636 30524 22642
rect 30472 22578 30524 22584
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 30380 22568 30432 22574
rect 30380 22510 30432 22516
rect 30392 22098 30420 22510
rect 31220 22234 31248 23054
rect 32232 22778 32260 23122
rect 32324 23118 32352 24142
rect 32600 24138 32628 24618
rect 32588 24132 32640 24138
rect 32588 24074 32640 24080
rect 32680 24064 32732 24070
rect 32680 24006 32732 24012
rect 32692 23866 32720 24006
rect 32680 23860 32732 23866
rect 32680 23802 32732 23808
rect 32784 23746 32812 26302
rect 33324 26250 33376 26256
rect 33796 25294 33824 26726
rect 34072 26586 34100 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 34060 26580 34112 26586
rect 34060 26522 34112 26528
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33324 25220 33376 25226
rect 33324 25162 33376 25168
rect 33336 24954 33364 25162
rect 33324 24948 33376 24954
rect 33324 24890 33376 24896
rect 33796 24818 33824 25230
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 33140 24404 33192 24410
rect 33140 24346 33192 24352
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32956 24200 33008 24206
rect 32956 24142 33008 24148
rect 32600 23718 32812 23746
rect 32600 23594 32628 23718
rect 32588 23588 32640 23594
rect 32588 23530 32640 23536
rect 32404 23180 32456 23186
rect 32404 23122 32456 23128
rect 32312 23112 32364 23118
rect 32312 23054 32364 23060
rect 32220 22772 32272 22778
rect 32220 22714 32272 22720
rect 32416 22438 32444 23122
rect 32600 22982 32628 23530
rect 32876 23322 32904 24142
rect 32968 23798 32996 24142
rect 33048 24064 33100 24070
rect 33048 24006 33100 24012
rect 32956 23792 33008 23798
rect 32956 23734 33008 23740
rect 33060 23662 33088 24006
rect 33048 23656 33100 23662
rect 33048 23598 33100 23604
rect 32864 23316 32916 23322
rect 32864 23258 32916 23264
rect 32956 23316 33008 23322
rect 32956 23258 33008 23264
rect 32876 23050 32904 23258
rect 32864 23044 32916 23050
rect 32864 22986 32916 22992
rect 32588 22976 32640 22982
rect 32588 22918 32640 22924
rect 32968 22574 32996 23258
rect 32956 22568 33008 22574
rect 32956 22510 33008 22516
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 32588 22432 32640 22438
rect 32588 22374 32640 22380
rect 31208 22228 31260 22234
rect 31208 22170 31260 22176
rect 30380 22092 30432 22098
rect 30380 22034 30432 22040
rect 32140 21962 32168 22374
rect 32416 22250 32444 22374
rect 32416 22234 32536 22250
rect 32416 22228 32548 22234
rect 32416 22222 32496 22228
rect 32496 22170 32548 22176
rect 32128 21956 32180 21962
rect 32128 21898 32180 21904
rect 31852 21888 31904 21894
rect 31852 21830 31904 21836
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30208 21146 30236 21286
rect 29276 21140 29328 21146
rect 29276 21082 29328 21088
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 29552 21140 29604 21146
rect 29552 21082 29604 21088
rect 30196 21140 30248 21146
rect 30196 21082 30248 21088
rect 29184 21072 29236 21078
rect 29184 21014 29236 21020
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28460 20534 28488 20810
rect 29196 20602 29224 21014
rect 29276 20800 29328 20806
rect 29276 20742 29328 20748
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 30472 20800 30524 20806
rect 30472 20742 30524 20748
rect 30564 20800 30616 20806
rect 30564 20742 30616 20748
rect 29184 20596 29236 20602
rect 29184 20538 29236 20544
rect 28448 20528 28500 20534
rect 28448 20470 28500 20476
rect 29288 20466 29316 20742
rect 30116 20466 30144 20742
rect 29276 20460 29328 20466
rect 29276 20402 29328 20408
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28540 20256 28592 20262
rect 28540 20198 28592 20204
rect 28552 20058 28580 20198
rect 28540 20052 28592 20058
rect 28540 19994 28592 20000
rect 28080 19440 28132 19446
rect 28080 19382 28132 19388
rect 27632 19230 27752 19258
rect 27724 19174 27752 19230
rect 27712 19168 27764 19174
rect 27712 19110 27764 19116
rect 27724 18834 27752 19110
rect 27712 18828 27764 18834
rect 27712 18770 27764 18776
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27632 17882 27660 18158
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27724 17134 27752 18770
rect 28092 18766 28120 19382
rect 28724 18896 28776 18902
rect 28724 18838 28776 18844
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 28736 18426 28764 18838
rect 28828 18834 28856 20334
rect 29092 20256 29144 20262
rect 29092 20198 29144 20204
rect 29104 20058 29132 20198
rect 29092 20052 29144 20058
rect 29092 19994 29144 20000
rect 29288 19854 29316 20402
rect 29368 20052 29420 20058
rect 29368 19994 29420 20000
rect 29380 19854 29408 19994
rect 29736 19984 29788 19990
rect 29736 19926 29788 19932
rect 29276 19848 29328 19854
rect 29276 19790 29328 19796
rect 29368 19848 29420 19854
rect 29368 19790 29420 19796
rect 29748 19514 29776 19926
rect 30116 19718 30144 20402
rect 30484 20330 30512 20742
rect 30576 20466 30604 20742
rect 30564 20460 30616 20466
rect 30564 20402 30616 20408
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 30472 20324 30524 20330
rect 30472 20266 30524 20272
rect 30484 20058 30512 20266
rect 30472 20052 30524 20058
rect 30472 19994 30524 20000
rect 30104 19712 30156 19718
rect 30104 19654 30156 19660
rect 30564 19712 30616 19718
rect 30564 19654 30616 19660
rect 29736 19508 29788 19514
rect 29736 19450 29788 19456
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 29932 18970 29960 19314
rect 30116 19310 30144 19654
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 29920 18964 29972 18970
rect 29920 18906 29972 18912
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29196 18426 29224 18702
rect 30300 18698 30328 19314
rect 30576 18902 30604 19654
rect 30656 19508 30708 19514
rect 30656 19450 30708 19456
rect 30564 18896 30616 18902
rect 30564 18838 30616 18844
rect 29644 18692 29696 18698
rect 29644 18634 29696 18640
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27896 17128 27948 17134
rect 27896 17070 27948 17076
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27158 16688 27214 16697
rect 27158 16623 27214 16632
rect 27172 15910 27200 16623
rect 27632 16590 27660 16934
rect 27908 16794 27936 17070
rect 27896 16788 27948 16794
rect 27896 16730 27948 16736
rect 28000 16658 28028 17614
rect 28276 17338 28304 17614
rect 28264 17332 28316 17338
rect 28264 17274 28316 17280
rect 29656 17202 29684 18634
rect 29736 18624 29788 18630
rect 29736 18566 29788 18572
rect 29748 17338 29776 18566
rect 30300 18426 30328 18634
rect 30288 18420 30340 18426
rect 30288 18362 30340 18368
rect 30300 17746 30328 18362
rect 30668 17746 30696 19450
rect 31404 19446 31432 20402
rect 31864 19514 31892 21830
rect 32036 21480 32088 21486
rect 32036 21422 32088 21428
rect 32048 20942 32076 21422
rect 32036 20936 32088 20942
rect 32036 20878 32088 20884
rect 32048 19854 32076 20878
rect 32128 20868 32180 20874
rect 32128 20810 32180 20816
rect 32140 20602 32168 20810
rect 32128 20596 32180 20602
rect 32128 20538 32180 20544
rect 32600 20346 32628 22374
rect 33048 21956 33100 21962
rect 33048 21898 33100 21904
rect 33060 21486 33088 21898
rect 33048 21480 33100 21486
rect 33048 21422 33100 21428
rect 33152 21078 33180 24346
rect 33888 23662 33916 26386
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 35532 25288 35584 25294
rect 35532 25230 35584 25236
rect 37280 25288 37332 25294
rect 37280 25230 37332 25236
rect 34336 24812 34388 24818
rect 34336 24754 34388 24760
rect 34520 24812 34572 24818
rect 34520 24754 34572 24760
rect 34348 24206 34376 24754
rect 34532 24410 34560 24754
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34520 24404 34572 24410
rect 34520 24346 34572 24352
rect 35544 24206 35572 25230
rect 36176 25152 36228 25158
rect 36176 25094 36228 25100
rect 36188 24886 36216 25094
rect 36176 24880 36228 24886
rect 36176 24822 36228 24828
rect 35992 24608 36044 24614
rect 35992 24550 36044 24556
rect 36084 24608 36136 24614
rect 36084 24550 36136 24556
rect 36004 24206 36032 24550
rect 34336 24200 34388 24206
rect 34336 24142 34388 24148
rect 35164 24200 35216 24206
rect 35164 24142 35216 24148
rect 35532 24200 35584 24206
rect 35532 24142 35584 24148
rect 35992 24200 36044 24206
rect 35992 24142 36044 24148
rect 34060 24132 34112 24138
rect 34060 24074 34112 24080
rect 33876 23656 33928 23662
rect 33876 23598 33928 23604
rect 34072 23594 34100 24074
rect 34152 23724 34204 23730
rect 34152 23666 34204 23672
rect 34060 23588 34112 23594
rect 34060 23530 34112 23536
rect 34164 23118 34192 23666
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 34152 23112 34204 23118
rect 34152 23054 34204 23060
rect 33244 22234 33272 23054
rect 34244 23044 34296 23050
rect 34244 22986 34296 22992
rect 34256 22778 34284 22986
rect 34244 22772 34296 22778
rect 34244 22714 34296 22720
rect 34348 22710 34376 24142
rect 35176 23866 35204 24142
rect 35164 23860 35216 23866
rect 35164 23802 35216 23808
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35544 23322 35572 24142
rect 36096 23662 36124 24550
rect 37292 24410 37320 25230
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 37924 24608 37976 24614
rect 37924 24550 37976 24556
rect 37936 24410 37964 24550
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 37280 24404 37332 24410
rect 37280 24346 37332 24352
rect 37924 24404 37976 24410
rect 37924 24346 37976 24352
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 37096 24200 37148 24206
rect 37096 24142 37148 24148
rect 36268 23792 36320 23798
rect 36268 23734 36320 23740
rect 36084 23656 36136 23662
rect 36084 23598 36136 23604
rect 35348 23316 35400 23322
rect 35348 23258 35400 23264
rect 35532 23316 35584 23322
rect 35532 23258 35584 23264
rect 34428 23112 34480 23118
rect 34428 23054 34480 23060
rect 33876 22704 33928 22710
rect 33876 22646 33928 22652
rect 34336 22704 34388 22710
rect 34336 22646 34388 22652
rect 33324 22636 33376 22642
rect 33324 22578 33376 22584
rect 33232 22228 33284 22234
rect 33232 22170 33284 22176
rect 33336 22030 33364 22578
rect 33888 22166 33916 22646
rect 33876 22160 33928 22166
rect 33876 22102 33928 22108
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 33888 21622 33916 22102
rect 34440 22098 34468 23054
rect 34520 22636 34572 22642
rect 34520 22578 34572 22584
rect 34532 22166 34560 22578
rect 35360 22506 35388 23258
rect 36096 23202 36124 23598
rect 36096 23174 36216 23202
rect 36188 23118 36216 23174
rect 36084 23112 36136 23118
rect 36084 23054 36136 23060
rect 36176 23112 36228 23118
rect 36176 23054 36228 23060
rect 35440 22976 35492 22982
rect 35440 22918 35492 22924
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35348 22500 35400 22506
rect 35348 22442 35400 22448
rect 35256 22432 35308 22438
rect 35308 22380 35388 22386
rect 35256 22374 35388 22380
rect 35268 22358 35388 22374
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34520 22160 34572 22166
rect 34520 22102 34572 22108
rect 34796 22160 34848 22166
rect 34796 22102 34848 22108
rect 34428 22092 34480 22098
rect 34428 22034 34480 22040
rect 34808 22030 34836 22102
rect 35164 22094 35216 22098
rect 35360 22094 35388 22358
rect 35164 22092 35388 22094
rect 35216 22066 35388 22092
rect 35164 22034 35216 22040
rect 35452 22030 35480 22918
rect 35544 22166 35572 22918
rect 36096 22778 36124 23054
rect 36084 22772 36136 22778
rect 36084 22714 36136 22720
rect 35624 22568 35676 22574
rect 35624 22510 35676 22516
rect 35532 22160 35584 22166
rect 35532 22102 35584 22108
rect 35636 22098 35664 22510
rect 35992 22432 36044 22438
rect 35992 22374 36044 22380
rect 35624 22092 35676 22098
rect 35624 22034 35676 22040
rect 35900 22092 35952 22098
rect 35900 22034 35952 22040
rect 34796 22024 34848 22030
rect 35440 22024 35492 22030
rect 34796 21966 34848 21972
rect 35360 21984 35440 22012
rect 35360 21690 35388 21984
rect 35440 21966 35492 21972
rect 35808 21888 35860 21894
rect 35808 21830 35860 21836
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 33876 21616 33928 21622
rect 33876 21558 33928 21564
rect 35440 21616 35492 21622
rect 35440 21558 35492 21564
rect 34244 21548 34296 21554
rect 34244 21490 34296 21496
rect 34256 21146 34284 21490
rect 35348 21344 35400 21350
rect 35348 21286 35400 21292
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34244 21140 34296 21146
rect 34244 21082 34296 21088
rect 33140 21072 33192 21078
rect 33140 21014 33192 21020
rect 33876 21072 33928 21078
rect 33876 21014 33928 21020
rect 33888 20942 33916 21014
rect 35360 21010 35388 21286
rect 35452 21010 35480 21558
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35348 21004 35400 21010
rect 35348 20946 35400 20952
rect 35440 21004 35492 21010
rect 35440 20946 35492 20952
rect 33876 20936 33928 20942
rect 33876 20878 33928 20884
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 32864 20800 32916 20806
rect 32864 20742 32916 20748
rect 35072 20800 35124 20806
rect 35072 20742 35124 20748
rect 32876 20466 32904 20742
rect 33140 20528 33192 20534
rect 33140 20470 33192 20476
rect 32864 20460 32916 20466
rect 32864 20402 32916 20408
rect 32600 20318 32812 20346
rect 32036 19848 32088 19854
rect 32036 19790 32088 19796
rect 31852 19508 31904 19514
rect 31852 19450 31904 19456
rect 31392 19440 31444 19446
rect 31392 19382 31444 19388
rect 31668 19440 31720 19446
rect 31668 19382 31720 19388
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30760 18834 30788 19110
rect 31404 18970 31432 19382
rect 31680 19334 31708 19382
rect 31944 19372 31996 19378
rect 31680 19306 31800 19334
rect 31944 19314 31996 19320
rect 31772 18970 31800 19306
rect 31392 18964 31444 18970
rect 31392 18906 31444 18912
rect 31760 18964 31812 18970
rect 31760 18906 31812 18912
rect 30840 18896 30892 18902
rect 30840 18838 30892 18844
rect 30748 18828 30800 18834
rect 30748 18770 30800 18776
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30656 17740 30708 17746
rect 30656 17682 30708 17688
rect 29828 17536 29880 17542
rect 29828 17478 29880 17484
rect 29840 17338 29868 17478
rect 29736 17332 29788 17338
rect 29736 17274 29788 17280
rect 29828 17332 29880 17338
rect 29828 17274 29880 17280
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 28264 16992 28316 16998
rect 28264 16934 28316 16940
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27434 15056 27490 15065
rect 27068 15020 27120 15026
rect 27540 15042 27568 15302
rect 27490 15026 27568 15042
rect 27632 15026 27660 16526
rect 27816 16250 27844 16526
rect 27804 16244 27856 16250
rect 27804 16186 27856 16192
rect 27816 15706 27844 16186
rect 28000 16182 28028 16594
rect 27988 16176 28040 16182
rect 27988 16118 28040 16124
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 27804 15496 27856 15502
rect 27804 15438 27856 15444
rect 27490 15020 27580 15026
rect 27490 15014 27528 15020
rect 27434 14991 27490 15000
rect 27068 14962 27120 14968
rect 27528 14962 27580 14968
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27816 14822 27844 15438
rect 28000 15026 28028 16118
rect 28276 16114 28304 16934
rect 30668 16794 30696 17682
rect 30852 17678 30880 18838
rect 31668 18828 31720 18834
rect 31668 18770 31720 18776
rect 31208 18216 31260 18222
rect 31208 18158 31260 18164
rect 31024 18080 31076 18086
rect 31024 18022 31076 18028
rect 31036 17678 31064 18022
rect 31220 17882 31248 18158
rect 31208 17876 31260 17882
rect 31208 17818 31260 17824
rect 30748 17672 30800 17678
rect 30748 17614 30800 17620
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 31484 17672 31536 17678
rect 31484 17614 31536 17620
rect 30760 17134 30788 17614
rect 30748 17128 30800 17134
rect 30748 17070 30800 17076
rect 31496 16794 31524 17614
rect 30656 16788 30708 16794
rect 30656 16730 30708 16736
rect 31484 16788 31536 16794
rect 31484 16730 31536 16736
rect 30668 16640 30696 16730
rect 30668 16612 30788 16640
rect 29920 16584 29972 16590
rect 29920 16526 29972 16532
rect 30104 16584 30156 16590
rect 30104 16526 30156 16532
rect 28540 16516 28592 16522
rect 28540 16458 28592 16464
rect 28552 16250 28580 16458
rect 29828 16448 29880 16454
rect 29828 16390 29880 16396
rect 28540 16244 28592 16250
rect 28540 16186 28592 16192
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 29840 16046 29868 16390
rect 29932 16250 29960 16526
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 29828 16040 29880 16046
rect 29828 15982 29880 15988
rect 29840 15502 29868 15982
rect 29932 15706 29960 16186
rect 30116 16182 30144 16526
rect 30760 16522 30788 16612
rect 30748 16516 30800 16522
rect 30748 16458 30800 16464
rect 30840 16448 30892 16454
rect 30840 16390 30892 16396
rect 30104 16176 30156 16182
rect 30104 16118 30156 16124
rect 29920 15700 29972 15706
rect 29920 15642 29972 15648
rect 30116 15570 30144 16118
rect 30852 16046 30880 16390
rect 31496 16046 31524 16730
rect 31680 16574 31708 18770
rect 31956 18290 31984 19314
rect 32600 18834 32628 20318
rect 32680 20256 32732 20262
rect 32680 20198 32732 20204
rect 32692 19378 32720 20198
rect 32784 20058 32812 20318
rect 32864 20256 32916 20262
rect 32864 20198 32916 20204
rect 32772 20052 32824 20058
rect 32772 19994 32824 20000
rect 32876 19786 32904 20198
rect 32864 19780 32916 19786
rect 32864 19722 32916 19728
rect 32956 19780 33008 19786
rect 32956 19722 33008 19728
rect 32772 19712 32824 19718
rect 32772 19654 32824 19660
rect 32784 19514 32812 19654
rect 32968 19514 32996 19722
rect 32772 19508 32824 19514
rect 32772 19450 32824 19456
rect 32956 19508 33008 19514
rect 32956 19450 33008 19456
rect 32680 19372 32732 19378
rect 32680 19314 32732 19320
rect 32680 19168 32732 19174
rect 32680 19110 32732 19116
rect 32588 18828 32640 18834
rect 32588 18770 32640 18776
rect 32692 18766 32720 19110
rect 32968 18834 32996 19450
rect 33152 19378 33180 20470
rect 35084 20466 35112 20742
rect 35360 20602 35388 20810
rect 35452 20602 35480 20946
rect 35728 20874 35756 21286
rect 35532 20868 35584 20874
rect 35532 20810 35584 20816
rect 35716 20868 35768 20874
rect 35716 20810 35768 20816
rect 35348 20596 35400 20602
rect 35348 20538 35400 20544
rect 35440 20596 35492 20602
rect 35440 20538 35492 20544
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 35072 20460 35124 20466
rect 35072 20402 35124 20408
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 33692 20256 33744 20262
rect 33692 20198 33744 20204
rect 33704 19786 33732 20198
rect 33692 19780 33744 19786
rect 33692 19722 33744 19728
rect 33416 19712 33468 19718
rect 33416 19654 33468 19660
rect 33428 19446 33456 19654
rect 34532 19446 34560 20402
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20058 35388 20402
rect 35452 20058 35480 20538
rect 35544 20466 35572 20810
rect 35624 20528 35676 20534
rect 35624 20470 35676 20476
rect 35532 20460 35584 20466
rect 35532 20402 35584 20408
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 35440 20052 35492 20058
rect 35440 19994 35492 20000
rect 35256 19916 35308 19922
rect 35256 19858 35308 19864
rect 34612 19780 34664 19786
rect 34612 19722 34664 19728
rect 33416 19440 33468 19446
rect 33416 19382 33468 19388
rect 34520 19440 34572 19446
rect 34520 19382 34572 19388
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 34624 19310 34652 19722
rect 34888 19712 34940 19718
rect 35164 19712 35216 19718
rect 34888 19654 34940 19660
rect 35084 19660 35164 19666
rect 35084 19654 35216 19660
rect 34612 19304 34664 19310
rect 34612 19246 34664 19252
rect 34624 18970 34652 19246
rect 34900 19174 34928 19654
rect 35084 19638 35204 19654
rect 35084 19446 35112 19638
rect 35268 19446 35296 19858
rect 35636 19802 35664 20470
rect 35820 20466 35848 21830
rect 35912 21146 35940 22034
rect 36004 21962 36032 22374
rect 36188 22234 36216 23054
rect 36280 23050 36308 23734
rect 36372 23730 36400 24142
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36360 23588 36412 23594
rect 36360 23530 36412 23536
rect 36268 23044 36320 23050
rect 36268 22986 36320 22992
rect 36176 22228 36228 22234
rect 36176 22170 36228 22176
rect 35992 21956 36044 21962
rect 35992 21898 36044 21904
rect 36268 21888 36320 21894
rect 36268 21830 36320 21836
rect 36280 21690 36308 21830
rect 36268 21684 36320 21690
rect 36268 21626 36320 21632
rect 35900 21140 35952 21146
rect 35900 21082 35952 21088
rect 35808 20460 35860 20466
rect 35808 20402 35860 20408
rect 36084 20460 36136 20466
rect 36084 20402 36136 20408
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 35900 20256 35952 20262
rect 35900 20198 35952 20204
rect 35912 19854 35940 20198
rect 36096 20058 36124 20402
rect 36084 20052 36136 20058
rect 36084 19994 36136 20000
rect 36188 19922 36216 20402
rect 36176 19916 36228 19922
rect 36176 19858 36228 19864
rect 35544 19774 35664 19802
rect 35900 19848 35952 19854
rect 35900 19790 35952 19796
rect 35544 19718 35572 19774
rect 35532 19712 35584 19718
rect 35532 19654 35584 19660
rect 35624 19712 35676 19718
rect 35624 19654 35676 19660
rect 35072 19440 35124 19446
rect 35072 19382 35124 19388
rect 35256 19440 35308 19446
rect 35636 19394 35664 19654
rect 35256 19382 35308 19388
rect 35084 19310 35112 19382
rect 35544 19378 35664 19394
rect 35532 19372 35664 19378
rect 35584 19366 35664 19372
rect 35532 19314 35584 19320
rect 35072 19304 35124 19310
rect 35072 19246 35124 19252
rect 34796 19168 34848 19174
rect 34796 19110 34848 19116
rect 34888 19168 34940 19174
rect 34888 19110 34940 19116
rect 33968 18964 34020 18970
rect 33968 18906 34020 18912
rect 34612 18964 34664 18970
rect 34612 18906 34664 18912
rect 32956 18828 33008 18834
rect 32956 18770 33008 18776
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 31944 18284 31996 18290
rect 31944 18226 31996 18232
rect 33980 17814 34008 18906
rect 34808 18766 34836 19110
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34980 18896 35032 18902
rect 34980 18838 35032 18844
rect 34796 18760 34848 18766
rect 34796 18702 34848 18708
rect 34992 18358 35020 18838
rect 34980 18352 35032 18358
rect 34980 18294 35032 18300
rect 35348 18284 35400 18290
rect 35348 18226 35400 18232
rect 34796 18080 34848 18086
rect 34796 18022 34848 18028
rect 33968 17808 34020 17814
rect 33968 17750 34020 17756
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 33796 17270 33824 17478
rect 33980 17270 34008 17750
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 33784 17264 33836 17270
rect 33784 17206 33836 17212
rect 33968 17264 34020 17270
rect 33968 17206 34020 17212
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 31864 16658 31892 17138
rect 34532 17134 34560 17614
rect 34704 17536 34756 17542
rect 34704 17478 34756 17484
rect 34716 17338 34744 17478
rect 34808 17338 34836 18022
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17882 35388 18226
rect 35912 17882 35940 19790
rect 36372 18290 36400 23530
rect 36464 23186 36492 24006
rect 37108 23730 37136 24142
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 36544 23724 36596 23730
rect 36544 23666 36596 23672
rect 37096 23724 37148 23730
rect 37096 23666 37148 23672
rect 36556 23254 36584 23666
rect 36728 23656 36780 23662
rect 36728 23598 36780 23604
rect 36820 23656 36872 23662
rect 36820 23598 36872 23604
rect 36636 23588 36688 23594
rect 36636 23530 36688 23536
rect 36648 23322 36676 23530
rect 36636 23316 36688 23322
rect 36636 23258 36688 23264
rect 36544 23248 36596 23254
rect 36544 23190 36596 23196
rect 36452 23180 36504 23186
rect 36452 23122 36504 23128
rect 36556 22166 36584 23190
rect 36740 23186 36768 23598
rect 36728 23180 36780 23186
rect 36728 23122 36780 23128
rect 36636 23112 36688 23118
rect 36636 23054 36688 23060
rect 36544 22160 36596 22166
rect 36544 22102 36596 22108
rect 36556 21842 36584 22102
rect 36648 22098 36676 23054
rect 36636 22092 36688 22098
rect 36740 22094 36768 23122
rect 36832 22930 36860 23598
rect 37280 23520 37332 23526
rect 37280 23462 37332 23468
rect 37292 23118 37320 23462
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 37280 23112 37332 23118
rect 37280 23054 37332 23060
rect 38384 22976 38436 22982
rect 36832 22902 37044 22930
rect 38384 22918 38436 22924
rect 36740 22066 36860 22094
rect 36636 22034 36688 22040
rect 36728 22024 36780 22030
rect 36728 21966 36780 21972
rect 36556 21814 36676 21842
rect 36648 21554 36676 21814
rect 36740 21622 36768 21966
rect 36832 21894 36860 22066
rect 36912 21956 36964 21962
rect 36912 21898 36964 21904
rect 36820 21888 36872 21894
rect 36820 21830 36872 21836
rect 36728 21616 36780 21622
rect 36728 21558 36780 21564
rect 36636 21548 36688 21554
rect 36636 21490 36688 21496
rect 36924 21418 36952 21898
rect 36912 21412 36964 21418
rect 36912 21354 36964 21360
rect 36728 20460 36780 20466
rect 36728 20402 36780 20408
rect 36740 18902 36768 20402
rect 37016 19922 37044 22902
rect 38396 22778 38424 22918
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 38384 22772 38436 22778
rect 38384 22714 38436 22720
rect 38016 22704 38068 22710
rect 38016 22646 38068 22652
rect 38028 22234 38056 22646
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 38016 22228 38068 22234
rect 38016 22170 38068 22176
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 37188 20936 37240 20942
rect 37188 20878 37240 20884
rect 38660 20936 38712 20942
rect 38660 20878 38712 20884
rect 37200 20602 37228 20878
rect 37832 20800 37884 20806
rect 37832 20742 37884 20748
rect 37924 20800 37976 20806
rect 37924 20742 37976 20748
rect 37188 20596 37240 20602
rect 37188 20538 37240 20544
rect 37844 20534 37872 20742
rect 37832 20528 37884 20534
rect 37832 20470 37884 20476
rect 37936 20466 37964 20742
rect 38672 20602 38700 20878
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 38660 20596 38712 20602
rect 38660 20538 38712 20544
rect 37924 20460 37976 20466
rect 37924 20402 37976 20408
rect 37280 20392 37332 20398
rect 37280 20334 37332 20340
rect 37188 20256 37240 20262
rect 37188 20198 37240 20204
rect 37200 20058 37228 20198
rect 37188 20052 37240 20058
rect 37188 19994 37240 20000
rect 37004 19916 37056 19922
rect 37004 19858 37056 19864
rect 37016 19802 37044 19858
rect 37016 19774 37136 19802
rect 37004 19712 37056 19718
rect 37004 19654 37056 19660
rect 37016 19514 37044 19654
rect 37004 19508 37056 19514
rect 37004 19450 37056 19456
rect 36728 18896 36780 18902
rect 36728 18838 36780 18844
rect 36636 18624 36688 18630
rect 36636 18566 36688 18572
rect 36648 18358 36676 18566
rect 36740 18426 36768 18838
rect 37004 18624 37056 18630
rect 37004 18566 37056 18572
rect 37016 18426 37044 18566
rect 36728 18420 36780 18426
rect 36728 18362 36780 18368
rect 37004 18420 37056 18426
rect 37004 18362 37056 18368
rect 36636 18352 36688 18358
rect 36636 18294 36688 18300
rect 36084 18284 36136 18290
rect 36084 18226 36136 18232
rect 36360 18284 36412 18290
rect 36360 18226 36412 18232
rect 36452 18284 36504 18290
rect 36452 18226 36504 18232
rect 36728 18284 36780 18290
rect 36728 18226 36780 18232
rect 36912 18284 36964 18290
rect 36912 18226 36964 18232
rect 35348 17876 35400 17882
rect 35348 17818 35400 17824
rect 35900 17876 35952 17882
rect 35900 17818 35952 17824
rect 36096 17814 36124 18226
rect 36084 17808 36136 17814
rect 36084 17750 36136 17756
rect 36464 17678 36492 18226
rect 36452 17672 36504 17678
rect 36452 17614 36504 17620
rect 36740 17610 36768 18226
rect 36924 17678 36952 18226
rect 36820 17672 36872 17678
rect 36820 17614 36872 17620
rect 36912 17672 36964 17678
rect 36912 17614 36964 17620
rect 36728 17604 36780 17610
rect 36728 17546 36780 17552
rect 36832 17338 36860 17614
rect 34612 17332 34664 17338
rect 34612 17274 34664 17280
rect 34704 17332 34756 17338
rect 34704 17274 34756 17280
rect 34796 17332 34848 17338
rect 34796 17274 34848 17280
rect 36820 17332 36872 17338
rect 36820 17274 36872 17280
rect 34520 17128 34572 17134
rect 34520 17070 34572 17076
rect 33416 16992 33468 16998
rect 33416 16934 33468 16940
rect 31852 16652 31904 16658
rect 31852 16594 31904 16600
rect 31680 16546 31800 16574
rect 31772 16114 31800 16546
rect 31760 16108 31812 16114
rect 31760 16050 31812 16056
rect 30840 16040 30892 16046
rect 30840 15982 30892 15988
rect 31484 16040 31536 16046
rect 31484 15982 31536 15988
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30760 15570 30788 15846
rect 30852 15638 30880 15982
rect 30840 15632 30892 15638
rect 30840 15574 30892 15580
rect 30104 15564 30156 15570
rect 30104 15506 30156 15512
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 28448 15360 28500 15366
rect 28448 15302 28500 15308
rect 29552 15360 29604 15366
rect 29552 15302 29604 15308
rect 29920 15360 29972 15366
rect 29920 15302 29972 15308
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27804 14816 27856 14822
rect 27804 14758 27856 14764
rect 27448 14618 27476 14758
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 28184 14550 28212 14962
rect 27620 14544 27672 14550
rect 27620 14486 27672 14492
rect 28172 14544 28224 14550
rect 28172 14486 28224 14492
rect 27344 14476 27396 14482
rect 27344 14418 27396 14424
rect 26882 14104 26938 14113
rect 26882 14039 26938 14048
rect 27356 13954 27384 14418
rect 27632 14346 27660 14486
rect 28460 14414 28488 15302
rect 29564 15094 29592 15302
rect 29552 15088 29604 15094
rect 29552 15030 29604 15036
rect 28448 14408 28500 14414
rect 28448 14350 28500 14356
rect 27620 14340 27672 14346
rect 27620 14282 27672 14288
rect 27264 13938 27384 13954
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 27252 13932 27384 13938
rect 27304 13926 27384 13932
rect 27252 13874 27304 13880
rect 26988 13394 27016 13874
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 27632 13326 27660 14282
rect 29552 14272 29604 14278
rect 29552 14214 29604 14220
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29564 14006 29592 14214
rect 29656 14074 29684 14214
rect 29644 14068 29696 14074
rect 29644 14010 29696 14016
rect 29552 14000 29604 14006
rect 29552 13942 29604 13948
rect 28356 13728 28408 13734
rect 28356 13670 28408 13676
rect 28368 13394 28396 13670
rect 29092 13456 29144 13462
rect 29092 13398 29144 13404
rect 28356 13388 28408 13394
rect 28356 13330 28408 13336
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26056 12708 26108 12714
rect 26056 12650 26108 12656
rect 25964 12436 26016 12442
rect 25964 12378 26016 12384
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25976 11354 26004 11562
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 25964 11008 26016 11014
rect 25964 10950 26016 10956
rect 25976 10674 26004 10950
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 26056 10056 26108 10062
rect 26160 10010 26188 12718
rect 26700 12436 26752 12442
rect 27632 12434 27660 13262
rect 28172 13184 28224 13190
rect 28172 13126 28224 13132
rect 27632 12406 27752 12434
rect 26700 12378 26752 12384
rect 26712 10742 26740 12378
rect 27252 12300 27304 12306
rect 27252 12242 27304 12248
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26804 11286 26832 11834
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 26792 11280 26844 11286
rect 26792 11222 26844 11228
rect 26700 10736 26752 10742
rect 26700 10678 26752 10684
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26424 10464 26476 10470
rect 26424 10406 26476 10412
rect 26108 10004 26188 10010
rect 26056 9998 26188 10004
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24952 9988 25004 9994
rect 24952 9930 25004 9936
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 22480 9178 22600 9194
rect 22468 9172 22600 9178
rect 22520 9166 22600 9172
rect 22468 9114 22520 9120
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 23124 9042 23152 9318
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21192 7478 21220 7686
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21836 6798 21864 7822
rect 21928 7274 21956 8434
rect 22020 7546 22048 8978
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 22664 8634 22692 8842
rect 23676 8634 23704 8842
rect 23860 8634 23888 9930
rect 24964 9722 24992 9930
rect 25148 9874 25176 9930
rect 25056 9846 25176 9874
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24412 9178 24440 9454
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22756 7886 22784 8434
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 22848 7478 22876 7686
rect 23676 7546 23704 7686
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22836 7472 22888 7478
rect 22836 7414 22888 7420
rect 21916 7268 21968 7274
rect 21916 7210 21968 7216
rect 22204 6866 22232 7414
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23584 6458 23612 6734
rect 23860 6458 23888 8570
rect 24688 8430 24716 9318
rect 24780 9178 24808 9522
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24964 8566 24992 9522
rect 25056 9382 25084 9846
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25056 8634 25084 9318
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 24952 8560 25004 8566
rect 24952 8502 25004 8508
rect 24964 8430 24992 8502
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24952 8424 25004 8430
rect 25240 8378 25268 9658
rect 25320 9036 25372 9042
rect 25516 9024 25544 9930
rect 25608 9178 25636 9998
rect 25700 9722 25728 9998
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25792 9586 25820 9998
rect 26068 9982 26188 9998
rect 26344 9926 26372 10406
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26240 9648 26292 9654
rect 26240 9590 26292 9596
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 25884 9178 25912 9522
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25372 8996 25544 9024
rect 25320 8978 25372 8984
rect 25332 8498 25360 8978
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 24952 8366 25004 8372
rect 24136 7886 24164 8366
rect 25056 8350 25636 8378
rect 25884 8362 25912 9114
rect 25976 8974 26004 9454
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24136 7546 24164 7822
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24136 7274 24164 7482
rect 24780 7478 24808 7958
rect 24768 7472 24820 7478
rect 25056 7426 25084 8350
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25148 7886 25176 8230
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 24768 7414 24820 7420
rect 24964 7410 25084 7426
rect 25240 7410 25268 8230
rect 25608 7818 25636 8350
rect 25872 8356 25924 8362
rect 25872 8298 25924 8304
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 25884 7410 25912 8298
rect 25964 8288 26016 8294
rect 25964 8230 26016 8236
rect 25976 7478 26004 8230
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 26148 7880 26200 7886
rect 26252 7868 26280 9590
rect 26344 9382 26372 9862
rect 26436 9654 26464 10406
rect 26528 10266 26556 10610
rect 26712 10606 26740 10678
rect 27172 10674 27200 11698
rect 27264 11218 27292 12242
rect 27724 12238 27752 12406
rect 27712 12232 27764 12238
rect 27712 12174 27764 12180
rect 28184 11898 28212 13126
rect 29104 12918 29132 13398
rect 29932 13326 29960 15302
rect 30024 15162 30052 15438
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 30116 13190 30144 15506
rect 30760 14958 30788 15506
rect 31496 15502 31524 15982
rect 31300 15496 31352 15502
rect 31300 15438 31352 15444
rect 31484 15496 31536 15502
rect 31484 15438 31536 15444
rect 30932 15360 30984 15366
rect 30932 15302 30984 15308
rect 30944 15162 30972 15302
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 31312 14958 31340 15438
rect 31772 15094 31800 16050
rect 31760 15088 31812 15094
rect 31760 15030 31812 15036
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 31300 14952 31352 14958
rect 31300 14894 31352 14900
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 30840 14816 30892 14822
rect 30840 14758 30892 14764
rect 30380 14408 30432 14414
rect 30380 14350 30432 14356
rect 30392 13530 30420 14350
rect 30564 13796 30616 13802
rect 30564 13738 30616 13744
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30576 13326 30604 13738
rect 30668 13530 30696 14758
rect 30852 14618 30880 14758
rect 30840 14612 30892 14618
rect 30840 14554 30892 14560
rect 31208 13864 31260 13870
rect 31208 13806 31260 13812
rect 31024 13728 31076 13734
rect 31024 13670 31076 13676
rect 31036 13530 31064 13670
rect 30656 13524 30708 13530
rect 30656 13466 30708 13472
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 30564 13320 30616 13326
rect 30564 13262 30616 13268
rect 30104 13184 30156 13190
rect 30104 13126 30156 13132
rect 30668 12918 30696 13466
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 28356 12912 28408 12918
rect 28356 12854 28408 12860
rect 29092 12912 29144 12918
rect 29092 12854 29144 12860
rect 30656 12912 30708 12918
rect 30656 12854 30708 12860
rect 28264 12640 28316 12646
rect 28264 12582 28316 12588
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 28080 11688 28132 11694
rect 28080 11630 28132 11636
rect 27252 11212 27304 11218
rect 27252 11154 27304 11160
rect 28092 10674 28120 11630
rect 28276 11014 28304 12582
rect 28264 11008 28316 11014
rect 28264 10950 28316 10956
rect 28276 10742 28304 10950
rect 28368 10810 28396 12854
rect 30944 12850 30972 13262
rect 31220 12850 31248 13806
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 28540 12776 28592 12782
rect 28540 12718 28592 12724
rect 29092 12776 29144 12782
rect 29092 12718 29144 12724
rect 28552 12646 28580 12718
rect 28540 12640 28592 12646
rect 28540 12582 28592 12588
rect 28552 12238 28580 12582
rect 29104 12434 29132 12718
rect 29184 12640 29236 12646
rect 29184 12582 29236 12588
rect 29012 12406 29132 12434
rect 29012 12306 29040 12406
rect 29000 12300 29052 12306
rect 29000 12242 29052 12248
rect 28540 12232 28592 12238
rect 28540 12174 28592 12180
rect 29012 11762 29040 12242
rect 29092 12232 29144 12238
rect 29196 12220 29224 12582
rect 30392 12442 30420 12786
rect 30656 12640 30708 12646
rect 30656 12582 30708 12588
rect 30380 12436 30432 12442
rect 30380 12378 30432 12384
rect 29144 12192 29224 12220
rect 29092 12174 29144 12180
rect 30012 11824 30064 11830
rect 30012 11766 30064 11772
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 28816 11688 28868 11694
rect 28816 11630 28868 11636
rect 28828 11354 28856 11630
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28172 10736 28224 10742
rect 28172 10678 28224 10684
rect 28264 10736 28316 10742
rect 28264 10678 28316 10684
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 26700 10600 26752 10606
rect 26700 10542 26752 10548
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 26712 9722 26740 9998
rect 27816 9722 27844 10406
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 27804 9716 27856 9722
rect 27804 9658 27856 9664
rect 26424 9648 26476 9654
rect 26424 9590 26476 9596
rect 27816 9602 27844 9658
rect 27160 9580 27212 9586
rect 27816 9574 27936 9602
rect 27160 9522 27212 9528
rect 26424 9512 26476 9518
rect 26424 9454 26476 9460
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26436 9178 26464 9454
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26528 9178 26556 9318
rect 27172 9178 27200 9522
rect 27804 9512 27856 9518
rect 27804 9454 27856 9460
rect 27436 9376 27488 9382
rect 27436 9318 27488 9324
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 26516 9172 26568 9178
rect 26516 9114 26568 9120
rect 27160 9172 27212 9178
rect 27160 9114 27212 9120
rect 26528 8974 26556 9114
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 26200 7840 26280 7868
rect 26148 7822 26200 7828
rect 26068 7546 26096 7822
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 25964 7472 26016 7478
rect 25964 7414 26016 7420
rect 24952 7404 25084 7410
rect 25004 7398 25084 7404
rect 25228 7404 25280 7410
rect 24952 7346 25004 7352
rect 25228 7346 25280 7352
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 26528 7342 26556 8910
rect 27172 8430 27200 9114
rect 27344 8900 27396 8906
rect 27344 8842 27396 8848
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27264 8566 27292 8774
rect 27252 8560 27304 8566
rect 27252 8502 27304 8508
rect 27160 8424 27212 8430
rect 27080 8372 27160 8378
rect 27080 8366 27212 8372
rect 27080 8350 27200 8366
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26516 7336 26568 7342
rect 26516 7278 26568 7284
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 24216 7268 24268 7274
rect 24216 7210 24268 7216
rect 24228 6866 24256 7210
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24412 7002 24440 7142
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 26528 6730 26556 7278
rect 26620 6730 26648 7822
rect 27080 7342 27108 8350
rect 27356 8294 27384 8842
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 27160 7540 27212 7546
rect 27160 7482 27212 7488
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27172 6798 27200 7482
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27356 7002 27384 7346
rect 27344 6996 27396 7002
rect 27344 6938 27396 6944
rect 27448 6866 27476 9318
rect 27816 9178 27844 9454
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27528 8900 27580 8906
rect 27528 8842 27580 8848
rect 27540 7886 27568 8842
rect 27908 7886 27936 9574
rect 28184 8498 28212 10678
rect 29012 10674 29040 11698
rect 30024 11354 30052 11766
rect 30668 11694 30696 12582
rect 30944 12238 30972 12786
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 30748 12164 30800 12170
rect 30748 12106 30800 12112
rect 30760 11898 30788 12106
rect 31116 12096 31168 12102
rect 31116 12038 31168 12044
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 31024 11552 31076 11558
rect 31024 11494 31076 11500
rect 30012 11348 30064 11354
rect 30012 11290 30064 11296
rect 30300 11218 30328 11494
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 29276 11008 29328 11014
rect 29276 10950 29328 10956
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 28816 9920 28868 9926
rect 28816 9862 28868 9868
rect 28828 9654 28856 9862
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 29012 9518 29040 10610
rect 29288 10062 29316 10950
rect 31036 10742 31064 11494
rect 30472 10736 30524 10742
rect 30472 10678 30524 10684
rect 31024 10736 31076 10742
rect 31024 10678 31076 10684
rect 30484 10266 30512 10678
rect 30472 10260 30524 10266
rect 30472 10202 30524 10208
rect 31128 10062 31156 12038
rect 31220 11150 31248 12174
rect 31300 12096 31352 12102
rect 31300 12038 31352 12044
rect 31312 11898 31340 12038
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 31300 11756 31352 11762
rect 31300 11698 31352 11704
rect 31312 11354 31340 11698
rect 31404 11694 31432 12582
rect 31864 12186 31892 16594
rect 33428 16114 33456 16934
rect 34532 16658 34560 17070
rect 34520 16652 34572 16658
rect 34520 16594 34572 16600
rect 34624 16114 34652 17274
rect 36832 17134 36860 17274
rect 37108 17270 37136 19774
rect 37292 19378 37320 20334
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 37280 19372 37332 19378
rect 37280 19314 37332 19320
rect 37188 18760 37240 18766
rect 37188 18702 37240 18708
rect 37200 18290 37228 18702
rect 37292 18290 37320 19314
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 38292 18692 38344 18698
rect 38292 18634 38344 18640
rect 37188 18284 37240 18290
rect 37188 18226 37240 18232
rect 37280 18284 37332 18290
rect 37280 18226 37332 18232
rect 38304 17882 38332 18634
rect 38476 18624 38528 18630
rect 38476 18566 38528 18572
rect 38488 18086 38516 18566
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 38476 18080 38528 18086
rect 38476 18022 38528 18028
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 38292 17876 38344 17882
rect 38292 17818 38344 17824
rect 37188 17672 37240 17678
rect 37188 17614 37240 17620
rect 37832 17672 37884 17678
rect 37832 17614 37884 17620
rect 37096 17264 37148 17270
rect 37096 17206 37148 17212
rect 36820 17128 36872 17134
rect 36820 17070 36872 17076
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 35348 16244 35400 16250
rect 35348 16186 35400 16192
rect 33416 16108 33468 16114
rect 33416 16050 33468 16056
rect 34060 16108 34112 16114
rect 34060 16050 34112 16056
rect 34612 16108 34664 16114
rect 34612 16050 34664 16056
rect 32036 15904 32088 15910
rect 32036 15846 32088 15852
rect 32496 15904 32548 15910
rect 32496 15846 32548 15852
rect 33324 15904 33376 15910
rect 33324 15846 33376 15852
rect 32048 15502 32076 15846
rect 32508 15706 32536 15846
rect 32496 15700 32548 15706
rect 32496 15642 32548 15648
rect 32036 15496 32088 15502
rect 32036 15438 32088 15444
rect 33336 15434 33364 15846
rect 33324 15428 33376 15434
rect 33324 15370 33376 15376
rect 33232 15360 33284 15366
rect 33232 15302 33284 15308
rect 33244 15094 33272 15302
rect 33232 15088 33284 15094
rect 33232 15030 33284 15036
rect 33428 15026 33456 16050
rect 34072 15706 34100 16050
rect 34704 15972 34756 15978
rect 34704 15914 34756 15920
rect 34612 15904 34664 15910
rect 34612 15846 34664 15852
rect 34060 15700 34112 15706
rect 34060 15642 34112 15648
rect 34624 15502 34652 15846
rect 34716 15706 34744 15914
rect 34704 15700 34756 15706
rect 34704 15642 34756 15648
rect 34808 15502 34836 16186
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15706 35388 16186
rect 35348 15700 35400 15706
rect 35348 15642 35400 15648
rect 33784 15496 33836 15502
rect 33784 15438 33836 15444
rect 33876 15496 33928 15502
rect 33876 15438 33928 15444
rect 34336 15496 34388 15502
rect 34336 15438 34388 15444
rect 34612 15496 34664 15502
rect 34612 15438 34664 15444
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 33692 15360 33744 15366
rect 33692 15302 33744 15308
rect 33416 15020 33468 15026
rect 33416 14962 33468 14968
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 32588 14816 32640 14822
rect 32588 14758 32640 14764
rect 31944 14272 31996 14278
rect 31944 14214 31996 14220
rect 31956 12434 31984 14214
rect 32600 13938 32628 14758
rect 33612 14550 33640 14962
rect 33600 14544 33652 14550
rect 33600 14486 33652 14492
rect 33508 14340 33560 14346
rect 33508 14282 33560 14288
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 32680 13864 32732 13870
rect 32680 13806 32732 13812
rect 32496 13252 32548 13258
rect 32496 13194 32548 13200
rect 32508 12986 32536 13194
rect 32496 12980 32548 12986
rect 32496 12922 32548 12928
rect 31956 12406 32352 12434
rect 31864 12158 31984 12186
rect 31760 12096 31812 12102
rect 31760 12038 31812 12044
rect 31852 12096 31904 12102
rect 31852 12038 31904 12044
rect 31392 11688 31444 11694
rect 31392 11630 31444 11636
rect 31668 11688 31720 11694
rect 31668 11630 31720 11636
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31208 11144 31260 11150
rect 31208 11086 31260 11092
rect 31404 10266 31432 11630
rect 31680 11150 31708 11630
rect 31772 11558 31800 12038
rect 31760 11552 31812 11558
rect 31760 11494 31812 11500
rect 31772 11354 31800 11494
rect 31864 11354 31892 12038
rect 31760 11348 31812 11354
rect 31760 11290 31812 11296
rect 31852 11348 31904 11354
rect 31852 11290 31904 11296
rect 31956 11286 31984 12158
rect 31944 11280 31996 11286
rect 31944 11222 31996 11228
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31496 10742 31524 11086
rect 31576 11076 31628 11082
rect 31576 11018 31628 11024
rect 31588 10962 31616 11018
rect 31864 10962 31892 11086
rect 32324 11082 32352 12406
rect 32692 12374 32720 13806
rect 33140 13728 33192 13734
rect 33140 13670 33192 13676
rect 33152 13258 33180 13670
rect 33520 13394 33548 14282
rect 33508 13388 33560 13394
rect 33508 13330 33560 13336
rect 33140 13252 33192 13258
rect 33140 13194 33192 13200
rect 33704 12442 33732 15302
rect 33796 15162 33824 15438
rect 33784 15156 33836 15162
rect 33784 15098 33836 15104
rect 33888 15042 33916 15438
rect 34348 15094 34376 15438
rect 35348 15428 35400 15434
rect 35348 15370 35400 15376
rect 35360 15162 35388 15370
rect 36452 15360 36504 15366
rect 36452 15302 36504 15308
rect 36464 15162 36492 15302
rect 37108 15162 37136 17206
rect 37200 17134 37228 17614
rect 37844 17338 37872 17614
rect 37924 17604 37976 17610
rect 37924 17546 37976 17552
rect 37832 17332 37884 17338
rect 37832 17274 37884 17280
rect 37936 17134 37964 17546
rect 38304 17338 38332 17818
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 38292 17332 38344 17338
rect 38292 17274 38344 17280
rect 37188 17128 37240 17134
rect 37188 17070 37240 17076
rect 37924 17128 37976 17134
rect 37924 17070 37976 17076
rect 37936 16794 37964 17070
rect 38108 16992 38160 16998
rect 38108 16934 38160 16940
rect 37924 16788 37976 16794
rect 37924 16730 37976 16736
rect 38120 16590 38148 16934
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 38108 16584 38160 16590
rect 38108 16526 38160 16532
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 37372 15904 37424 15910
rect 37372 15846 37424 15852
rect 37384 15502 37412 15846
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 68296 15502 68324 27814
rect 37372 15496 37424 15502
rect 37372 15438 37424 15444
rect 68284 15496 68336 15502
rect 68284 15438 68336 15444
rect 37280 15360 37332 15366
rect 37280 15302 37332 15308
rect 35348 15156 35400 15162
rect 35348 15098 35400 15104
rect 36452 15156 36504 15162
rect 36452 15098 36504 15104
rect 37096 15156 37148 15162
rect 37096 15098 37148 15104
rect 33796 15014 33916 15042
rect 34336 15088 34388 15094
rect 34336 15030 34388 15036
rect 35716 15020 35768 15026
rect 33796 14414 33824 15014
rect 35716 14962 35768 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35728 14618 35756 14962
rect 37292 14822 37320 15302
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 67640 14952 67692 14958
rect 67640 14894 67692 14900
rect 37280 14816 37332 14822
rect 37280 14758 37332 14764
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 35716 14612 35768 14618
rect 35716 14554 35768 14560
rect 33784 14408 33836 14414
rect 33784 14350 33836 14356
rect 33796 14074 33824 14350
rect 35348 14340 35400 14346
rect 35348 14282 35400 14288
rect 34336 14272 34388 14278
rect 34336 14214 34388 14220
rect 33784 14068 33836 14074
rect 33784 14010 33836 14016
rect 34348 14006 34376 14214
rect 34336 14000 34388 14006
rect 34336 13942 34388 13948
rect 35360 13870 35388 14282
rect 36084 14272 36136 14278
rect 36084 14214 36136 14220
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 34796 13864 34848 13870
rect 34796 13806 34848 13812
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 34152 13728 34204 13734
rect 34152 13670 34204 13676
rect 34164 13258 34192 13670
rect 34808 13530 34836 13806
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34428 13524 34480 13530
rect 34428 13466 34480 13472
rect 34796 13524 34848 13530
rect 34796 13466 34848 13472
rect 34152 13252 34204 13258
rect 34152 13194 34204 13200
rect 34164 12918 34192 13194
rect 34440 12986 34468 13466
rect 34612 13252 34664 13258
rect 34612 13194 34664 13200
rect 34428 12980 34480 12986
rect 34428 12922 34480 12928
rect 34152 12912 34204 12918
rect 34440 12866 34468 12922
rect 34152 12854 34204 12860
rect 33968 12640 34020 12646
rect 33968 12582 34020 12588
rect 33692 12436 33744 12442
rect 33692 12378 33744 12384
rect 33980 12374 34008 12582
rect 34164 12442 34192 12854
rect 34244 12844 34296 12850
rect 34244 12786 34296 12792
rect 34348 12838 34468 12866
rect 34256 12442 34284 12786
rect 34152 12436 34204 12442
rect 34152 12378 34204 12384
rect 34244 12436 34296 12442
rect 34244 12378 34296 12384
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 33324 12368 33376 12374
rect 33324 12310 33376 12316
rect 33876 12368 33928 12374
rect 33876 12310 33928 12316
rect 33968 12368 34020 12374
rect 34348 12322 34376 12838
rect 34428 12708 34480 12714
rect 34428 12650 34480 12656
rect 33968 12310 34020 12316
rect 32864 12300 32916 12306
rect 32864 12242 32916 12248
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32496 11552 32548 11558
rect 32496 11494 32548 11500
rect 32508 11150 32536 11494
rect 32600 11218 32628 12038
rect 32876 11762 32904 12242
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32772 11756 32824 11762
rect 32772 11698 32824 11704
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 32784 11642 32812 11698
rect 32692 11614 32812 11642
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32312 11076 32364 11082
rect 32312 11018 32364 11024
rect 31588 10934 31892 10962
rect 31484 10736 31536 10742
rect 31484 10678 31536 10684
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31588 10130 31616 10934
rect 32692 10742 32720 11614
rect 32772 11552 32824 11558
rect 32772 11494 32824 11500
rect 32864 11552 32916 11558
rect 32864 11494 32916 11500
rect 32784 11286 32812 11494
rect 32772 11280 32824 11286
rect 32772 11222 32824 11228
rect 32680 10736 32732 10742
rect 32680 10678 32732 10684
rect 32876 10538 32904 11494
rect 32968 10810 32996 12174
rect 33140 11892 33192 11898
rect 33192 11852 33272 11880
rect 33140 11834 33192 11840
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 33152 11082 33180 11698
rect 33244 11626 33272 11852
rect 33232 11620 33284 11626
rect 33232 11562 33284 11568
rect 33140 11076 33192 11082
rect 33140 11018 33192 11024
rect 32956 10804 33008 10810
rect 32956 10746 33008 10752
rect 32864 10532 32916 10538
rect 32864 10474 32916 10480
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 31576 10124 31628 10130
rect 31576 10066 31628 10072
rect 31944 10124 31996 10130
rect 31944 10066 31996 10072
rect 32404 10124 32456 10130
rect 32404 10066 32456 10072
rect 29276 10056 29328 10062
rect 29276 9998 29328 10004
rect 30288 10056 30340 10062
rect 30288 9998 30340 10004
rect 31116 10056 31168 10062
rect 31116 9998 31168 10004
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29000 9512 29052 9518
rect 29000 9454 29052 9460
rect 28908 8900 28960 8906
rect 28828 8860 28908 8888
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 28540 8832 28592 8838
rect 28540 8774 28592 8780
rect 28276 8498 28304 8774
rect 28552 8498 28580 8774
rect 28828 8498 28856 8860
rect 28908 8842 28960 8848
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28540 8492 28592 8498
rect 28540 8434 28592 8440
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28908 8492 28960 8498
rect 29012 8480 29040 9454
rect 29564 9110 29592 9522
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29748 9178 29776 9318
rect 29736 9172 29788 9178
rect 29736 9114 29788 9120
rect 29552 9104 29604 9110
rect 29552 9046 29604 9052
rect 29644 9104 29696 9110
rect 29840 9058 29868 9318
rect 29696 9052 29868 9058
rect 29644 9046 29868 9052
rect 29276 8900 29328 8906
rect 29276 8842 29328 8848
rect 29288 8566 29316 8842
rect 29276 8560 29328 8566
rect 29276 8502 29328 8508
rect 28960 8452 29040 8480
rect 28908 8434 28960 8440
rect 28184 8090 28212 8434
rect 28276 8362 28304 8434
rect 28264 8356 28316 8362
rect 28264 8298 28316 8304
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 27540 7546 27568 7822
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27816 7478 27844 7686
rect 27804 7472 27856 7478
rect 27804 7414 27856 7420
rect 27908 7410 27936 7822
rect 28080 7472 28132 7478
rect 28080 7414 28132 7420
rect 27896 7404 27948 7410
rect 27896 7346 27948 7352
rect 27804 7336 27856 7342
rect 27804 7278 27856 7284
rect 27436 6860 27488 6866
rect 27436 6802 27488 6808
rect 27160 6792 27212 6798
rect 27160 6734 27212 6740
rect 26056 6724 26108 6730
rect 26056 6666 26108 6672
rect 26516 6724 26568 6730
rect 26516 6666 26568 6672
rect 26608 6724 26660 6730
rect 26608 6666 26660 6672
rect 27712 6724 27764 6730
rect 27712 6666 27764 6672
rect 26068 6458 26096 6666
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 26528 6322 26556 6666
rect 27724 6458 27752 6666
rect 27712 6452 27764 6458
rect 27712 6394 27764 6400
rect 27816 6390 27844 7278
rect 27988 7268 28040 7274
rect 27988 7210 28040 7216
rect 28000 6390 28028 7210
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 27988 6384 28040 6390
rect 27988 6326 28040 6332
rect 28092 6322 28120 7414
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28184 6390 28212 7142
rect 28828 6934 28856 8434
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29196 7886 29224 8230
rect 29564 8090 29592 9046
rect 29656 9042 29868 9046
rect 29656 9036 29880 9042
rect 29656 9030 29828 9036
rect 29828 8978 29880 8984
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 30208 8090 30236 8502
rect 30300 8294 30328 9998
rect 30932 9920 30984 9926
rect 30932 9862 30984 9868
rect 30748 9512 30800 9518
rect 30748 9454 30800 9460
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 30668 8634 30696 8910
rect 30760 8634 30788 9454
rect 30944 8634 30972 9862
rect 31128 9722 31156 9998
rect 31116 9716 31168 9722
rect 31116 9658 31168 9664
rect 31956 9654 31984 10066
rect 32416 9722 32444 10066
rect 32588 9920 32640 9926
rect 32588 9862 32640 9868
rect 32600 9722 32628 9862
rect 32404 9716 32456 9722
rect 32404 9658 32456 9664
rect 32588 9716 32640 9722
rect 32588 9658 32640 9664
rect 32692 9654 32720 10202
rect 33140 10192 33192 10198
rect 33244 10180 33272 11562
rect 33336 11150 33364 12310
rect 33888 12238 33916 12310
rect 34256 12294 34376 12322
rect 34256 12238 34284 12294
rect 33416 12232 33468 12238
rect 33416 12174 33468 12180
rect 33876 12232 33928 12238
rect 33876 12174 33928 12180
rect 34244 12232 34296 12238
rect 34440 12186 34468 12650
rect 34520 12640 34572 12646
rect 34520 12582 34572 12588
rect 34532 12306 34560 12582
rect 34520 12300 34572 12306
rect 34520 12242 34572 12248
rect 34244 12174 34296 12180
rect 33428 11830 33456 12174
rect 34348 12158 34468 12186
rect 33600 12096 33652 12102
rect 33600 12038 33652 12044
rect 33416 11824 33468 11830
rect 33416 11766 33468 11772
rect 33612 11558 33640 12038
rect 33692 11756 33744 11762
rect 33692 11698 33744 11704
rect 33600 11552 33652 11558
rect 33600 11494 33652 11500
rect 33704 11218 33732 11698
rect 34348 11354 34376 12158
rect 34624 11898 34652 13194
rect 35360 12782 35388 13806
rect 35452 13530 35480 13874
rect 35440 13524 35492 13530
rect 35440 13466 35492 13472
rect 34796 12776 34848 12782
rect 34796 12718 34848 12724
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 34808 12102 34836 12718
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35256 12164 35308 12170
rect 35256 12106 35308 12112
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 35268 11898 35296 12106
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 35256 11892 35308 11898
rect 35256 11834 35308 11840
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 34428 11688 34480 11694
rect 34428 11630 34480 11636
rect 34336 11348 34388 11354
rect 34336 11290 34388 11296
rect 34348 11218 34376 11290
rect 33692 11212 33744 11218
rect 33692 11154 33744 11160
rect 34336 11212 34388 11218
rect 34336 11154 34388 11160
rect 33324 11144 33376 11150
rect 33324 11086 33376 11092
rect 33192 10152 33272 10180
rect 33140 10134 33192 10140
rect 33152 10062 33180 10134
rect 32864 10056 32916 10062
rect 32864 9998 32916 10004
rect 33140 10056 33192 10062
rect 33140 9998 33192 10004
rect 32876 9722 32904 9998
rect 32864 9716 32916 9722
rect 32864 9658 32916 9664
rect 31208 9648 31260 9654
rect 31208 9590 31260 9596
rect 31944 9648 31996 9654
rect 32680 9648 32732 9654
rect 31944 9590 31996 9596
rect 32586 9616 32642 9625
rect 31220 9178 31248 9590
rect 32680 9590 32732 9596
rect 32586 9551 32588 9560
rect 32640 9551 32642 9560
rect 32588 9522 32640 9528
rect 32220 9376 32272 9382
rect 32220 9318 32272 9324
rect 31208 9172 31260 9178
rect 31208 9114 31260 9120
rect 32232 9042 32260 9318
rect 32220 9036 32272 9042
rect 32220 8978 32272 8984
rect 33244 8906 33272 10152
rect 33336 10130 33364 11086
rect 33600 11008 33652 11014
rect 33600 10950 33652 10956
rect 33416 10736 33468 10742
rect 33416 10678 33468 10684
rect 33428 10198 33456 10678
rect 33416 10192 33468 10198
rect 33468 10152 33548 10180
rect 33416 10134 33468 10140
rect 33324 10124 33376 10130
rect 33324 10066 33376 10072
rect 33336 9042 33364 10066
rect 33416 9920 33468 9926
rect 33416 9862 33468 9868
rect 33428 9722 33456 9862
rect 33416 9716 33468 9722
rect 33416 9658 33468 9664
rect 33416 9376 33468 9382
rect 33414 9344 33416 9353
rect 33468 9344 33470 9353
rect 33414 9279 33470 9288
rect 33520 9110 33548 10152
rect 33612 9654 33640 10950
rect 33704 10062 33732 11154
rect 34244 11144 34296 11150
rect 34244 11086 34296 11092
rect 34256 10266 34284 11086
rect 34440 10538 34468 11630
rect 34520 11144 34572 11150
rect 34520 11086 34572 11092
rect 34612 11144 34664 11150
rect 34612 11086 34664 11092
rect 34532 10810 34560 11086
rect 34520 10804 34572 10810
rect 34520 10746 34572 10752
rect 34428 10532 34480 10538
rect 34428 10474 34480 10480
rect 33784 10260 33836 10266
rect 33784 10202 33836 10208
rect 34244 10260 34296 10266
rect 34244 10202 34296 10208
rect 33692 10056 33744 10062
rect 33692 9998 33744 10004
rect 33600 9648 33652 9654
rect 33598 9616 33600 9625
rect 33652 9616 33654 9625
rect 33598 9551 33654 9560
rect 33508 9104 33560 9110
rect 33508 9046 33560 9052
rect 33324 9036 33376 9042
rect 33324 8978 33376 8984
rect 33704 8974 33732 9998
rect 33796 9450 33824 10202
rect 34244 9648 34296 9654
rect 34244 9590 34296 9596
rect 33968 9580 34020 9586
rect 33968 9522 34020 9528
rect 33980 9466 34008 9522
rect 33784 9444 33836 9450
rect 33784 9386 33836 9392
rect 33888 9438 34008 9466
rect 33888 9178 33916 9438
rect 34256 9353 34284 9590
rect 34242 9344 34298 9353
rect 34242 9279 34298 9288
rect 33876 9172 33928 9178
rect 33876 9114 33928 9120
rect 34624 9110 34652 11086
rect 34704 11008 34756 11014
rect 34704 10950 34756 10956
rect 34716 10742 34744 10950
rect 34704 10736 34756 10742
rect 34704 10678 34756 10684
rect 34808 10470 34836 11698
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35360 11234 35388 12718
rect 35452 12238 35480 13466
rect 35532 13320 35584 13326
rect 35532 13262 35584 13268
rect 35544 12374 35572 13262
rect 35808 13252 35860 13258
rect 35808 13194 35860 13200
rect 35992 13252 36044 13258
rect 35992 13194 36044 13200
rect 35820 12986 35848 13194
rect 35808 12980 35860 12986
rect 35808 12922 35860 12928
rect 35900 12912 35952 12918
rect 35900 12854 35952 12860
rect 35912 12442 35940 12854
rect 35900 12436 35952 12442
rect 35900 12378 35952 12384
rect 35532 12368 35584 12374
rect 35532 12310 35584 12316
rect 36004 12238 36032 13194
rect 36096 12238 36124 14214
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 36176 13932 36228 13938
rect 36176 13874 36228 13880
rect 36188 13462 36216 13874
rect 36360 13864 36412 13870
rect 36360 13806 36412 13812
rect 36268 13728 36320 13734
rect 36268 13670 36320 13676
rect 36176 13456 36228 13462
rect 36176 13398 36228 13404
rect 36280 13326 36308 13670
rect 36372 13394 36400 13806
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 36360 13388 36412 13394
rect 36360 13330 36412 13336
rect 36268 13320 36320 13326
rect 36268 13262 36320 13268
rect 36176 13252 36228 13258
rect 36176 13194 36228 13200
rect 35440 12232 35492 12238
rect 35440 12174 35492 12180
rect 35992 12232 36044 12238
rect 35992 12174 36044 12180
rect 36084 12232 36136 12238
rect 36084 12174 36136 12180
rect 35440 11892 35492 11898
rect 35440 11834 35492 11840
rect 35268 11218 35388 11234
rect 35256 11212 35388 11218
rect 35308 11206 35388 11212
rect 35256 11154 35308 11160
rect 35072 11144 35124 11150
rect 35124 11104 35204 11132
rect 35072 11086 35124 11092
rect 35176 10810 35204 11104
rect 35452 10810 35480 11834
rect 36188 11218 36216 13194
rect 36728 13184 36780 13190
rect 36728 13126 36780 13132
rect 36820 13184 36872 13190
rect 36820 13126 36872 13132
rect 36740 13002 36768 13126
rect 36648 12974 36768 13002
rect 36360 12912 36412 12918
rect 36360 12854 36412 12860
rect 36372 12442 36400 12854
rect 36360 12436 36412 12442
rect 36360 12378 36412 12384
rect 36648 12238 36676 12974
rect 36832 12646 36860 13126
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 36820 12640 36872 12646
rect 36820 12582 36872 12588
rect 37280 12640 37332 12646
rect 37280 12582 37332 12588
rect 37292 12306 37320 12582
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 37280 12300 37332 12306
rect 37280 12242 37332 12248
rect 36268 12232 36320 12238
rect 36268 12174 36320 12180
rect 36636 12232 36688 12238
rect 36636 12174 36688 12180
rect 36176 11212 36228 11218
rect 36176 11154 36228 11160
rect 35900 11008 35952 11014
rect 35900 10950 35952 10956
rect 35912 10810 35940 10950
rect 35164 10804 35216 10810
rect 35164 10746 35216 10752
rect 35440 10804 35492 10810
rect 35440 10746 35492 10752
rect 35900 10804 35952 10810
rect 35900 10746 35952 10752
rect 36280 10674 36308 12174
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 36820 11076 36872 11082
rect 36820 11018 36872 11024
rect 36544 11008 36596 11014
rect 36544 10950 36596 10956
rect 36268 10668 36320 10674
rect 36268 10610 36320 10616
rect 36556 10606 36584 10950
rect 36832 10810 36860 11018
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 36820 10804 36872 10810
rect 36820 10746 36872 10752
rect 35992 10600 36044 10606
rect 35992 10542 36044 10548
rect 36544 10600 36596 10606
rect 36544 10542 36596 10548
rect 34796 10464 34848 10470
rect 34796 10406 34848 10412
rect 34808 10062 34836 10406
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35256 10124 35308 10130
rect 35256 10066 35308 10072
rect 34796 10056 34848 10062
rect 34796 9998 34848 10004
rect 34704 9920 34756 9926
rect 34704 9862 34756 9868
rect 34716 9518 34744 9862
rect 34704 9512 34756 9518
rect 34704 9454 34756 9460
rect 34808 9178 34836 9998
rect 35268 9722 35296 10066
rect 35532 9920 35584 9926
rect 35532 9862 35584 9868
rect 35256 9716 35308 9722
rect 35256 9658 35308 9664
rect 35544 9382 35572 9862
rect 36004 9586 36032 10542
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 34796 9172 34848 9178
rect 34796 9114 34848 9120
rect 34612 9104 34664 9110
rect 34612 9046 34664 9052
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 32036 8900 32088 8906
rect 32036 8842 32088 8848
rect 33232 8900 33284 8906
rect 33232 8842 33284 8848
rect 31208 8832 31260 8838
rect 31208 8774 31260 8780
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30748 8628 30800 8634
rect 30748 8570 30800 8576
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 31220 8430 31248 8774
rect 32048 8634 32076 8842
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 32036 8628 32088 8634
rect 32036 8570 32088 8576
rect 31208 8424 31260 8430
rect 31208 8366 31260 8372
rect 30288 8288 30340 8294
rect 30288 8230 30340 8236
rect 29552 8084 29604 8090
rect 29552 8026 29604 8032
rect 30196 8084 30248 8090
rect 30196 8026 30248 8032
rect 30300 7886 30328 8230
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 29184 7880 29236 7886
rect 29184 7822 29236 7828
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 29736 7812 29788 7818
rect 29736 7754 29788 7760
rect 28816 6928 28868 6934
rect 28816 6870 28868 6876
rect 28264 6860 28316 6866
rect 28264 6802 28316 6808
rect 28172 6384 28224 6390
rect 28172 6326 28224 6332
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 28080 6316 28132 6322
rect 28080 6258 28132 6264
rect 28276 6186 28304 6802
rect 29748 6798 29776 7754
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 29460 6656 29512 6662
rect 29460 6598 29512 6604
rect 29472 6254 29500 6598
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 29460 6248 29512 6254
rect 29460 6190 29512 6196
rect 28264 6180 28316 6186
rect 28264 6122 28316 6128
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 43260 2848 43312 2854
rect 43260 2790 43312 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 43272 2446 43300 2790
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 67652 2446 67680 14894
rect 68468 10056 68520 10062
rect 68468 9998 68520 10004
rect 68480 9625 68508 9998
rect 68466 9616 68522 9625
rect 68466 9551 68522 9560
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 43260 2440 43312 2446
rect 43260 2382 43312 2388
rect 67640 2440 67692 2446
rect 67640 2382 67692 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 26528 1306 26556 2382
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 68008 2304 68060 2310
rect 68008 2246 68060 2252
rect 26436 1278 26556 1306
rect 26436 800 26464 1278
rect 43824 800 43852 2246
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 18 0 74 800
rect 8390 0 8446 800
rect 17406 0 17462 800
rect 26422 0 26478 800
rect 34794 0 34850 800
rect 43810 0 43866 800
rect 52826 0 52882 800
rect 61198 0 61254 800
rect 68020 105 68048 2246
rect 68006 96 68062 105
rect 68006 31 68062 40
<< via2 >>
rect 19580 67482 19636 67484
rect 19660 67482 19716 67484
rect 19740 67482 19796 67484
rect 19820 67482 19876 67484
rect 19580 67430 19626 67482
rect 19626 67430 19636 67482
rect 19660 67430 19690 67482
rect 19690 67430 19702 67482
rect 19702 67430 19716 67482
rect 19740 67430 19754 67482
rect 19754 67430 19766 67482
rect 19766 67430 19796 67482
rect 19820 67430 19830 67482
rect 19830 67430 19876 67482
rect 19580 67428 19636 67430
rect 19660 67428 19716 67430
rect 19740 67428 19796 67430
rect 19820 67428 19876 67430
rect 50300 67482 50356 67484
rect 50380 67482 50436 67484
rect 50460 67482 50516 67484
rect 50540 67482 50596 67484
rect 50300 67430 50346 67482
rect 50346 67430 50356 67482
rect 50380 67430 50410 67482
rect 50410 67430 50422 67482
rect 50422 67430 50436 67482
rect 50460 67430 50474 67482
rect 50474 67430 50486 67482
rect 50486 67430 50516 67482
rect 50540 67430 50550 67482
rect 50550 67430 50596 67482
rect 50300 67428 50356 67430
rect 50380 67428 50436 67430
rect 50460 67428 50516 67430
rect 50540 67428 50596 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 19580 66394 19636 66396
rect 19660 66394 19716 66396
rect 19740 66394 19796 66396
rect 19820 66394 19876 66396
rect 19580 66342 19626 66394
rect 19626 66342 19636 66394
rect 19660 66342 19690 66394
rect 19690 66342 19702 66394
rect 19702 66342 19716 66394
rect 19740 66342 19754 66394
rect 19754 66342 19766 66394
rect 19766 66342 19796 66394
rect 19820 66342 19830 66394
rect 19830 66342 19876 66394
rect 19580 66340 19636 66342
rect 19660 66340 19716 66342
rect 19740 66340 19796 66342
rect 19820 66340 19876 66342
rect 50300 66394 50356 66396
rect 50380 66394 50436 66396
rect 50460 66394 50516 66396
rect 50540 66394 50596 66396
rect 50300 66342 50346 66394
rect 50346 66342 50356 66394
rect 50380 66342 50410 66394
rect 50410 66342 50422 66394
rect 50422 66342 50436 66394
rect 50460 66342 50474 66394
rect 50474 66342 50486 66394
rect 50486 66342 50516 66394
rect 50540 66342 50550 66394
rect 50550 66342 50596 66394
rect 50300 66340 50356 66342
rect 50380 66340 50436 66342
rect 50460 66340 50516 66342
rect 50540 66340 50596 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 19580 65306 19636 65308
rect 19660 65306 19716 65308
rect 19740 65306 19796 65308
rect 19820 65306 19876 65308
rect 19580 65254 19626 65306
rect 19626 65254 19636 65306
rect 19660 65254 19690 65306
rect 19690 65254 19702 65306
rect 19702 65254 19716 65306
rect 19740 65254 19754 65306
rect 19754 65254 19766 65306
rect 19766 65254 19796 65306
rect 19820 65254 19830 65306
rect 19830 65254 19876 65306
rect 19580 65252 19636 65254
rect 19660 65252 19716 65254
rect 19740 65252 19796 65254
rect 19820 65252 19876 65254
rect 50300 65306 50356 65308
rect 50380 65306 50436 65308
rect 50460 65306 50516 65308
rect 50540 65306 50596 65308
rect 50300 65254 50346 65306
rect 50346 65254 50356 65306
rect 50380 65254 50410 65306
rect 50410 65254 50422 65306
rect 50422 65254 50436 65306
rect 50460 65254 50474 65306
rect 50474 65254 50486 65306
rect 50486 65254 50516 65306
rect 50540 65254 50550 65306
rect 50550 65254 50596 65306
rect 50300 65252 50356 65254
rect 50380 65252 50436 65254
rect 50460 65252 50516 65254
rect 50540 65252 50596 65254
rect 1398 64776 1454 64832
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 34940 64762 34996 64764
rect 35020 64762 35076 64764
rect 35100 64762 35156 64764
rect 35180 64762 35236 64764
rect 34940 64710 34986 64762
rect 34986 64710 34996 64762
rect 35020 64710 35050 64762
rect 35050 64710 35062 64762
rect 35062 64710 35076 64762
rect 35100 64710 35114 64762
rect 35114 64710 35126 64762
rect 35126 64710 35156 64762
rect 35180 64710 35190 64762
rect 35190 64710 35236 64762
rect 34940 64708 34996 64710
rect 35020 64708 35076 64710
rect 35100 64708 35156 64710
rect 35180 64708 35236 64710
rect 65660 64762 65716 64764
rect 65740 64762 65796 64764
rect 65820 64762 65876 64764
rect 65900 64762 65956 64764
rect 65660 64710 65706 64762
rect 65706 64710 65716 64762
rect 65740 64710 65770 64762
rect 65770 64710 65782 64762
rect 65782 64710 65796 64762
rect 65820 64710 65834 64762
rect 65834 64710 65846 64762
rect 65846 64710 65876 64762
rect 65900 64710 65910 64762
rect 65910 64710 65956 64762
rect 65660 64708 65716 64710
rect 65740 64708 65796 64710
rect 65820 64708 65876 64710
rect 65900 64708 65956 64710
rect 19580 64218 19636 64220
rect 19660 64218 19716 64220
rect 19740 64218 19796 64220
rect 19820 64218 19876 64220
rect 19580 64166 19626 64218
rect 19626 64166 19636 64218
rect 19660 64166 19690 64218
rect 19690 64166 19702 64218
rect 19702 64166 19716 64218
rect 19740 64166 19754 64218
rect 19754 64166 19766 64218
rect 19766 64166 19796 64218
rect 19820 64166 19830 64218
rect 19830 64166 19876 64218
rect 19580 64164 19636 64166
rect 19660 64164 19716 64166
rect 19740 64164 19796 64166
rect 19820 64164 19876 64166
rect 50300 64218 50356 64220
rect 50380 64218 50436 64220
rect 50460 64218 50516 64220
rect 50540 64218 50596 64220
rect 50300 64166 50346 64218
rect 50346 64166 50356 64218
rect 50380 64166 50410 64218
rect 50410 64166 50422 64218
rect 50422 64166 50436 64218
rect 50460 64166 50474 64218
rect 50474 64166 50486 64218
rect 50486 64166 50516 64218
rect 50540 64166 50550 64218
rect 50550 64166 50596 64218
rect 50300 64164 50356 64166
rect 50380 64164 50436 64166
rect 50460 64164 50516 64166
rect 50540 64164 50596 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 34940 63674 34996 63676
rect 35020 63674 35076 63676
rect 35100 63674 35156 63676
rect 35180 63674 35236 63676
rect 34940 63622 34986 63674
rect 34986 63622 34996 63674
rect 35020 63622 35050 63674
rect 35050 63622 35062 63674
rect 35062 63622 35076 63674
rect 35100 63622 35114 63674
rect 35114 63622 35126 63674
rect 35126 63622 35156 63674
rect 35180 63622 35190 63674
rect 35190 63622 35236 63674
rect 34940 63620 34996 63622
rect 35020 63620 35076 63622
rect 35100 63620 35156 63622
rect 35180 63620 35236 63622
rect 65660 63674 65716 63676
rect 65740 63674 65796 63676
rect 65820 63674 65876 63676
rect 65900 63674 65956 63676
rect 65660 63622 65706 63674
rect 65706 63622 65716 63674
rect 65740 63622 65770 63674
rect 65770 63622 65782 63674
rect 65782 63622 65796 63674
rect 65820 63622 65834 63674
rect 65834 63622 65846 63674
rect 65846 63622 65876 63674
rect 65900 63622 65910 63674
rect 65910 63622 65956 63674
rect 65660 63620 65716 63622
rect 65740 63620 65796 63622
rect 65820 63620 65876 63622
rect 65900 63620 65956 63622
rect 19580 63130 19636 63132
rect 19660 63130 19716 63132
rect 19740 63130 19796 63132
rect 19820 63130 19876 63132
rect 19580 63078 19626 63130
rect 19626 63078 19636 63130
rect 19660 63078 19690 63130
rect 19690 63078 19702 63130
rect 19702 63078 19716 63130
rect 19740 63078 19754 63130
rect 19754 63078 19766 63130
rect 19766 63078 19796 63130
rect 19820 63078 19830 63130
rect 19830 63078 19876 63130
rect 19580 63076 19636 63078
rect 19660 63076 19716 63078
rect 19740 63076 19796 63078
rect 19820 63076 19876 63078
rect 50300 63130 50356 63132
rect 50380 63130 50436 63132
rect 50460 63130 50516 63132
rect 50540 63130 50596 63132
rect 50300 63078 50346 63130
rect 50346 63078 50356 63130
rect 50380 63078 50410 63130
rect 50410 63078 50422 63130
rect 50422 63078 50436 63130
rect 50460 63078 50474 63130
rect 50474 63078 50486 63130
rect 50486 63078 50516 63130
rect 50540 63078 50550 63130
rect 50550 63078 50596 63130
rect 50300 63076 50356 63078
rect 50380 63076 50436 63078
rect 50460 63076 50516 63078
rect 50540 63076 50596 63078
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 34940 62586 34996 62588
rect 35020 62586 35076 62588
rect 35100 62586 35156 62588
rect 35180 62586 35236 62588
rect 34940 62534 34986 62586
rect 34986 62534 34996 62586
rect 35020 62534 35050 62586
rect 35050 62534 35062 62586
rect 35062 62534 35076 62586
rect 35100 62534 35114 62586
rect 35114 62534 35126 62586
rect 35126 62534 35156 62586
rect 35180 62534 35190 62586
rect 35190 62534 35236 62586
rect 34940 62532 34996 62534
rect 35020 62532 35076 62534
rect 35100 62532 35156 62534
rect 35180 62532 35236 62534
rect 65660 62586 65716 62588
rect 65740 62586 65796 62588
rect 65820 62586 65876 62588
rect 65900 62586 65956 62588
rect 65660 62534 65706 62586
rect 65706 62534 65716 62586
rect 65740 62534 65770 62586
rect 65770 62534 65782 62586
rect 65782 62534 65796 62586
rect 65820 62534 65834 62586
rect 65834 62534 65846 62586
rect 65846 62534 65876 62586
rect 65900 62534 65910 62586
rect 65910 62534 65956 62586
rect 65660 62532 65716 62534
rect 65740 62532 65796 62534
rect 65820 62532 65876 62534
rect 65900 62532 65956 62534
rect 19580 62042 19636 62044
rect 19660 62042 19716 62044
rect 19740 62042 19796 62044
rect 19820 62042 19876 62044
rect 19580 61990 19626 62042
rect 19626 61990 19636 62042
rect 19660 61990 19690 62042
rect 19690 61990 19702 62042
rect 19702 61990 19716 62042
rect 19740 61990 19754 62042
rect 19754 61990 19766 62042
rect 19766 61990 19796 62042
rect 19820 61990 19830 62042
rect 19830 61990 19876 62042
rect 19580 61988 19636 61990
rect 19660 61988 19716 61990
rect 19740 61988 19796 61990
rect 19820 61988 19876 61990
rect 50300 62042 50356 62044
rect 50380 62042 50436 62044
rect 50460 62042 50516 62044
rect 50540 62042 50596 62044
rect 50300 61990 50346 62042
rect 50346 61990 50356 62042
rect 50380 61990 50410 62042
rect 50410 61990 50422 62042
rect 50422 61990 50436 62042
rect 50460 61990 50474 62042
rect 50474 61990 50486 62042
rect 50486 61990 50516 62042
rect 50540 61990 50550 62042
rect 50550 61990 50596 62042
rect 50300 61988 50356 61990
rect 50380 61988 50436 61990
rect 50460 61988 50516 61990
rect 50540 61988 50596 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 65660 61498 65716 61500
rect 65740 61498 65796 61500
rect 65820 61498 65876 61500
rect 65900 61498 65956 61500
rect 65660 61446 65706 61498
rect 65706 61446 65716 61498
rect 65740 61446 65770 61498
rect 65770 61446 65782 61498
rect 65782 61446 65796 61498
rect 65820 61446 65834 61498
rect 65834 61446 65846 61498
rect 65846 61446 65876 61498
rect 65900 61446 65910 61498
rect 65910 61446 65956 61498
rect 65660 61444 65716 61446
rect 65740 61444 65796 61446
rect 65820 61444 65876 61446
rect 65900 61444 65956 61446
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 65660 60410 65716 60412
rect 65740 60410 65796 60412
rect 65820 60410 65876 60412
rect 65900 60410 65956 60412
rect 65660 60358 65706 60410
rect 65706 60358 65716 60410
rect 65740 60358 65770 60410
rect 65770 60358 65782 60410
rect 65782 60358 65796 60410
rect 65820 60358 65834 60410
rect 65834 60358 65846 60410
rect 65846 60358 65876 60410
rect 65900 60358 65910 60410
rect 65910 60358 65956 60410
rect 65660 60356 65716 60358
rect 65740 60356 65796 60358
rect 65820 60356 65876 60358
rect 65900 60356 65956 60358
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 65660 59322 65716 59324
rect 65740 59322 65796 59324
rect 65820 59322 65876 59324
rect 65900 59322 65956 59324
rect 65660 59270 65706 59322
rect 65706 59270 65716 59322
rect 65740 59270 65770 59322
rect 65770 59270 65782 59322
rect 65782 59270 65796 59322
rect 65820 59270 65834 59322
rect 65834 59270 65846 59322
rect 65846 59270 65876 59322
rect 65900 59270 65910 59322
rect 65910 59270 65956 59322
rect 65660 59268 65716 59270
rect 65740 59268 65796 59270
rect 65820 59268 65876 59270
rect 65900 59268 65956 59270
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 65660 58234 65716 58236
rect 65740 58234 65796 58236
rect 65820 58234 65876 58236
rect 65900 58234 65956 58236
rect 65660 58182 65706 58234
rect 65706 58182 65716 58234
rect 65740 58182 65770 58234
rect 65770 58182 65782 58234
rect 65782 58182 65796 58234
rect 65820 58182 65834 58234
rect 65834 58182 65846 58234
rect 65846 58182 65876 58234
rect 65900 58182 65910 58234
rect 65910 58182 65956 58234
rect 65660 58180 65716 58182
rect 65740 58180 65796 58182
rect 65820 58180 65876 58182
rect 65900 58180 65956 58182
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 68466 55800 68522 55856
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 938 46316 940 46336
rect 940 46316 992 46336
rect 992 46316 994 46336
rect 938 46280 994 46316
rect 938 36760 994 36816
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4066 18400 4122 18456
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 13910 20460 13966 20496
rect 13910 20440 13912 20460
rect 13912 20440 13964 20460
rect 13964 20440 13966 20460
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 16302 19372 16358 19408
rect 16302 19352 16304 19372
rect 16304 19352 16356 19372
rect 16356 19352 16358 19372
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 18878 17212 18880 17232
rect 18880 17212 18932 17232
rect 18932 17212 18934 17232
rect 18878 17176 18934 17212
rect 18970 17040 19026 17096
rect 20166 19352 20222 19408
rect 20810 19352 20866 19408
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19246 16632 19302 16688
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 18878 14864 18934 14920
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 17038 9580 17094 9616
rect 17038 9560 17040 9580
rect 17040 9560 17092 9580
rect 17092 9560 17094 9580
rect 19338 11736 19394 11792
rect 18510 9560 18566 9616
rect 18510 9444 18566 9480
rect 18510 9424 18512 9444
rect 18512 9424 18564 9444
rect 18564 9424 18566 9444
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19154 9424 19210 9480
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 18694 8628 18750 8664
rect 18694 8608 18696 8628
rect 18696 8608 18748 8628
rect 18748 8608 18750 8628
rect 19154 8608 19210 8664
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 22558 20440 22614 20496
rect 21822 11772 21824 11792
rect 21824 11772 21876 11792
rect 21876 11772 21878 11792
rect 21822 11736 21878 11772
rect 23110 17212 23112 17232
rect 23112 17212 23164 17232
rect 23164 17212 23166 17232
rect 23110 17176 23166 17212
rect 23478 17040 23534 17096
rect 23662 14068 23718 14104
rect 23662 14048 23664 14068
rect 23664 14048 23716 14068
rect 23716 14048 23718 14068
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 68834 27920 68890 27976
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 30470 26444 30526 26480
rect 30470 26424 30472 26444
rect 30472 26424 30524 26444
rect 30524 26424 30526 26444
rect 24122 15020 24178 15056
rect 24122 15000 24124 15020
rect 24124 15000 24176 15020
rect 24176 15000 24178 15020
rect 24766 14864 24822 14920
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 33046 26444 33102 26480
rect 33046 26424 33048 26444
rect 33048 26424 33100 26444
rect 33100 26424 33102 26444
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 27158 16632 27214 16688
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 27434 15000 27490 15056
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 26882 14048 26938 14104
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 32586 9580 32642 9616
rect 32586 9560 32588 9580
rect 32588 9560 32640 9580
rect 32640 9560 32642 9580
rect 33414 9324 33416 9344
rect 33416 9324 33468 9344
rect 33468 9324 33470 9344
rect 33414 9288 33470 9324
rect 33598 9596 33600 9616
rect 33600 9596 33652 9616
rect 33652 9596 33654 9616
rect 33598 9560 33654 9596
rect 34242 9288 34298 9344
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 68466 9560 68522 9616
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 68006 40 68062 96
<< metal3 >>
rect 19570 67488 19886 67489
rect 19570 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19886 67488
rect 19570 67423 19886 67424
rect 50290 67488 50606 67489
rect 50290 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50606 67488
rect 50290 67423 50606 67424
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 19570 66400 19886 66401
rect 19570 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19886 66400
rect 19570 66335 19886 66336
rect 50290 66400 50606 66401
rect 50290 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50606 66400
rect 50290 66335 50606 66336
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 19570 65312 19886 65313
rect 19570 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19886 65312
rect 19570 65247 19886 65248
rect 50290 65312 50606 65313
rect 50290 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50606 65312
rect 69200 65288 70000 65408
rect 50290 65247 50606 65248
rect 1393 64834 1459 64837
rect 798 64832 1459 64834
rect 798 64776 1398 64832
rect 1454 64776 1459 64832
rect 798 64774 1459 64776
rect 798 64728 858 64774
rect 1393 64771 1459 64774
rect 0 64638 858 64728
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 34930 64768 35246 64769
rect 34930 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35246 64768
rect 34930 64703 35246 64704
rect 65650 64768 65966 64769
rect 65650 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65966 64768
rect 65650 64703 65966 64704
rect 0 64608 800 64638
rect 19570 64224 19886 64225
rect 19570 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19886 64224
rect 19570 64159 19886 64160
rect 50290 64224 50606 64225
rect 50290 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50606 64224
rect 50290 64159 50606 64160
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 34930 63680 35246 63681
rect 34930 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35246 63680
rect 34930 63615 35246 63616
rect 65650 63680 65966 63681
rect 65650 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65966 63680
rect 65650 63615 65966 63616
rect 19570 63136 19886 63137
rect 19570 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19886 63136
rect 19570 63071 19886 63072
rect 50290 63136 50606 63137
rect 50290 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50606 63136
rect 50290 63071 50606 63072
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 34930 62592 35246 62593
rect 34930 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35246 62592
rect 34930 62527 35246 62528
rect 65650 62592 65966 62593
rect 65650 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65966 62592
rect 65650 62527 65966 62528
rect 19570 62048 19886 62049
rect 19570 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19886 62048
rect 19570 61983 19886 61984
rect 50290 62048 50606 62049
rect 50290 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50606 62048
rect 50290 61983 50606 61984
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 34930 61439 35246 61440
rect 65650 61504 65966 61505
rect 65650 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65966 61504
rect 65650 61439 65966 61440
rect 19570 60960 19886 60961
rect 19570 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19886 60960
rect 19570 60895 19886 60896
rect 50290 60960 50606 60961
rect 50290 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50606 60960
rect 50290 60895 50606 60896
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 34930 60351 35246 60352
rect 65650 60416 65966 60417
rect 65650 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65966 60416
rect 65650 60351 65966 60352
rect 19570 59872 19886 59873
rect 19570 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19886 59872
rect 19570 59807 19886 59808
rect 50290 59872 50606 59873
rect 50290 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50606 59872
rect 50290 59807 50606 59808
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 34930 59328 35246 59329
rect 34930 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35246 59328
rect 34930 59263 35246 59264
rect 65650 59328 65966 59329
rect 65650 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65966 59328
rect 65650 59263 65966 59264
rect 19570 58784 19886 58785
rect 19570 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19886 58784
rect 19570 58719 19886 58720
rect 50290 58784 50606 58785
rect 50290 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50606 58784
rect 50290 58719 50606 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 34930 58240 35246 58241
rect 34930 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35246 58240
rect 34930 58175 35246 58176
rect 65650 58240 65966 58241
rect 65650 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65966 58240
rect 65650 58175 65966 58176
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 65650 55999 65966 56000
rect 0 55768 800 55888
rect 68461 55858 68527 55861
rect 69200 55858 70000 55888
rect 68461 55856 70000 55858
rect 68461 55800 68466 55856
rect 68522 55800 70000 55856
rect 68461 55798 70000 55800
rect 68461 55795 68527 55798
rect 69200 55768 70000 55798
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 65650 53823 65966 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 65650 48383 65966 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 0 46338 800 46368
rect 933 46338 999 46341
rect 0 46336 999 46338
rect 0 46280 938 46336
rect 994 46280 999 46336
rect 0 46278 999 46280
rect 0 46248 800 46278
rect 933 46275 999 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 69200 46248 70000 46368
rect 65650 46207 65966 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 65650 44031 65966 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 65650 42943 65966 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 69200 37408 70000 37528
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 0 27888 800 28008
rect 68829 27978 68895 27981
rect 69200 27978 70000 28008
rect 68829 27976 70000 27978
rect 68829 27920 68834 27976
rect 68890 27920 70000 27976
rect 68829 27918 70000 27920
rect 68829 27915 68895 27918
rect 69200 27888 70000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 30465 26482 30531 26485
rect 33041 26482 33107 26485
rect 30465 26480 33107 26482
rect 30465 26424 30470 26480
rect 30526 26424 33046 26480
rect 33102 26424 33107 26480
rect 30465 26422 33107 26424
rect 30465 26419 30531 26422
rect 33041 26419 33107 26422
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 13905 20498 13971 20501
rect 22553 20498 22619 20501
rect 13905 20496 22619 20498
rect 13905 20440 13910 20496
rect 13966 20440 22558 20496
rect 22614 20440 22619 20496
rect 13905 20438 22619 20440
rect 13905 20435 13971 20438
rect 22553 20435 22619 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 16297 19410 16363 19413
rect 20161 19410 20227 19413
rect 20805 19410 20871 19413
rect 16297 19408 20871 19410
rect 16297 19352 16302 19408
rect 16358 19352 20166 19408
rect 20222 19352 20810 19408
rect 20866 19352 20871 19408
rect 16297 19350 20871 19352
rect 16297 19347 16363 19350
rect 20161 19347 20227 19350
rect 20805 19347 20871 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 19570 18528 19886 18529
rect 0 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 4061 18458 4127 18461
rect 0 18456 4127 18458
rect 0 18400 4066 18456
rect 4122 18400 4127 18456
rect 0 18398 4127 18400
rect 0 18368 800 18398
rect 4061 18395 4127 18398
rect 69200 18368 70000 18488
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 18873 17234 18939 17237
rect 23105 17234 23171 17237
rect 18873 17232 23171 17234
rect 18873 17176 18878 17232
rect 18934 17176 23110 17232
rect 23166 17176 23171 17232
rect 18873 17174 23171 17176
rect 18873 17171 18939 17174
rect 23105 17171 23171 17174
rect 18965 17098 19031 17101
rect 23473 17098 23539 17101
rect 18965 17096 23539 17098
rect 18965 17040 18970 17096
rect 19026 17040 23478 17096
rect 23534 17040 23539 17096
rect 18965 17038 23539 17040
rect 18965 17035 19031 17038
rect 23473 17035 23539 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 19241 16690 19307 16693
rect 27153 16690 27219 16693
rect 19241 16688 27219 16690
rect 19241 16632 19246 16688
rect 19302 16632 27158 16688
rect 27214 16632 27219 16688
rect 19241 16630 27219 16632
rect 19241 16627 19307 16630
rect 27153 16627 27219 16630
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 24117 15058 24183 15061
rect 27429 15058 27495 15061
rect 24117 15056 27495 15058
rect 24117 15000 24122 15056
rect 24178 15000 27434 15056
rect 27490 15000 27495 15056
rect 24117 14998 27495 15000
rect 24117 14995 24183 14998
rect 27429 14995 27495 14998
rect 18873 14922 18939 14925
rect 24761 14922 24827 14925
rect 18873 14920 24827 14922
rect 18873 14864 18878 14920
rect 18934 14864 24766 14920
rect 24822 14864 24827 14920
rect 18873 14862 24827 14864
rect 18873 14859 18939 14862
rect 24761 14859 24827 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 23657 14106 23723 14109
rect 26877 14106 26943 14109
rect 23657 14104 26943 14106
rect 23657 14048 23662 14104
rect 23718 14048 26882 14104
rect 26938 14048 26943 14104
rect 23657 14046 26943 14048
rect 23657 14043 23723 14046
rect 26877 14043 26943 14046
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 19333 11794 19399 11797
rect 21817 11794 21883 11797
rect 19333 11792 21883 11794
rect 19333 11736 19338 11792
rect 19394 11736 21822 11792
rect 21878 11736 21883 11792
rect 19333 11734 21883 11736
rect 19333 11731 19399 11734
rect 21817 11731 21883 11734
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 17033 9618 17099 9621
rect 18505 9618 18571 9621
rect 17033 9616 18571 9618
rect 17033 9560 17038 9616
rect 17094 9560 18510 9616
rect 18566 9560 18571 9616
rect 17033 9558 18571 9560
rect 17033 9555 17099 9558
rect 18505 9555 18571 9558
rect 32581 9618 32647 9621
rect 33593 9618 33659 9621
rect 32581 9616 33659 9618
rect 32581 9560 32586 9616
rect 32642 9560 33598 9616
rect 33654 9560 33659 9616
rect 32581 9558 33659 9560
rect 32581 9555 32647 9558
rect 33593 9555 33659 9558
rect 68461 9618 68527 9621
rect 69200 9618 70000 9648
rect 68461 9616 70000 9618
rect 68461 9560 68466 9616
rect 68522 9560 70000 9616
rect 68461 9558 70000 9560
rect 68461 9555 68527 9558
rect 69200 9528 70000 9558
rect 18505 9482 18571 9485
rect 19149 9482 19215 9485
rect 18505 9480 19215 9482
rect 18505 9424 18510 9480
rect 18566 9424 19154 9480
rect 19210 9424 19215 9480
rect 18505 9422 19215 9424
rect 18505 9419 18571 9422
rect 19149 9419 19215 9422
rect 33409 9346 33475 9349
rect 34237 9346 34303 9349
rect 33409 9344 34303 9346
rect 33409 9288 33414 9344
rect 33470 9288 34242 9344
rect 34298 9288 34303 9344
rect 33409 9286 34303 9288
rect 33409 9283 33475 9286
rect 34237 9283 34303 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 0 8848 800 8968
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 18689 8666 18755 8669
rect 19149 8666 19215 8669
rect 18689 8664 19215 8666
rect 18689 8608 18694 8664
rect 18750 8608 19154 8664
rect 19210 8608 19215 8664
rect 18689 8606 19215 8608
rect 18689 8603 18755 8606
rect 19149 8603 19215 8606
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 68001 98 68067 101
rect 69200 98 70000 128
rect 68001 96 70000 98
rect 68001 40 68006 96
rect 68062 40 70000 96
rect 68001 38 70000 40
rect 68001 35 68067 38
rect 69200 8 70000 38
<< via3 >>
rect 19576 67484 19640 67488
rect 19576 67428 19580 67484
rect 19580 67428 19636 67484
rect 19636 67428 19640 67484
rect 19576 67424 19640 67428
rect 19656 67484 19720 67488
rect 19656 67428 19660 67484
rect 19660 67428 19716 67484
rect 19716 67428 19720 67484
rect 19656 67424 19720 67428
rect 19736 67484 19800 67488
rect 19736 67428 19740 67484
rect 19740 67428 19796 67484
rect 19796 67428 19800 67484
rect 19736 67424 19800 67428
rect 19816 67484 19880 67488
rect 19816 67428 19820 67484
rect 19820 67428 19876 67484
rect 19876 67428 19880 67484
rect 19816 67424 19880 67428
rect 50296 67484 50360 67488
rect 50296 67428 50300 67484
rect 50300 67428 50356 67484
rect 50356 67428 50360 67484
rect 50296 67424 50360 67428
rect 50376 67484 50440 67488
rect 50376 67428 50380 67484
rect 50380 67428 50436 67484
rect 50436 67428 50440 67484
rect 50376 67424 50440 67428
rect 50456 67484 50520 67488
rect 50456 67428 50460 67484
rect 50460 67428 50516 67484
rect 50516 67428 50520 67484
rect 50456 67424 50520 67428
rect 50536 67484 50600 67488
rect 50536 67428 50540 67484
rect 50540 67428 50596 67484
rect 50596 67428 50600 67484
rect 50536 67424 50600 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 19576 66396 19640 66400
rect 19576 66340 19580 66396
rect 19580 66340 19636 66396
rect 19636 66340 19640 66396
rect 19576 66336 19640 66340
rect 19656 66396 19720 66400
rect 19656 66340 19660 66396
rect 19660 66340 19716 66396
rect 19716 66340 19720 66396
rect 19656 66336 19720 66340
rect 19736 66396 19800 66400
rect 19736 66340 19740 66396
rect 19740 66340 19796 66396
rect 19796 66340 19800 66396
rect 19736 66336 19800 66340
rect 19816 66396 19880 66400
rect 19816 66340 19820 66396
rect 19820 66340 19876 66396
rect 19876 66340 19880 66396
rect 19816 66336 19880 66340
rect 50296 66396 50360 66400
rect 50296 66340 50300 66396
rect 50300 66340 50356 66396
rect 50356 66340 50360 66396
rect 50296 66336 50360 66340
rect 50376 66396 50440 66400
rect 50376 66340 50380 66396
rect 50380 66340 50436 66396
rect 50436 66340 50440 66396
rect 50376 66336 50440 66340
rect 50456 66396 50520 66400
rect 50456 66340 50460 66396
rect 50460 66340 50516 66396
rect 50516 66340 50520 66396
rect 50456 66336 50520 66340
rect 50536 66396 50600 66400
rect 50536 66340 50540 66396
rect 50540 66340 50596 66396
rect 50596 66340 50600 66396
rect 50536 66336 50600 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 19576 65308 19640 65312
rect 19576 65252 19580 65308
rect 19580 65252 19636 65308
rect 19636 65252 19640 65308
rect 19576 65248 19640 65252
rect 19656 65308 19720 65312
rect 19656 65252 19660 65308
rect 19660 65252 19716 65308
rect 19716 65252 19720 65308
rect 19656 65248 19720 65252
rect 19736 65308 19800 65312
rect 19736 65252 19740 65308
rect 19740 65252 19796 65308
rect 19796 65252 19800 65308
rect 19736 65248 19800 65252
rect 19816 65308 19880 65312
rect 19816 65252 19820 65308
rect 19820 65252 19876 65308
rect 19876 65252 19880 65308
rect 19816 65248 19880 65252
rect 50296 65308 50360 65312
rect 50296 65252 50300 65308
rect 50300 65252 50356 65308
rect 50356 65252 50360 65308
rect 50296 65248 50360 65252
rect 50376 65308 50440 65312
rect 50376 65252 50380 65308
rect 50380 65252 50436 65308
rect 50436 65252 50440 65308
rect 50376 65248 50440 65252
rect 50456 65308 50520 65312
rect 50456 65252 50460 65308
rect 50460 65252 50516 65308
rect 50516 65252 50520 65308
rect 50456 65248 50520 65252
rect 50536 65308 50600 65312
rect 50536 65252 50540 65308
rect 50540 65252 50596 65308
rect 50596 65252 50600 65308
rect 50536 65248 50600 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 34936 64764 35000 64768
rect 34936 64708 34940 64764
rect 34940 64708 34996 64764
rect 34996 64708 35000 64764
rect 34936 64704 35000 64708
rect 35016 64764 35080 64768
rect 35016 64708 35020 64764
rect 35020 64708 35076 64764
rect 35076 64708 35080 64764
rect 35016 64704 35080 64708
rect 35096 64764 35160 64768
rect 35096 64708 35100 64764
rect 35100 64708 35156 64764
rect 35156 64708 35160 64764
rect 35096 64704 35160 64708
rect 35176 64764 35240 64768
rect 35176 64708 35180 64764
rect 35180 64708 35236 64764
rect 35236 64708 35240 64764
rect 35176 64704 35240 64708
rect 65656 64764 65720 64768
rect 65656 64708 65660 64764
rect 65660 64708 65716 64764
rect 65716 64708 65720 64764
rect 65656 64704 65720 64708
rect 65736 64764 65800 64768
rect 65736 64708 65740 64764
rect 65740 64708 65796 64764
rect 65796 64708 65800 64764
rect 65736 64704 65800 64708
rect 65816 64764 65880 64768
rect 65816 64708 65820 64764
rect 65820 64708 65876 64764
rect 65876 64708 65880 64764
rect 65816 64704 65880 64708
rect 65896 64764 65960 64768
rect 65896 64708 65900 64764
rect 65900 64708 65956 64764
rect 65956 64708 65960 64764
rect 65896 64704 65960 64708
rect 19576 64220 19640 64224
rect 19576 64164 19580 64220
rect 19580 64164 19636 64220
rect 19636 64164 19640 64220
rect 19576 64160 19640 64164
rect 19656 64220 19720 64224
rect 19656 64164 19660 64220
rect 19660 64164 19716 64220
rect 19716 64164 19720 64220
rect 19656 64160 19720 64164
rect 19736 64220 19800 64224
rect 19736 64164 19740 64220
rect 19740 64164 19796 64220
rect 19796 64164 19800 64220
rect 19736 64160 19800 64164
rect 19816 64220 19880 64224
rect 19816 64164 19820 64220
rect 19820 64164 19876 64220
rect 19876 64164 19880 64220
rect 19816 64160 19880 64164
rect 50296 64220 50360 64224
rect 50296 64164 50300 64220
rect 50300 64164 50356 64220
rect 50356 64164 50360 64220
rect 50296 64160 50360 64164
rect 50376 64220 50440 64224
rect 50376 64164 50380 64220
rect 50380 64164 50436 64220
rect 50436 64164 50440 64220
rect 50376 64160 50440 64164
rect 50456 64220 50520 64224
rect 50456 64164 50460 64220
rect 50460 64164 50516 64220
rect 50516 64164 50520 64220
rect 50456 64160 50520 64164
rect 50536 64220 50600 64224
rect 50536 64164 50540 64220
rect 50540 64164 50596 64220
rect 50596 64164 50600 64220
rect 50536 64160 50600 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 34936 63676 35000 63680
rect 34936 63620 34940 63676
rect 34940 63620 34996 63676
rect 34996 63620 35000 63676
rect 34936 63616 35000 63620
rect 35016 63676 35080 63680
rect 35016 63620 35020 63676
rect 35020 63620 35076 63676
rect 35076 63620 35080 63676
rect 35016 63616 35080 63620
rect 35096 63676 35160 63680
rect 35096 63620 35100 63676
rect 35100 63620 35156 63676
rect 35156 63620 35160 63676
rect 35096 63616 35160 63620
rect 35176 63676 35240 63680
rect 35176 63620 35180 63676
rect 35180 63620 35236 63676
rect 35236 63620 35240 63676
rect 35176 63616 35240 63620
rect 65656 63676 65720 63680
rect 65656 63620 65660 63676
rect 65660 63620 65716 63676
rect 65716 63620 65720 63676
rect 65656 63616 65720 63620
rect 65736 63676 65800 63680
rect 65736 63620 65740 63676
rect 65740 63620 65796 63676
rect 65796 63620 65800 63676
rect 65736 63616 65800 63620
rect 65816 63676 65880 63680
rect 65816 63620 65820 63676
rect 65820 63620 65876 63676
rect 65876 63620 65880 63676
rect 65816 63616 65880 63620
rect 65896 63676 65960 63680
rect 65896 63620 65900 63676
rect 65900 63620 65956 63676
rect 65956 63620 65960 63676
rect 65896 63616 65960 63620
rect 19576 63132 19640 63136
rect 19576 63076 19580 63132
rect 19580 63076 19636 63132
rect 19636 63076 19640 63132
rect 19576 63072 19640 63076
rect 19656 63132 19720 63136
rect 19656 63076 19660 63132
rect 19660 63076 19716 63132
rect 19716 63076 19720 63132
rect 19656 63072 19720 63076
rect 19736 63132 19800 63136
rect 19736 63076 19740 63132
rect 19740 63076 19796 63132
rect 19796 63076 19800 63132
rect 19736 63072 19800 63076
rect 19816 63132 19880 63136
rect 19816 63076 19820 63132
rect 19820 63076 19876 63132
rect 19876 63076 19880 63132
rect 19816 63072 19880 63076
rect 50296 63132 50360 63136
rect 50296 63076 50300 63132
rect 50300 63076 50356 63132
rect 50356 63076 50360 63132
rect 50296 63072 50360 63076
rect 50376 63132 50440 63136
rect 50376 63076 50380 63132
rect 50380 63076 50436 63132
rect 50436 63076 50440 63132
rect 50376 63072 50440 63076
rect 50456 63132 50520 63136
rect 50456 63076 50460 63132
rect 50460 63076 50516 63132
rect 50516 63076 50520 63132
rect 50456 63072 50520 63076
rect 50536 63132 50600 63136
rect 50536 63076 50540 63132
rect 50540 63076 50596 63132
rect 50596 63076 50600 63132
rect 50536 63072 50600 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 34936 62588 35000 62592
rect 34936 62532 34940 62588
rect 34940 62532 34996 62588
rect 34996 62532 35000 62588
rect 34936 62528 35000 62532
rect 35016 62588 35080 62592
rect 35016 62532 35020 62588
rect 35020 62532 35076 62588
rect 35076 62532 35080 62588
rect 35016 62528 35080 62532
rect 35096 62588 35160 62592
rect 35096 62532 35100 62588
rect 35100 62532 35156 62588
rect 35156 62532 35160 62588
rect 35096 62528 35160 62532
rect 35176 62588 35240 62592
rect 35176 62532 35180 62588
rect 35180 62532 35236 62588
rect 35236 62532 35240 62588
rect 35176 62528 35240 62532
rect 65656 62588 65720 62592
rect 65656 62532 65660 62588
rect 65660 62532 65716 62588
rect 65716 62532 65720 62588
rect 65656 62528 65720 62532
rect 65736 62588 65800 62592
rect 65736 62532 65740 62588
rect 65740 62532 65796 62588
rect 65796 62532 65800 62588
rect 65736 62528 65800 62532
rect 65816 62588 65880 62592
rect 65816 62532 65820 62588
rect 65820 62532 65876 62588
rect 65876 62532 65880 62588
rect 65816 62528 65880 62532
rect 65896 62588 65960 62592
rect 65896 62532 65900 62588
rect 65900 62532 65956 62588
rect 65956 62532 65960 62588
rect 65896 62528 65960 62532
rect 19576 62044 19640 62048
rect 19576 61988 19580 62044
rect 19580 61988 19636 62044
rect 19636 61988 19640 62044
rect 19576 61984 19640 61988
rect 19656 62044 19720 62048
rect 19656 61988 19660 62044
rect 19660 61988 19716 62044
rect 19716 61988 19720 62044
rect 19656 61984 19720 61988
rect 19736 62044 19800 62048
rect 19736 61988 19740 62044
rect 19740 61988 19796 62044
rect 19796 61988 19800 62044
rect 19736 61984 19800 61988
rect 19816 62044 19880 62048
rect 19816 61988 19820 62044
rect 19820 61988 19876 62044
rect 19876 61988 19880 62044
rect 19816 61984 19880 61988
rect 50296 62044 50360 62048
rect 50296 61988 50300 62044
rect 50300 61988 50356 62044
rect 50356 61988 50360 62044
rect 50296 61984 50360 61988
rect 50376 62044 50440 62048
rect 50376 61988 50380 62044
rect 50380 61988 50436 62044
rect 50436 61988 50440 62044
rect 50376 61984 50440 61988
rect 50456 62044 50520 62048
rect 50456 61988 50460 62044
rect 50460 61988 50516 62044
rect 50516 61988 50520 62044
rect 50456 61984 50520 61988
rect 50536 62044 50600 62048
rect 50536 61988 50540 62044
rect 50540 61988 50596 62044
rect 50596 61988 50600 62044
rect 50536 61984 50600 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 65656 61500 65720 61504
rect 65656 61444 65660 61500
rect 65660 61444 65716 61500
rect 65716 61444 65720 61500
rect 65656 61440 65720 61444
rect 65736 61500 65800 61504
rect 65736 61444 65740 61500
rect 65740 61444 65796 61500
rect 65796 61444 65800 61500
rect 65736 61440 65800 61444
rect 65816 61500 65880 61504
rect 65816 61444 65820 61500
rect 65820 61444 65876 61500
rect 65876 61444 65880 61500
rect 65816 61440 65880 61444
rect 65896 61500 65960 61504
rect 65896 61444 65900 61500
rect 65900 61444 65956 61500
rect 65956 61444 65960 61500
rect 65896 61440 65960 61444
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 65656 60412 65720 60416
rect 65656 60356 65660 60412
rect 65660 60356 65716 60412
rect 65716 60356 65720 60412
rect 65656 60352 65720 60356
rect 65736 60412 65800 60416
rect 65736 60356 65740 60412
rect 65740 60356 65796 60412
rect 65796 60356 65800 60412
rect 65736 60352 65800 60356
rect 65816 60412 65880 60416
rect 65816 60356 65820 60412
rect 65820 60356 65876 60412
rect 65876 60356 65880 60412
rect 65816 60352 65880 60356
rect 65896 60412 65960 60416
rect 65896 60356 65900 60412
rect 65900 60356 65956 60412
rect 65956 60356 65960 60412
rect 65896 60352 65960 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 65656 59324 65720 59328
rect 65656 59268 65660 59324
rect 65660 59268 65716 59324
rect 65716 59268 65720 59324
rect 65656 59264 65720 59268
rect 65736 59324 65800 59328
rect 65736 59268 65740 59324
rect 65740 59268 65796 59324
rect 65796 59268 65800 59324
rect 65736 59264 65800 59268
rect 65816 59324 65880 59328
rect 65816 59268 65820 59324
rect 65820 59268 65876 59324
rect 65876 59268 65880 59324
rect 65816 59264 65880 59268
rect 65896 59324 65960 59328
rect 65896 59268 65900 59324
rect 65900 59268 65956 59324
rect 65956 59268 65960 59324
rect 65896 59264 65960 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 65656 58236 65720 58240
rect 65656 58180 65660 58236
rect 65660 58180 65716 58236
rect 65716 58180 65720 58236
rect 65656 58176 65720 58180
rect 65736 58236 65800 58240
rect 65736 58180 65740 58236
rect 65740 58180 65796 58236
rect 65796 58180 65800 58236
rect 65736 58176 65800 58180
rect 65816 58236 65880 58240
rect 65816 58180 65820 58236
rect 65820 58180 65876 58236
rect 65876 58180 65880 58236
rect 65816 58176 65880 58180
rect 65896 58236 65960 58240
rect 65896 58180 65900 58236
rect 65900 58180 65956 58236
rect 65956 58180 65960 58236
rect 65896 58176 65960 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 66944 4528 67504
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 65856 4528 66880
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 67488 19888 67504
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 66400 19888 67424
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 65312 19888 66336
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 64224 19888 65248
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 63136 19888 64160
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 62048 19888 63072
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 60960 19888 61984
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 66944 35248 67504
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 65856 35248 66880
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 64768 35248 65792
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 63680 35248 64704
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 62592 35248 63616
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 61504 35248 62528
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 67488 50608 67504
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 66400 50608 67424
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 65312 50608 66336
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 64224 50608 65248
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 63136 50608 64160
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 62048 50608 63072
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 60960 50608 61984
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 66944 65968 67504
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 65856 65968 66880
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 64768 65968 65792
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 63680 65968 64704
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 62592 65968 63616
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 61504 65968 62528
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 60416 65968 61440
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 59328 65968 60352
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 58240 65968 59264
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 57152 65968 58176
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__or4b_1  _0611_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34316 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0612_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0613_
timestamp 1688980957
transform -1 0 34040 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0614_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0615_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0616_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33396 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0617_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35144 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0618_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34132 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0619_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35972 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0620_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31188 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0621_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36156 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0622_
timestamp 1688980957
transform 1 0 36616 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0623_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35328 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0624_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35420 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0625_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0626_
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1688980957
transform 1 0 30820 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0628_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0629_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34040 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0630_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0631_
timestamp 1688980957
transform 1 0 34776 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0632_
timestamp 1688980957
transform -1 0 35236 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1688980957
transform 1 0 35420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0634_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33396 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0635_
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0636_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32292 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0637_
timestamp 1688980957
transform 1 0 32660 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0638_
timestamp 1688980957
transform 1 0 32200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0639_
timestamp 1688980957
transform -1 0 31648 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0640_
timestamp 1688980957
transform -1 0 31924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0641_
timestamp 1688980957
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform 1 0 30912 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1688980957
transform 1 0 30728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0644_
timestamp 1688980957
transform 1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0645_
timestamp 1688980957
transform 1 0 21620 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _0646_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0647_
timestamp 1688980957
transform 1 0 16836 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0648_
timestamp 1688980957
transform 1 0 22632 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0649_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0650_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0651_
timestamp 1688980957
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0652_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22264 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0653_
timestamp 1688980957
transform 1 0 25944 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0654_
timestamp 1688980957
transform -1 0 27140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0655_
timestamp 1688980957
transform -1 0 26864 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0656_
timestamp 1688980957
transform -1 0 26772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0657_
timestamp 1688980957
transform -1 0 27232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0658_
timestamp 1688980957
transform -1 0 26404 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0659_
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0660_
timestamp 1688980957
transform 1 0 26404 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0661_
timestamp 1688980957
transform 1 0 27324 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0662_
timestamp 1688980957
transform -1 0 29256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0663_
timestamp 1688980957
transform -1 0 28244 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0664_
timestamp 1688980957
transform 1 0 29348 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1688980957
transform -1 0 28244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0666_
timestamp 1688980957
transform 1 0 28244 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0667_
timestamp 1688980957
transform 1 0 28520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0668_
timestamp 1688980957
transform -1 0 26864 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0669_
timestamp 1688980957
transform 1 0 26956 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0670_
timestamp 1688980957
transform -1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0671_
timestamp 1688980957
transform -1 0 28244 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1688980957
transform -1 0 27784 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0673_
timestamp 1688980957
transform 1 0 28336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0674_
timestamp 1688980957
transform 1 0 27692 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1688980957
transform -1 0 26128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0676_
timestamp 1688980957
transform -1 0 25208 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0677_
timestamp 1688980957
transform 1 0 25116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0678_
timestamp 1688980957
transform -1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0679_
timestamp 1688980957
transform -1 0 26036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0680_
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0681_
timestamp 1688980957
transform -1 0 25760 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0682_
timestamp 1688980957
transform 1 0 24472 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0683_
timestamp 1688980957
transform 1 0 23736 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1688980957
transform 1 0 23092 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1688980957
transform -1 0 23184 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0686_
timestamp 1688980957
transform -1 0 24196 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0687_
timestamp 1688980957
transform -1 0 22816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0688_
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0689_
timestamp 1688980957
transform -1 0 23000 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0690_
timestamp 1688980957
transform 1 0 22632 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0691_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23460 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0692_
timestamp 1688980957
transform -1 0 23368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0693_
timestamp 1688980957
transform 1 0 23184 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0694_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21896 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1688980957
transform 1 0 17020 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0696_
timestamp 1688980957
transform -1 0 19136 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1688980957
transform 1 0 18676 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0698_
timestamp 1688980957
transform -1 0 20516 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0699_
timestamp 1688980957
transform -1 0 20056 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0700_
timestamp 1688980957
transform -1 0 20516 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0701_
timestamp 1688980957
transform 1 0 20332 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0702_
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0703_
timestamp 1688980957
transform -1 0 21620 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0704_
timestamp 1688980957
transform 1 0 20148 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1688980957
transform -1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0706_
timestamp 1688980957
transform -1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0707_
timestamp 1688980957
transform -1 0 22264 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0708_
timestamp 1688980957
transform -1 0 19136 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0710_
timestamp 1688980957
transform -1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0711_
timestamp 1688980957
transform -1 0 19596 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0712_
timestamp 1688980957
transform 1 0 17848 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1688980957
transform -1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0714_
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0715_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0716_
timestamp 1688980957
transform 1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0717_
timestamp 1688980957
transform -1 0 17388 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0718_
timestamp 1688980957
transform 1 0 18032 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0719_
timestamp 1688980957
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0720_
timestamp 1688980957
transform -1 0 18860 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 1688980957
transform 1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 1688980957
transform -1 0 16468 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1688980957
transform -1 0 16192 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1688980957
transform 1 0 10948 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1688980957
transform -1 0 15548 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0727_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12052 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1688980957
transform -1 0 13340 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0729_
timestamp 1688980957
transform -1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0730_
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1688980957
transform -1 0 13248 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0732_
timestamp 1688980957
transform 1 0 15180 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1688980957
transform -1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0734_
timestamp 1688980957
transform -1 0 23460 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1688980957
transform -1 0 22816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 1688980957
transform 1 0 22264 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0737_
timestamp 1688980957
transform -1 0 21068 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0738_
timestamp 1688980957
transform 1 0 21804 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0739_
timestamp 1688980957
transform -1 0 21804 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0740_
timestamp 1688980957
transform -1 0 21620 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0741_
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1688980957
transform 1 0 19688 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 1688980957
transform 1 0 19504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0744_
timestamp 1688980957
transform -1 0 21712 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0745_
timestamp 1688980957
transform 1 0 19780 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0746_
timestamp 1688980957
transform 1 0 21988 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0747_
timestamp 1688980957
transform 1 0 23184 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0748_
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0749_
timestamp 1688980957
transform -1 0 22448 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0750_
timestamp 1688980957
transform -1 0 22908 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0751_
timestamp 1688980957
transform 1 0 23000 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0752_
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0753_
timestamp 1688980957
transform 1 0 22172 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1688980957
transform 1 0 25392 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0755_
timestamp 1688980957
transform 1 0 25668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0756_
timestamp 1688980957
transform -1 0 25208 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0757_
timestamp 1688980957
transform -1 0 25392 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0758_
timestamp 1688980957
transform -1 0 25116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1688980957
transform -1 0 25668 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0760_
timestamp 1688980957
transform -1 0 24748 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0761_
timestamp 1688980957
transform 1 0 20700 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0762_
timestamp 1688980957
transform 1 0 20424 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0763_
timestamp 1688980957
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1688980957
transform 1 0 12696 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0765_
timestamp 1688980957
transform -1 0 13248 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1688980957
transform -1 0 14352 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0767_
timestamp 1688980957
transform -1 0 11408 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0768_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11408 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0769_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0770_
timestamp 1688980957
transform 1 0 12052 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0771_
timestamp 1688980957
transform 1 0 13156 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0772_
timestamp 1688980957
transform -1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0773_
timestamp 1688980957
transform 1 0 10488 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0774_
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0776_
timestamp 1688980957
transform 1 0 13616 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0778_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _0779_
timestamp 1688980957
transform -1 0 13340 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0780_
timestamp 1688980957
transform -1 0 12696 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1688980957
transform 1 0 12328 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0782_
timestamp 1688980957
transform -1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0783_
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0784_
timestamp 1688980957
transform 1 0 11960 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0785_
timestamp 1688980957
transform -1 0 11408 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0786_
timestamp 1688980957
transform -1 0 10580 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0787_
timestamp 1688980957
transform 1 0 11316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0788_
timestamp 1688980957
transform -1 0 11316 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1688980957
transform 1 0 11592 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0790_
timestamp 1688980957
transform -1 0 11592 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0791_
timestamp 1688980957
transform -1 0 11132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1688980957
transform -1 0 11408 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0793_
timestamp 1688980957
transform 1 0 10212 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0794_
timestamp 1688980957
transform 1 0 9752 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0795_
timestamp 1688980957
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0796_
timestamp 1688980957
transform 1 0 11868 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0797_
timestamp 1688980957
transform -1 0 11776 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0798_
timestamp 1688980957
transform 1 0 11592 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0799_
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1688980957
transform 1 0 9200 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 1688980957
transform 1 0 8464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0802_
timestamp 1688980957
transform -1 0 12328 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0803_
timestamp 1688980957
transform -1 0 11316 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0804_
timestamp 1688980957
transform -1 0 10120 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0805_
timestamp 1688980957
transform -1 0 10120 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1688980957
transform -1 0 11960 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0807_
timestamp 1688980957
transform 1 0 11224 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0808_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0809_
timestamp 1688980957
transform 1 0 10212 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0811_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0812_
timestamp 1688980957
transform -1 0 10212 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1688980957
transform -1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1688980957
transform -1 0 11592 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0816_
timestamp 1688980957
transform 1 0 10212 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1688980957
transform 1 0 9016 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0818_
timestamp 1688980957
transform 1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1688980957
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0820_
timestamp 1688980957
transform -1 0 10948 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0821_
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0822_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0823_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9384 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0825_
timestamp 1688980957
transform 1 0 12512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0826_
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0828_
timestamp 1688980957
transform -1 0 12788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0830_
timestamp 1688980957
transform 1 0 10672 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0831_
timestamp 1688980957
transform 1 0 29900 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1688980957
transform -1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1688980957
transform -1 0 31004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0834_
timestamp 1688980957
transform -1 0 30728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 1688980957
transform 1 0 25392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0836_
timestamp 1688980957
transform 1 0 24564 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0837_
timestamp 1688980957
transform 1 0 25300 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1688980957
transform 1 0 13984 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0839_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18400 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0840_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0841_
timestamp 1688980957
transform 1 0 17664 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1688980957
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0843_
timestamp 1688980957
transform 1 0 27508 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0844_
timestamp 1688980957
transform 1 0 26312 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0845_
timestamp 1688980957
transform 1 0 26404 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0846_
timestamp 1688980957
transform 1 0 28060 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0847_
timestamp 1688980957
transform 1 0 17572 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0848_
timestamp 1688980957
transform -1 0 18676 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0851_
timestamp 1688980957
transform 1 0 18216 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1688980957
transform 1 0 26956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0853_
timestamp 1688980957
transform -1 0 26404 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0854_
timestamp 1688980957
transform 1 0 22448 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0855_
timestamp 1688980957
transform 1 0 21804 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0856_
timestamp 1688980957
transform 1 0 21344 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0857_
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0858_
timestamp 1688980957
transform 1 0 23460 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0859_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0860_
timestamp 1688980957
transform -1 0 27876 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1688980957
transform -1 0 28244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1688980957
transform 1 0 20700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0864_
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1688980957
transform -1 0 23276 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0866_
timestamp 1688980957
transform -1 0 22908 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0868_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1688980957
transform -1 0 34224 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0870_
timestamp 1688980957
transform 1 0 23552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0871_
timestamp 1688980957
transform 1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0872_
timestamp 1688980957
transform 1 0 23368 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0873_
timestamp 1688980957
transform 1 0 19044 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0874_
timestamp 1688980957
transform -1 0 14996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0875_
timestamp 1688980957
transform -1 0 21712 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0876_
timestamp 1688980957
transform 1 0 20516 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0877_
timestamp 1688980957
transform 1 0 20792 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1688980957
transform -1 0 37444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0879_
timestamp 1688980957
transform 1 0 30728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0880_
timestamp 1688980957
transform 1 0 30452 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0881_
timestamp 1688980957
transform 1 0 31556 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0882_
timestamp 1688980957
transform 1 0 35328 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0883_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27692 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0884_
timestamp 1688980957
transform 1 0 28152 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0885_
timestamp 1688980957
transform -1 0 32016 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0886_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30912 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0887_
timestamp 1688980957
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0888_
timestamp 1688980957
transform -1 0 29808 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 1688980957
transform -1 0 29440 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0890_
timestamp 1688980957
transform 1 0 28888 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0891_
timestamp 1688980957
transform 1 0 29348 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1688980957
transform 1 0 28704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1688980957
transform -1 0 30728 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _0894_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29624 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0895_
timestamp 1688980957
transform -1 0 30176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0896_
timestamp 1688980957
transform 1 0 20792 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0897_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27876 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0898_
timestamp 1688980957
transform -1 0 36708 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1688980957
transform -1 0 36248 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_2  _0900_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 37168 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0901_
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 1688980957
transform -1 0 35328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0903_
timestamp 1688980957
transform 1 0 34868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1688980957
transform 1 0 33764 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1688980957
transform 1 0 34224 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0906_
timestamp 1688980957
transform -1 0 35788 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0907_
timestamp 1688980957
transform -1 0 35236 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0908_
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0909_
timestamp 1688980957
transform -1 0 35788 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0910_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36156 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0911_
timestamp 1688980957
transform -1 0 26128 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1688980957
transform -1 0 26036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0913_
timestamp 1688980957
transform -1 0 15824 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1688980957
transform -1 0 15456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0915_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 1688980957
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1688980957
transform -1 0 17848 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0918_
timestamp 1688980957
transform 1 0 16652 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 1688980957
transform 1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0920_
timestamp 1688980957
transform 1 0 18768 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0921_
timestamp 1688980957
transform 1 0 19964 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0922_
timestamp 1688980957
transform -1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0923_
timestamp 1688980957
transform -1 0 16560 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0924_
timestamp 1688980957
transform -1 0 19228 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1688980957
transform -1 0 19136 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1688980957
transform 1 0 23276 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0927_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0928_
timestamp 1688980957
transform 1 0 17480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp 1688980957
transform -1 0 18216 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0930_
timestamp 1688980957
transform 1 0 17848 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1688980957
transform -1 0 18584 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0932_
timestamp 1688980957
transform -1 0 22540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0933_
timestamp 1688980957
transform -1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0934_
timestamp 1688980957
transform -1 0 23736 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0935_
timestamp 1688980957
transform 1 0 23000 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0936_
timestamp 1688980957
transform -1 0 24748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0937_
timestamp 1688980957
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 1688980957
transform 1 0 26036 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1688980957
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0941_
timestamp 1688980957
transform 1 0 19596 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0942_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20056 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1688980957
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0944_
timestamp 1688980957
transform 1 0 24564 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp 1688980957
transform 1 0 22448 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 1688980957
transform 1 0 21620 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0947_
timestamp 1688980957
transform 1 0 14904 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 1688980957
transform 1 0 13064 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0949_
timestamp 1688980957
transform -1 0 13156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 1688980957
transform 1 0 13156 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_1  _0951_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12880 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0952_
timestamp 1688980957
transform 1 0 12604 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0953_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13064 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0954_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0955_
timestamp 1688980957
transform 1 0 24932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1688980957
transform -1 0 25760 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0957_
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0958_
timestamp 1688980957
transform 1 0 25576 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0959_
timestamp 1688980957
transform -1 0 25852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0960_
timestamp 1688980957
transform 1 0 24564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0961_
timestamp 1688980957
transform 1 0 22264 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0962_
timestamp 1688980957
transform -1 0 27508 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1688980957
transform 1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1688980957
transform -1 0 26772 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0965_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25576 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0966_
timestamp 1688980957
transform -1 0 26036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0967_
timestamp 1688980957
transform -1 0 25484 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0968_
timestamp 1688980957
transform -1 0 25576 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _0969_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1688980957
transform 1 0 34224 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1688980957
transform 1 0 32568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0972_
timestamp 1688980957
transform -1 0 31924 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0973_
timestamp 1688980957
transform -1 0 35328 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 1688980957
transform -1 0 32752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0975_
timestamp 1688980957
transform -1 0 33580 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0976_
timestamp 1688980957
transform 1 0 32476 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _0977_
timestamp 1688980957
transform 1 0 32200 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1688980957
transform -1 0 19688 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0979_
timestamp 1688980957
transform -1 0 18216 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _0980_
timestamp 1688980957
transform 1 0 18768 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0981_
timestamp 1688980957
transform 1 0 18124 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0982_
timestamp 1688980957
transform -1 0 18768 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0983_
timestamp 1688980957
transform -1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0984_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23092 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0985_
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _0986_
timestamp 1688980957
transform 1 0 13248 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1688980957
transform 1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0988_
timestamp 1688980957
transform -1 0 13156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0989_
timestamp 1688980957
transform 1 0 11592 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _0990_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0991_
timestamp 1688980957
transform 1 0 13248 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _0992_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12512 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1688980957
transform 1 0 10488 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1688980957
transform 1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 1688980957
transform 1 0 14628 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1688980957
transform 1 0 14352 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0997_
timestamp 1688980957
transform 1 0 19596 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1688980957
transform -1 0 19504 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp 1688980957
transform -1 0 20056 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1688980957
transform 1 0 19688 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 1688980957
transform 1 0 27416 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1688980957
transform -1 0 26864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1003_
timestamp 1688980957
transform -1 0 30452 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1688980957
transform 1 0 29808 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1688980957
transform 1 0 16100 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1688980957
transform 1 0 18032 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1007_
timestamp 1688980957
transform 1 0 17480 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1688980957
transform 1 0 17940 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1009_
timestamp 1688980957
transform 1 0 25208 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1688980957
transform 1 0 25300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _1011_
timestamp 1688980957
transform 1 0 24932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1012_
timestamp 1688980957
transform 1 0 17572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1013_
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1688980957
transform -1 0 18952 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1015_
timestamp 1688980957
transform -1 0 17388 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1688980957
transform -1 0 16560 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1017_
timestamp 1688980957
transform -1 0 19780 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1688980957
transform -1 0 18768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1019_
timestamp 1688980957
transform 1 0 20332 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1688980957
transform -1 0 22080 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1021_
timestamp 1688980957
transform 1 0 28244 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1688980957
transform 1 0 29440 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1023_
timestamp 1688980957
transform -1 0 30452 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1688980957
transform -1 0 29440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1025_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1688980957
transform 1 0 13800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1027_
timestamp 1688980957
transform 1 0 20516 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1028_
timestamp 1688980957
transform -1 0 24840 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1688980957
transform -1 0 24012 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 1688980957
transform 1 0 23828 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1688980957
transform -1 0 24656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1032_
timestamp 1688980957
transform 1 0 20332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1033_
timestamp 1688980957
transform 1 0 27140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1034_
timestamp 1688980957
transform 1 0 30452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1035_
timestamp 1688980957
transform -1 0 36156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1036_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1037_
timestamp 1688980957
transform 1 0 32568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1038_
timestamp 1688980957
transform 1 0 33488 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1039_
timestamp 1688980957
transform -1 0 33304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1040_
timestamp 1688980957
transform -1 0 32936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1041_
timestamp 1688980957
transform 1 0 34868 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1042_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1043_
timestamp 1688980957
transform -1 0 36156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1044_
timestamp 1688980957
transform 1 0 37904 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1045_
timestamp 1688980957
transform -1 0 38364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1046_
timestamp 1688980957
transform 1 0 36340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1047_
timestamp 1688980957
transform 1 0 36984 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1688980957
transform 1 0 35052 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1049_
timestamp 1688980957
transform -1 0 35696 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1050_
timestamp 1688980957
transform -1 0 34592 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1051_
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1052_
timestamp 1688980957
transform -1 0 35696 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1053_
timestamp 1688980957
transform -1 0 37536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1054_
timestamp 1688980957
transform -1 0 36340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1055_
timestamp 1688980957
transform 1 0 35788 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1056_
timestamp 1688980957
transform 1 0 34960 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1057_
timestamp 1688980957
transform 1 0 35696 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1058_
timestamp 1688980957
transform -1 0 36800 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1059_
timestamp 1688980957
transform 1 0 36524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1060_
timestamp 1688980957
transform -1 0 36616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1061_
timestamp 1688980957
transform -1 0 36984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1062_
timestamp 1688980957
transform 1 0 33672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1063_
timestamp 1688980957
transform -1 0 31464 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1688980957
transform 1 0 29624 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1065_
timestamp 1688980957
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1066_
timestamp 1688980957
transform 1 0 30268 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1067_
timestamp 1688980957
transform -1 0 28796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 1688980957
transform -1 0 28704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1069_
timestamp 1688980957
transform 1 0 28704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 1688980957
transform -1 0 29992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1071_
timestamp 1688980957
transform 1 0 30268 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1072_
timestamp 1688980957
transform -1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1073_
timestamp 1688980957
transform 1 0 26772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1074_
timestamp 1688980957
transform -1 0 32016 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1075_
timestamp 1688980957
transform -1 0 26404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1076_
timestamp 1688980957
transform 1 0 24564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1077_
timestamp 1688980957
transform 1 0 25208 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1078_
timestamp 1688980957
transform -1 0 31096 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1079_
timestamp 1688980957
transform -1 0 31924 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1080_
timestamp 1688980957
transform 1 0 26680 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1081_
timestamp 1688980957
transform 1 0 30268 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1082_
timestamp 1688980957
transform -1 0 31096 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1083_
timestamp 1688980957
transform 1 0 29900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1084_
timestamp 1688980957
transform -1 0 34132 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1085_
timestamp 1688980957
transform -1 0 31832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1086_
timestamp 1688980957
transform 1 0 31004 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1087_
timestamp 1688980957
transform 1 0 32384 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1088_
timestamp 1688980957
transform 1 0 34132 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1089_
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1090_
timestamp 1688980957
transform -1 0 33028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1091_
timestamp 1688980957
transform 1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _1092_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32844 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1688980957
transform -1 0 31280 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1094_
timestamp 1688980957
transform 1 0 31280 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1095_
timestamp 1688980957
transform -1 0 32476 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1096_
timestamp 1688980957
transform 1 0 31924 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1097_
timestamp 1688980957
transform -1 0 33120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1098_
timestamp 1688980957
transform -1 0 33580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1099_
timestamp 1688980957
transform 1 0 32568 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1688980957
transform -1 0 32568 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1101_
timestamp 1688980957
transform 1 0 31280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1102_
timestamp 1688980957
transform -1 0 32200 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1103_
timestamp 1688980957
transform 1 0 30360 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1104_
timestamp 1688980957
transform 1 0 29900 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1105_
timestamp 1688980957
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1106_
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1107_
timestamp 1688980957
transform -1 0 28336 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1108_
timestamp 1688980957
transform 1 0 27600 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1688980957
transform -1 0 28612 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1110_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27600 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 1688980957
transform -1 0 26772 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1112_
timestamp 1688980957
transform -1 0 28060 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1113_
timestamp 1688980957
transform 1 0 27508 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1114_
timestamp 1688980957
transform -1 0 27692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1688980957
transform -1 0 26864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1116_
timestamp 1688980957
transform -1 0 27876 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1117_
timestamp 1688980957
transform -1 0 27416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1118_
timestamp 1688980957
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1119_
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1120_
timestamp 1688980957
transform 1 0 28612 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  _1121_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33212 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1123_
timestamp 1688980957
transform -1 0 31556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1124_
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1688980957
transform 1 0 29992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1688980957
transform -1 0 13340 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1688980957
transform -1 0 11776 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1688980957
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1688980957
transform 1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1688980957
transform 1 0 9292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1688980957
transform 1 0 8464 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1688980957
transform -1 0 8740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1688980957
transform 1 0 8464 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1134_
timestamp 1688980957
transform -1 0 15732 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1688980957
transform -1 0 9660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1688980957
transform -1 0 11132 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1137_
timestamp 1688980957
transform -1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1138_
timestamp 1688980957
transform -1 0 15272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1688980957
transform -1 0 15916 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1140_
timestamp 1688980957
transform 1 0 14352 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1688980957
transform 1 0 14628 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1688980957
transform -1 0 8832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 1688980957
transform 1 0 11592 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1688980957
transform 1 0 9476 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1688980957
transform 1 0 9292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1688980957
transform 1 0 11040 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1149_
timestamp 1688980957
transform -1 0 20608 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1150_
timestamp 1688980957
transform -1 0 14352 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1688980957
transform -1 0 16468 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1152_
timestamp 1688980957
transform -1 0 16560 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1153_
timestamp 1688980957
transform 1 0 14444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 1688980957
transform -1 0 15824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1155_
timestamp 1688980957
transform 1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1156_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1157_
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1158_
timestamp 1688980957
transform -1 0 15272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1159_
timestamp 1688980957
transform -1 0 14536 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1688980957
transform 1 0 21252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1688980957
transform 1 0 20976 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1163_
timestamp 1688980957
transform 1 0 24748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1688980957
transform 1 0 22632 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1688980957
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1688980957
transform -1 0 22080 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1167_
timestamp 1688980957
transform 1 0 20424 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1688980957
transform 1 0 18676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1688980957
transform -1 0 19504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1688980957
transform 1 0 19504 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1171_
timestamp 1688980957
transform 1 0 23000 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1172_
timestamp 1688980957
transform -1 0 20424 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1688980957
transform 1 0 23184 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1174_
timestamp 1688980957
transform -1 0 24104 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1176_
timestamp 1688980957
transform -1 0 17204 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1177_
timestamp 1688980957
transform -1 0 15272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1688980957
transform 1 0 14720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1179_
timestamp 1688980957
transform 1 0 14168 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1688980957
transform 1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1688980957
transform -1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1688980957
transform -1 0 16560 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1688980957
transform -1 0 16100 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1186_
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1688980957
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1688980957
transform -1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1688980957
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190_
timestamp 1688980957
transform -1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1191_
timestamp 1688980957
transform -1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1192_
timestamp 1688980957
transform -1 0 18308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1688980957
transform 1 0 20516 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1194_
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1195_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1196_
timestamp 1688980957
transform -1 0 24288 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1197_
timestamp 1688980957
transform 1 0 26404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198_
timestamp 1688980957
transform -1 0 25484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1199_
timestamp 1688980957
transform -1 0 25668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1688980957
transform 1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1688980957
transform 1 0 23368 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1688980957
transform 1 0 23552 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1203_
timestamp 1688980957
transform -1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1688980957
transform 1 0 22724 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1205_
timestamp 1688980957
transform 1 0 23184 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1206_
timestamp 1688980957
transform 1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1207_
timestamp 1688980957
transform -1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1208_
timestamp 1688980957
transform -1 0 29808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp 1688980957
transform -1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1688980957
transform -1 0 29348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1211_
timestamp 1688980957
transform -1 0 27508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1212_
timestamp 1688980957
transform -1 0 23920 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1688980957
transform 1 0 17572 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1688980957
transform -1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1215_
timestamp 1688980957
transform -1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1216_
timestamp 1688980957
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1217_
timestamp 1688980957
transform -1 0 28520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1218_
timestamp 1688980957
transform -1 0 31280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1219_
timestamp 1688980957
transform 1 0 30360 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1220_
timestamp 1688980957
transform 1 0 31464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1221_
timestamp 1688980957
transform -1 0 36064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1222_
timestamp 1688980957
transform 1 0 36708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1223_
timestamp 1688980957
transform 1 0 33028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1688980957
transform -1 0 34592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1688980957
transform 1 0 36248 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1226_
timestamp 1688980957
transform -1 0 32016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1227_
timestamp 1688980957
transform 1 0 30360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1228_
timestamp 1688980957
transform -1 0 28704 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1229_
timestamp 1688980957
transform -1 0 29992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1230_
timestamp 1688980957
transform -1 0 31188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1231_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31924 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1232_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19136 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp 1688980957
transform -1 0 19136 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 1688980957
transform -1 0 17664 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp 1688980957
transform -1 0 19780 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 1688980957
transform 1 0 16652 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp 1688980957
transform 1 0 19504 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp 1688980957
transform -1 0 26404 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1688980957
transform 1 0 22816 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1688980957
transform 1 0 20976 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1688980957
transform -1 0 25392 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1688980957
transform 1 0 24748 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 1688980957
transform 1 0 35604 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1688980957
transform 1 0 32016 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1688980957
transform 1 0 32936 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1688980957
transform 1 0 36156 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1688980957
transform 1 0 33764 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1688980957
transform 1 0 35696 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1688980957
transform 1 0 34224 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1688980957
transform 1 0 36984 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1688980957
transform 1 0 36616 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1688980957
transform 1 0 31464 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1688980957
transform 1 0 27508 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 1688980957
transform 1 0 27784 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1688980957
transform -1 0 31004 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 1688980957
transform -1 0 32016 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1688980957
transform 1 0 25300 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1688980957
transform -1 0 25208 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1688980957
transform 1 0 31372 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1688980957
transform -1 0 28428 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1688980957
transform 1 0 24840 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1688980957
transform -1 0 28060 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1688980957
transform 1 0 25392 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1688980957
transform 1 0 26404 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1688980957
transform 1 0 30360 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1688980957
transform 1 0 31832 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1688980957
transform -1 0 34500 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1688980957
transform -1 0 33948 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1688980957
transform 1 0 32568 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1688980957
transform 1 0 29900 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp 1688980957
transform -1 0 29164 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1688980957
transform 1 0 26036 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp 1688980957
transform 1 0 26036 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1688980957
transform 1 0 26128 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1688980957
transform 1 0 27968 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1280_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25024 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1281_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34224 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1688980957
transform 1 0 34960 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1688980957
transform -1 0 13984 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1286_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1688980957
transform 1 0 33396 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1688980957
transform 1 0 22816 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1688980957
transform -1 0 19964 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1688980957
transform -1 0 31004 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1688980957
transform 1 0 27232 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1688980957
transform -1 0 31280 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1688980957
transform -1 0 29440 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1688980957
transform 1 0 33396 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1688980957
transform 1 0 17020 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1688980957
transform 1 0 15088 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1688980957
transform -1 0 17664 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1688980957
transform -1 0 17480 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1688980957
transform 1 0 17572 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1688980957
transform -1 0 18032 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1304_
timestamp 1688980957
transform 1 0 28980 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1305_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1306_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10304 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1307_
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1308_
timestamp 1688980957
transform 1 0 11960 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1309_
timestamp 1688980957
transform 1 0 8372 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1310_
timestamp 1688980957
transform 1 0 7544 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1311_
timestamp 1688980957
transform 1 0 6992 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 1688980957
transform 1 0 7728 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 1688980957
transform 1 0 9568 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1688980957
transform -1 0 15180 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1688980957
transform -1 0 15548 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1317_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1318_
timestamp 1688980957
transform 1 0 7912 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1319_
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1320_
timestamp 1688980957
transform -1 0 11040 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1321_
timestamp 1688980957
transform 1 0 7912 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1322_
timestamp 1688980957
transform 1 0 7912 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1323_
timestamp 1688980957
transform 1 0 8280 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1324_
timestamp 1688980957
transform 1 0 10120 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1325_
timestamp 1688980957
transform 1 0 12144 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1326_
timestamp 1688980957
transform 1 0 13984 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1688980957
transform 1 0 13984 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1688980957
transform -1 0 16928 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1688980957
transform 1 0 14536 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _1330_
timestamp 1688980957
transform 1 0 13156 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1331_
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1332_
timestamp 1688980957
transform 1 0 20056 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1333_
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1334_
timestamp 1688980957
transform -1 0 25760 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1335_
timestamp 1688980957
transform 1 0 22172 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1336_
timestamp 1688980957
transform 1 0 23644 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 1688980957
transform 1 0 20424 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1338_
timestamp 1688980957
transform 1 0 17848 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1339_
timestamp 1688980957
transform 1 0 18124 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1340_
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1688980957
transform 1 0 19596 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1688980957
transform -1 0 23368 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1343_
timestamp 1688980957
transform 1 0 15272 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1688980957
transform 1 0 14536 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1688980957
transform -1 0 14720 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1688980957
transform 1 0 21344 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1688980957
transform 1 0 19780 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1688980957
transform -1 0 19136 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1688980957
transform -1 0 22632 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1350_
timestamp 1688980957
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1351_
timestamp 1688980957
transform 1 0 19228 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1352_
timestamp 1688980957
transform 1 0 20056 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1353_
timestamp 1688980957
transform 1 0 15548 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1354_
timestamp 1688980957
transform 1 0 14628 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1355_
timestamp 1688980957
transform 1 0 15364 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1356_
timestamp 1688980957
transform 1 0 14628 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1357_
timestamp 1688980957
transform 1 0 17296 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1358_
timestamp 1688980957
transform 1 0 19780 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1359_
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1360_
timestamp 1688980957
transform 1 0 20516 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1361_
timestamp 1688980957
transform 1 0 19136 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1688980957
transform 1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1688980957
transform -1 0 20332 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _1364_
timestamp 1688980957
transform 1 0 23000 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1688980957
transform -1 0 25760 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1688980957
transform 1 0 24564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1367_
timestamp 1688980957
transform -1 0 25116 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1368_
timestamp 1688980957
transform 1 0 22356 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1369_
timestamp 1688980957
transform 1 0 22724 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1370_
timestamp 1688980957
transform 1 0 22172 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1371_
timestamp 1688980957
transform 1 0 21896 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1372_
timestamp 1688980957
transform -1 0 26864 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1373_
timestamp 1688980957
transform 1 0 27416 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1374_
timestamp 1688980957
transform 1 0 27508 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1375_
timestamp 1688980957
transform 1 0 28888 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1376_
timestamp 1688980957
transform 1 0 27232 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1378_
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1688980957
transform 1 0 16560 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1688980957
transform 1 0 15088 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1381_
timestamp 1688980957
transform -1 0 29164 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1382_
timestamp 1688980957
transform 1 0 29900 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1383_
timestamp 1688980957
transform 1 0 29440 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1384_
timestamp 1688980957
transform 1 0 31280 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1385_
timestamp 1688980957
transform 1 0 33948 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1386_
timestamp 1688980957
transform 1 0 35236 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1387_
timestamp 1688980957
transform 1 0 32200 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1388_
timestamp 1688980957
transform -1 0 35144 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1389_
timestamp 1688980957
transform 1 0 35328 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1390_
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1688980957
transform 1 0 27968 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1688980957
transform -1 0 31464 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1688980957
transform -1 0 33580 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23092 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 1688980957
transform -1 0 15824 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform 1 0 13984 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform 1 0 20608 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform -1 0 13432 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform -1 0 13432 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform -1 0 19320 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform -1 0 27876 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 33580 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform -1 0 26864 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform -1 0 27968 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform 1 0 33304 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 32752 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_7 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13248 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_8
timestamp 1688980957
transform 1 0 68264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_9
timestamp 1688980957
transform -1 0 26772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_10
timestamp 1688980957
transform 1 0 68264 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_11
timestamp 1688980957
transform -1 0 30636 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_12
timestamp 1688980957
transform -1 0 39652 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_13
timestamp 1688980957
transform 1 0 1380 0 -1 65280
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_265 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_273
timestamp 1688980957
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_461 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_471
timestamp 1688980957
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_475
timestamp 1688980957
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_477
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_489
timestamp 1688980957
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 1688980957
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_505
timestamp 1688980957
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_517
timestamp 1688980957
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 1688980957
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_533
timestamp 1688980957
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_545
timestamp 1688980957
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 1688980957
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_561
timestamp 1688980957
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_573
timestamp 1688980957
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 1688980957
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_589
timestamp 1688980957
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_601
timestamp 1688980957
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 1688980957
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_617
timestamp 1688980957
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_629
timestamp 1688980957
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_641
timestamp 1688980957
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_645
timestamp 1688980957
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_657
timestamp 1688980957
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_669
timestamp 1688980957
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_673
timestamp 1688980957
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_685
timestamp 1688980957
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_697
timestamp 1688980957
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_701
timestamp 1688980957
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_713
timestamp 1688980957
transform 1 0 66700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_721
timestamp 1688980957
transform 1 0 67436 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_729
timestamp 1688980957
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_455
timestamp 1688980957
transform 1 0 42964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_459
timestamp 1688980957
transform 1 0 43332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_471
timestamp 1688980957
transform 1 0 44436 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_483
timestamp 1688980957
transform 1 0 45540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_495
timestamp 1688980957
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 1688980957
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_505
timestamp 1688980957
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_517
timestamp 1688980957
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_529
timestamp 1688980957
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_541
timestamp 1688980957
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_553
timestamp 1688980957
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 1688980957
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_561
timestamp 1688980957
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_573
timestamp 1688980957
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_585
timestamp 1688980957
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_597
timestamp 1688980957
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_609
timestamp 1688980957
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_615
timestamp 1688980957
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_617
timestamp 1688980957
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_629
timestamp 1688980957
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_641
timestamp 1688980957
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_653
timestamp 1688980957
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_665
timestamp 1688980957
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_671
timestamp 1688980957
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_673
timestamp 1688980957
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_685
timestamp 1688980957
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_697
timestamp 1688980957
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_709
timestamp 1688980957
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_721
timestamp 1688980957
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_727
timestamp 1688980957
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_729
timestamp 1688980957
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 1688980957
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 1688980957
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 1688980957
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 1688980957
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 1688980957
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1688980957
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1688980957
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 1688980957
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_569
timestamp 1688980957
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_581
timestamp 1688980957
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 1688980957
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_589
timestamp 1688980957
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_601
timestamp 1688980957
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_613
timestamp 1688980957
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_625
timestamp 1688980957
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_637
timestamp 1688980957
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_643
timestamp 1688980957
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_645
timestamp 1688980957
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_657
timestamp 1688980957
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_669
timestamp 1688980957
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_681
timestamp 1688980957
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_693
timestamp 1688980957
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_699
timestamp 1688980957
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_701
timestamp 1688980957
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_713
timestamp 1688980957
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_725
timestamp 1688980957
transform 1 0 67804 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 1688980957
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 1688980957
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 1688980957
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_505
timestamp 1688980957
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_517
timestamp 1688980957
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 1688980957
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 1688980957
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 1688980957
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 1688980957
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 1688980957
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 1688980957
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 1688980957
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_597
timestamp 1688980957
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_609
timestamp 1688980957
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1688980957
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_617
timestamp 1688980957
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_629
timestamp 1688980957
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_641
timestamp 1688980957
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_653
timestamp 1688980957
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_665
timestamp 1688980957
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_671
timestamp 1688980957
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_673
timestamp 1688980957
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_685
timestamp 1688980957
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_697
timestamp 1688980957
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_709
timestamp 1688980957
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_721
timestamp 1688980957
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_727
timestamp 1688980957
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_729
timestamp 1688980957
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 1688980957
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_501
timestamp 1688980957
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_513
timestamp 1688980957
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_525
timestamp 1688980957
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 1688980957
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 1688980957
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 1688980957
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 1688980957
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 1688980957
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 1688980957
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 1688980957
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1688980957
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1688980957
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1688980957
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_625
timestamp 1688980957
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_637
timestamp 1688980957
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_643
timestamp 1688980957
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_645
timestamp 1688980957
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_657
timestamp 1688980957
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_669
timestamp 1688980957
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_681
timestamp 1688980957
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_693
timestamp 1688980957
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_699
timestamp 1688980957
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_701
timestamp 1688980957
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_713
timestamp 1688980957
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_725
timestamp 1688980957
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 1688980957
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 1688980957
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 1688980957
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 1688980957
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_517
timestamp 1688980957
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_529
timestamp 1688980957
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_541
timestamp 1688980957
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 1688980957
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 1688980957
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 1688980957
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 1688980957
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 1688980957
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 1688980957
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 1688980957
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 1688980957
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_617
timestamp 1688980957
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_629
timestamp 1688980957
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_641
timestamp 1688980957
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_653
timestamp 1688980957
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_665
timestamp 1688980957
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_671
timestamp 1688980957
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_673
timestamp 1688980957
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_685
timestamp 1688980957
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_697
timestamp 1688980957
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_709
timestamp 1688980957
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_721
timestamp 1688980957
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_727
timestamp 1688980957
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_729
timestamp 1688980957
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_489
timestamp 1688980957
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_501
timestamp 1688980957
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_513
timestamp 1688980957
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_525
timestamp 1688980957
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 1688980957
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1688980957
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 1688980957
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 1688980957
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 1688980957
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 1688980957
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 1688980957
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1688980957
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1688980957
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1688980957
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_625
timestamp 1688980957
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_637
timestamp 1688980957
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_643
timestamp 1688980957
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_645
timestamp 1688980957
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_657
timestamp 1688980957
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_669
timestamp 1688980957
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_681
timestamp 1688980957
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_693
timestamp 1688980957
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_699
timestamp 1688980957
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_701
timestamp 1688980957
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_713
timestamp 1688980957
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_725
timestamp 1688980957
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_246
timestamp 1688980957
transform 1 0 23736 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_258
timestamp 1688980957
transform 1 0 24840 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_270
timestamp 1688980957
transform 1 0 25944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_274
timestamp 1688980957
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_299
timestamp 1688980957
transform 1 0 28612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_311
timestamp 1688980957
transform 1 0 29716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_323
timestamp 1688980957
transform 1 0 30820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_485
timestamp 1688980957
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_497
timestamp 1688980957
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_503
timestamp 1688980957
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_505
timestamp 1688980957
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_517
timestamp 1688980957
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_529
timestamp 1688980957
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_541
timestamp 1688980957
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_553
timestamp 1688980957
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 1688980957
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_561
timestamp 1688980957
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_573
timestamp 1688980957
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_585
timestamp 1688980957
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_597
timestamp 1688980957
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 1688980957
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 1688980957
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_617
timestamp 1688980957
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_629
timestamp 1688980957
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_641
timestamp 1688980957
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_653
timestamp 1688980957
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_665
timestamp 1688980957
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_671
timestamp 1688980957
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_673
timestamp 1688980957
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_685
timestamp 1688980957
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_697
timestamp 1688980957
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_709
timestamp 1688980957
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_721
timestamp 1688980957
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_727
timestamp 1688980957
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_729
timestamp 1688980957
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_185 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_190
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_226
timestamp 1688980957
transform 1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_259
timestamp 1688980957
transform 1 0 24932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_280
timestamp 1688980957
transform 1 0 26864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_306
timestamp 1688980957
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_312
timestamp 1688980957
transform 1 0 29808 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_324
timestamp 1688980957
transform 1 0 30912 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_336
timestamp 1688980957
transform 1 0 32016 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_348
timestamp 1688980957
transform 1 0 33120 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_360
timestamp 1688980957
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_489
timestamp 1688980957
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_501
timestamp 1688980957
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_513
timestamp 1688980957
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_525
timestamp 1688980957
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 1688980957
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_533
timestamp 1688980957
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_545
timestamp 1688980957
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_557
timestamp 1688980957
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 1688980957
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 1688980957
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 1688980957
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 1688980957
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 1688980957
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 1688980957
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_625
timestamp 1688980957
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_637
timestamp 1688980957
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_643
timestamp 1688980957
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_645
timestamp 1688980957
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_657
timestamp 1688980957
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_669
timestamp 1688980957
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_681
timestamp 1688980957
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_693
timestamp 1688980957
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_699
timestamp 1688980957
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_701
timestamp 1688980957
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_713
timestamp 1688980957
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_725
timestamp 1688980957
transform 1 0 67804 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1688980957
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_172
timestamp 1688980957
transform 1 0 16928 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_196
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_201
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_246
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_271
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_295
timestamp 1688980957
transform 1 0 28244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_307
timestamp 1688980957
transform 1 0 29348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_319
timestamp 1688980957
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_331
timestamp 1688980957
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 1688980957
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_485
timestamp 1688980957
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_497
timestamp 1688980957
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 1688980957
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 1688980957
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_517
timestamp 1688980957
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_529
timestamp 1688980957
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_541
timestamp 1688980957
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_553
timestamp 1688980957
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_559
timestamp 1688980957
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_561
timestamp 1688980957
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 1688980957
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 1688980957
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 1688980957
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 1688980957
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 1688980957
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_617
timestamp 1688980957
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_629
timestamp 1688980957
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_641
timestamp 1688980957
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_653
timestamp 1688980957
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_665
timestamp 1688980957
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_671
timestamp 1688980957
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_673
timestamp 1688980957
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_685
timestamp 1688980957
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_697
timestamp 1688980957
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_709
timestamp 1688980957
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_721
timestamp 1688980957
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_727
timestamp 1688980957
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_729
timestamp 1688980957
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_181
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_206
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_214
timestamp 1688980957
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_220
timestamp 1688980957
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_232
timestamp 1688980957
transform 1 0 22448 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_238
timestamp 1688980957
transform 1 0 23000 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_272
timestamp 1688980957
transform 1 0 26128 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_280
timestamp 1688980957
transform 1 0 26864 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_285
timestamp 1688980957
transform 1 0 27324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_297
timestamp 1688980957
transform 1 0 28428 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_306
timestamp 1688980957
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_318
timestamp 1688980957
transform 1 0 30360 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_330
timestamp 1688980957
transform 1 0 31464 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_342
timestamp 1688980957
transform 1 0 32568 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_354
timestamp 1688980957
transform 1 0 33672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_362
timestamp 1688980957
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 1688980957
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_489
timestamp 1688980957
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_501
timestamp 1688980957
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_513
timestamp 1688980957
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_525
timestamp 1688980957
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_531
timestamp 1688980957
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 1688980957
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 1688980957
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 1688980957
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 1688980957
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 1688980957
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 1688980957
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 1688980957
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 1688980957
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_613
timestamp 1688980957
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_625
timestamp 1688980957
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_637
timestamp 1688980957
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_643
timestamp 1688980957
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_645
timestamp 1688980957
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_657
timestamp 1688980957
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_669
timestamp 1688980957
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_681
timestamp 1688980957
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_693
timestamp 1688980957
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_699
timestamp 1688980957
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_701
timestamp 1688980957
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_713
timestamp 1688980957
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_725
timestamp 1688980957
transform 1 0 67804 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_178
timestamp 1688980957
transform 1 0 17480 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_186
timestamp 1688980957
transform 1 0 18216 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_204
timestamp 1688980957
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_218
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_236
timestamp 1688980957
transform 1 0 22816 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_245
timestamp 1688980957
transform 1 0 23644 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_275
timestamp 1688980957
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_287
timestamp 1688980957
transform 1 0 27508 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_291
timestamp 1688980957
transform 1 0 27876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_325
timestamp 1688980957
transform 1 0 31004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_333
timestamp 1688980957
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_473
timestamp 1688980957
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_485
timestamp 1688980957
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_497
timestamp 1688980957
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 1688980957
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_505
timestamp 1688980957
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 1688980957
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_529
timestamp 1688980957
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_541
timestamp 1688980957
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_553
timestamp 1688980957
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 1688980957
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 1688980957
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 1688980957
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 1688980957
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 1688980957
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 1688980957
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1688980957
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_617
timestamp 1688980957
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_629
timestamp 1688980957
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_641
timestamp 1688980957
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_653
timestamp 1688980957
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_665
timestamp 1688980957
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_671
timestamp 1688980957
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_673
timestamp 1688980957
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_685
timestamp 1688980957
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_697
timestamp 1688980957
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_709
timestamp 1688980957
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_721
timestamp 1688980957
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_727
timestamp 1688980957
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_729
timestamp 1688980957
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_159
timestamp 1688980957
transform 1 0 15732 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_163
timestamp 1688980957
transform 1 0 16100 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_171
timestamp 1688980957
transform 1 0 16836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_178
timestamp 1688980957
transform 1 0 17480 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_183
timestamp 1688980957
transform 1 0 17940 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_257
timestamp 1688980957
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_271
timestamp 1688980957
transform 1 0 26036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_283
timestamp 1688980957
transform 1 0 27140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_306
timestamp 1688980957
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_358
timestamp 1688980957
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 1688980957
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_489
timestamp 1688980957
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_501
timestamp 1688980957
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_513
timestamp 1688980957
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_525
timestamp 1688980957
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 1688980957
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 1688980957
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 1688980957
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 1688980957
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 1688980957
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 1688980957
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 1688980957
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 1688980957
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 1688980957
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 1688980957
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_625
timestamp 1688980957
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_637
timestamp 1688980957
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_643
timestamp 1688980957
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_645
timestamp 1688980957
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_657
timestamp 1688980957
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_669
timestamp 1688980957
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_681
timestamp 1688980957
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_693
timestamp 1688980957
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_699
timestamp 1688980957
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_701
timestamp 1688980957
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_713
timestamp 1688980957
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_725
timestamp 1688980957
transform 1 0 67804 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_184
timestamp 1688980957
transform 1 0 18032 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_196
timestamp 1688980957
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_208
timestamp 1688980957
transform 1 0 20240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_214
timestamp 1688980957
transform 1 0 20792 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_242
timestamp 1688980957
transform 1 0 23368 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_255
timestamp 1688980957
transform 1 0 24564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_266
timestamp 1688980957
transform 1 0 25576 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_312
timestamp 1688980957
transform 1 0 29808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_346
timestamp 1688980957
transform 1 0 32936 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_380
timestamp 1688980957
transform 1 0 36064 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1688980957
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 1688980957
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 1688980957
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 1688980957
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_473
timestamp 1688980957
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_485
timestamp 1688980957
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_497
timestamp 1688980957
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 1688980957
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 1688980957
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_517
timestamp 1688980957
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_529
timestamp 1688980957
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_541
timestamp 1688980957
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 1688980957
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 1688980957
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_561
timestamp 1688980957
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_573
timestamp 1688980957
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_585
timestamp 1688980957
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_597
timestamp 1688980957
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_609
timestamp 1688980957
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 1688980957
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_617
timestamp 1688980957
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_629
timestamp 1688980957
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_641
timestamp 1688980957
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_653
timestamp 1688980957
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_665
timestamp 1688980957
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_671
timestamp 1688980957
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_673
timestamp 1688980957
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_685
timestamp 1688980957
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_697
timestamp 1688980957
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_709
timestamp 1688980957
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_721
timestamp 1688980957
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_727
timestamp 1688980957
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_729
timestamp 1688980957
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_168
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_203
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_207
timestamp 1688980957
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_214
timestamp 1688980957
transform 1 0 20792 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_226
timestamp 1688980957
transform 1 0 21896 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_238
timestamp 1688980957
transform 1 0 23000 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_247
timestamp 1688980957
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_279
timestamp 1688980957
transform 1 0 26772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_291
timestamp 1688980957
transform 1 0 27876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_303
timestamp 1688980957
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_312
timestamp 1688980957
transform 1 0 29808 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_349
timestamp 1688980957
transform 1 0 33212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_358
timestamp 1688980957
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_376
timestamp 1688980957
transform 1 0 35696 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_388
timestamp 1688980957
transform 1 0 36800 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_400
timestamp 1688980957
transform 1 0 37904 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_412
timestamp 1688980957
transform 1 0 39008 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_433
timestamp 1688980957
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 1688980957
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_457
timestamp 1688980957
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_469
timestamp 1688980957
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 1688980957
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_477
timestamp 1688980957
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_489
timestamp 1688980957
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_501
timestamp 1688980957
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_513
timestamp 1688980957
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_525
timestamp 1688980957
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 1688980957
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_533
timestamp 1688980957
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_545
timestamp 1688980957
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_557
timestamp 1688980957
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_569
timestamp 1688980957
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_581
timestamp 1688980957
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_587
timestamp 1688980957
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_589
timestamp 1688980957
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_601
timestamp 1688980957
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_613
timestamp 1688980957
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_625
timestamp 1688980957
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_637
timestamp 1688980957
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_643
timestamp 1688980957
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_645
timestamp 1688980957
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_657
timestamp 1688980957
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_669
timestamp 1688980957
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_681
timestamp 1688980957
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_693
timestamp 1688980957
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_699
timestamp 1688980957
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_701
timestamp 1688980957
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_713
timestamp 1688980957
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_725
timestamp 1688980957
transform 1 0 67804 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_729
timestamp 1688980957
transform 1 0 68172 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_198
timestamp 1688980957
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_207
timestamp 1688980957
transform 1 0 20148 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_219
timestamp 1688980957
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_233
timestamp 1688980957
transform 1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_256
timestamp 1688980957
transform 1 0 24656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_284
timestamp 1688980957
transform 1 0 27232 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_288
timestamp 1688980957
transform 1 0 27600 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_298
timestamp 1688980957
transform 1 0 28520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_306
timestamp 1688980957
transform 1 0 29256 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_331
timestamp 1688980957
transform 1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_345
timestamp 1688980957
transform 1 0 32844 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_352
timestamp 1688980957
transform 1 0 33488 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_364
timestamp 1688980957
transform 1 0 34592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_371
timestamp 1688980957
transform 1 0 35236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1688980957
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 1688980957
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 1688980957
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_429
timestamp 1688980957
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_441
timestamp 1688980957
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_447
timestamp 1688980957
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_461
timestamp 1688980957
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_473
timestamp 1688980957
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_485
timestamp 1688980957
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_497
timestamp 1688980957
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_503
timestamp 1688980957
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_505
timestamp 1688980957
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_517
timestamp 1688980957
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_529
timestamp 1688980957
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_541
timestamp 1688980957
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_553
timestamp 1688980957
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_559
timestamp 1688980957
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_561
timestamp 1688980957
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_573
timestamp 1688980957
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_585
timestamp 1688980957
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_597
timestamp 1688980957
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_609
timestamp 1688980957
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_615
timestamp 1688980957
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_617
timestamp 1688980957
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_629
timestamp 1688980957
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_641
timestamp 1688980957
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_653
timestamp 1688980957
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_665
timestamp 1688980957
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_671
timestamp 1688980957
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_673
timestamp 1688980957
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_685
timestamp 1688980957
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_697
timestamp 1688980957
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_709
timestamp 1688980957
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_721
timestamp 1688980957
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_727
timestamp 1688980957
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_729
timestamp 1688980957
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_123
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_135
timestamp 1688980957
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_178
timestamp 1688980957
transform 1 0 17480 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_192
timestamp 1688980957
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_211
timestamp 1688980957
transform 1 0 20516 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_218
timestamp 1688980957
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_226
timestamp 1688980957
transform 1 0 21896 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_238
timestamp 1688980957
transform 1 0 23000 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_246
timestamp 1688980957
transform 1 0 23736 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_268
timestamp 1688980957
transform 1 0 25760 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_272
timestamp 1688980957
transform 1 0 26128 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_313
timestamp 1688980957
transform 1 0 29900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_317
timestamp 1688980957
transform 1 0 30268 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_325
timestamp 1688980957
transform 1 0 31004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_335
timestamp 1688980957
transform 1 0 31924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_353
timestamp 1688980957
transform 1 0 33580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_391
timestamp 1688980957
transform 1 0 37076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_403
timestamp 1688980957
transform 1 0 38180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_415
timestamp 1688980957
transform 1 0 39284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 1688980957
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 1688980957
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_445
timestamp 1688980957
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_457
timestamp 1688980957
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_469
timestamp 1688980957
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_475
timestamp 1688980957
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_477
timestamp 1688980957
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_489
timestamp 1688980957
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_501
timestamp 1688980957
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_513
timestamp 1688980957
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_525
timestamp 1688980957
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_531
timestamp 1688980957
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_533
timestamp 1688980957
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_545
timestamp 1688980957
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_557
timestamp 1688980957
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_569
timestamp 1688980957
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_581
timestamp 1688980957
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_587
timestamp 1688980957
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_589
timestamp 1688980957
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_601
timestamp 1688980957
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_613
timestamp 1688980957
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_625
timestamp 1688980957
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_637
timestamp 1688980957
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_643
timestamp 1688980957
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_645
timestamp 1688980957
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_657
timestamp 1688980957
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_669
timestamp 1688980957
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_681
timestamp 1688980957
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_693
timestamp 1688980957
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_699
timestamp 1688980957
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_701
timestamp 1688980957
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_713
timestamp 1688980957
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_725
timestamp 1688980957
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_116
timestamp 1688980957
transform 1 0 11776 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_128
timestamp 1688980957
transform 1 0 12880 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_132
timestamp 1688980957
transform 1 0 13248 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_144
timestamp 1688980957
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_148
timestamp 1688980957
transform 1 0 14720 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_160
timestamp 1688980957
transform 1 0 15824 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_164
timestamp 1688980957
transform 1 0 16192 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_186
timestamp 1688980957
transform 1 0 18216 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_194
timestamp 1688980957
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_219
timestamp 1688980957
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_230
timestamp 1688980957
transform 1 0 22264 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_239
timestamp 1688980957
transform 1 0 23092 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_269
timestamp 1688980957
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_324
timestamp 1688980957
transform 1 0 30912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_333
timestamp 1688980957
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_358
timestamp 1688980957
transform 1 0 34040 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_364
timestamp 1688980957
transform 1 0 34592 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 1688980957
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 1688980957
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_429
timestamp 1688980957
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_441
timestamp 1688980957
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 1688980957
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 1688980957
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_461
timestamp 1688980957
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_473
timestamp 1688980957
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_485
timestamp 1688980957
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_497
timestamp 1688980957
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_503
timestamp 1688980957
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_505
timestamp 1688980957
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_517
timestamp 1688980957
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_529
timestamp 1688980957
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_541
timestamp 1688980957
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_553
timestamp 1688980957
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_559
timestamp 1688980957
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_561
timestamp 1688980957
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_573
timestamp 1688980957
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_585
timestamp 1688980957
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_597
timestamp 1688980957
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_609
timestamp 1688980957
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 1688980957
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_617
timestamp 1688980957
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_629
timestamp 1688980957
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_641
timestamp 1688980957
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_653
timestamp 1688980957
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_665
timestamp 1688980957
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_671
timestamp 1688980957
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_673
timestamp 1688980957
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_685
timestamp 1688980957
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_697
timestamp 1688980957
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_709
timestamp 1688980957
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_721
timestamp 1688980957
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_727
timestamp 1688980957
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_729
timestamp 1688980957
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_92
timestamp 1688980957
transform 1 0 9568 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_107
timestamp 1688980957
transform 1 0 10948 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_115
timestamp 1688980957
transform 1 0 11684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_173
timestamp 1688980957
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_181
timestamp 1688980957
transform 1 0 17756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1688980957
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_206
timestamp 1688980957
transform 1 0 20056 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_228
timestamp 1688980957
transform 1 0 22080 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_239
timestamp 1688980957
transform 1 0 23092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_281
timestamp 1688980957
transform 1 0 26956 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_300
timestamp 1688980957
transform 1 0 28704 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_335
timestamp 1688980957
transform 1 0 31924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_344
timestamp 1688980957
transform 1 0 32752 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_352
timestamp 1688980957
transform 1 0 33488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_361
timestamp 1688980957
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_368
timestamp 1688980957
transform 1 0 34960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_379
timestamp 1688980957
transform 1 0 35972 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_385
timestamp 1688980957
transform 1 0 36524 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_397
timestamp 1688980957
transform 1 0 37628 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_409
timestamp 1688980957
transform 1 0 38732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_417
timestamp 1688980957
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 1688980957
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 1688980957
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_457
timestamp 1688980957
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_469
timestamp 1688980957
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 1688980957
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_477
timestamp 1688980957
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_489
timestamp 1688980957
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_501
timestamp 1688980957
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_513
timestamp 1688980957
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_525
timestamp 1688980957
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_531
timestamp 1688980957
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_533
timestamp 1688980957
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_545
timestamp 1688980957
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_557
timestamp 1688980957
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_569
timestamp 1688980957
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_581
timestamp 1688980957
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_587
timestamp 1688980957
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_589
timestamp 1688980957
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_601
timestamp 1688980957
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_613
timestamp 1688980957
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_625
timestamp 1688980957
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_637
timestamp 1688980957
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_643
timestamp 1688980957
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_645
timestamp 1688980957
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_657
timestamp 1688980957
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_669
timestamp 1688980957
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_681
timestamp 1688980957
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_693
timestamp 1688980957
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_699
timestamp 1688980957
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_701
timestamp 1688980957
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_713
timestamp 1688980957
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_725
timestamp 1688980957
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_77
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_99
timestamp 1688980957
transform 1 0 10212 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_107
timestamp 1688980957
transform 1 0 10948 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_130
timestamp 1688980957
transform 1 0 13064 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_151
timestamp 1688980957
transform 1 0 14996 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_163
timestamp 1688980957
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_184
timestamp 1688980957
transform 1 0 18032 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_248
timestamp 1688980957
transform 1 0 23920 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_254
timestamp 1688980957
transform 1 0 24472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_267
timestamp 1688980957
transform 1 0 25668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_322
timestamp 1688980957
transform 1 0 30728 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_333
timestamp 1688980957
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_343
timestamp 1688980957
transform 1 0 32660 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_347
timestamp 1688980957
transform 1 0 33028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_355
timestamp 1688980957
transform 1 0 33764 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_401
timestamp 1688980957
transform 1 0 37996 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_413
timestamp 1688980957
transform 1 0 39100 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_425
timestamp 1688980957
transform 1 0 40204 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_437
timestamp 1688980957
transform 1 0 41308 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_445
timestamp 1688980957
transform 1 0 42044 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_449
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_461
timestamp 1688980957
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_473
timestamp 1688980957
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_485
timestamp 1688980957
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_497
timestamp 1688980957
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_503
timestamp 1688980957
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_505
timestamp 1688980957
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_517
timestamp 1688980957
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_529
timestamp 1688980957
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_541
timestamp 1688980957
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_553
timestamp 1688980957
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_559
timestamp 1688980957
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_561
timestamp 1688980957
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_573
timestamp 1688980957
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_585
timestamp 1688980957
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_597
timestamp 1688980957
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_609
timestamp 1688980957
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_615
timestamp 1688980957
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_617
timestamp 1688980957
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_629
timestamp 1688980957
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_641
timestamp 1688980957
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_653
timestamp 1688980957
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_665
timestamp 1688980957
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_671
timestamp 1688980957
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_673
timestamp 1688980957
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_685
timestamp 1688980957
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_697
timestamp 1688980957
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_709
timestamp 1688980957
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_721
timestamp 1688980957
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_727
timestamp 1688980957
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_729
timestamp 1688980957
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_89
timestamp 1688980957
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_115
timestamp 1688980957
transform 1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_122
timestamp 1688980957
transform 1 0 12328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_130
timestamp 1688980957
transform 1 0 13064 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_136
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_149
timestamp 1688980957
transform 1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_187
timestamp 1688980957
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_205
timestamp 1688980957
transform 1 0 19964 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_227
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_231
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_241
timestamp 1688980957
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1688980957
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_291
timestamp 1688980957
transform 1 0 27876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_302
timestamp 1688980957
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_325
timestamp 1688980957
transform 1 0 31004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_337
timestamp 1688980957
transform 1 0 32108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_358
timestamp 1688980957
transform 1 0 34040 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1688980957
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_401
timestamp 1688980957
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_413
timestamp 1688980957
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_419
timestamp 1688980957
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_421
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_433
timestamp 1688980957
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_445
timestamp 1688980957
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_457
timestamp 1688980957
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_469
timestamp 1688980957
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_475
timestamp 1688980957
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_477
timestamp 1688980957
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_489
timestamp 1688980957
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_501
timestamp 1688980957
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_513
timestamp 1688980957
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_525
timestamp 1688980957
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_531
timestamp 1688980957
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_533
timestamp 1688980957
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_545
timestamp 1688980957
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_557
timestamp 1688980957
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_569
timestamp 1688980957
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_581
timestamp 1688980957
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_587
timestamp 1688980957
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_589
timestamp 1688980957
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_601
timestamp 1688980957
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_613
timestamp 1688980957
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_625
timestamp 1688980957
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_637
timestamp 1688980957
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_643
timestamp 1688980957
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_645
timestamp 1688980957
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_657
timestamp 1688980957
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_669
timestamp 1688980957
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_681
timestamp 1688980957
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_693
timestamp 1688980957
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_699
timestamp 1688980957
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_701
timestamp 1688980957
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_713
timestamp 1688980957
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_725
timestamp 1688980957
transform 1 0 67804 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_91
timestamp 1688980957
transform 1 0 9476 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_100
timestamp 1688980957
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1688980957
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_145
timestamp 1688980957
transform 1 0 14444 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_154
timestamp 1688980957
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1688980957
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_176
timestamp 1688980957
transform 1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_191
timestamp 1688980957
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_209
timestamp 1688980957
transform 1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_214
timestamp 1688980957
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_234
timestamp 1688980957
transform 1 0 22632 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_269
timestamp 1688980957
transform 1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_275
timestamp 1688980957
transform 1 0 26404 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_297
timestamp 1688980957
transform 1 0 28428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_341
timestamp 1688980957
transform 1 0 32476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_345
timestamp 1688980957
transform 1 0 32844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_370
timestamp 1688980957
transform 1 0 35144 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_382
timestamp 1688980957
transform 1 0 36248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_390
timestamp 1688980957
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 1688980957
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_417
timestamp 1688980957
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_429
timestamp 1688980957
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_441
timestamp 1688980957
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_447
timestamp 1688980957
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_461
timestamp 1688980957
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_473
timestamp 1688980957
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_485
timestamp 1688980957
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_497
timestamp 1688980957
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_503
timestamp 1688980957
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_505
timestamp 1688980957
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_517
timestamp 1688980957
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_529
timestamp 1688980957
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_541
timestamp 1688980957
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_553
timestamp 1688980957
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_559
timestamp 1688980957
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_561
timestamp 1688980957
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_573
timestamp 1688980957
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_585
timestamp 1688980957
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_597
timestamp 1688980957
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_609
timestamp 1688980957
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_615
timestamp 1688980957
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_617
timestamp 1688980957
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_629
timestamp 1688980957
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_641
timestamp 1688980957
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_653
timestamp 1688980957
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_665
timestamp 1688980957
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_671
timestamp 1688980957
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_673
timestamp 1688980957
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_685
timestamp 1688980957
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_697
timestamp 1688980957
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_709
timestamp 1688980957
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_721
timestamp 1688980957
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_727
timestamp 1688980957
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_729
timestamp 1688980957
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_105
timestamp 1688980957
transform 1 0 10764 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_114
timestamp 1688980957
transform 1 0 11592 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_118
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_144
timestamp 1688980957
transform 1 0 14352 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_162
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_168
timestamp 1688980957
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_176
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_187
timestamp 1688980957
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_216
timestamp 1688980957
transform 1 0 20976 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_234
timestamp 1688980957
transform 1 0 22632 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_242
timestamp 1688980957
transform 1 0 23368 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_279
timestamp 1688980957
transform 1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_295
timestamp 1688980957
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_315
timestamp 1688980957
transform 1 0 30084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_327
timestamp 1688980957
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_335
timestamp 1688980957
transform 1 0 31924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_343
timestamp 1688980957
transform 1 0 32660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_356
timestamp 1688980957
transform 1 0 33856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_360
timestamp 1688980957
transform 1 0 34224 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1688980957
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_401
timestamp 1688980957
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 1688980957
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1688980957
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_433
timestamp 1688980957
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_445
timestamp 1688980957
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_457
timestamp 1688980957
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_469
timestamp 1688980957
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_475
timestamp 1688980957
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_477
timestamp 1688980957
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_489
timestamp 1688980957
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_501
timestamp 1688980957
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_513
timestamp 1688980957
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_525
timestamp 1688980957
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_531
timestamp 1688980957
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_533
timestamp 1688980957
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_545
timestamp 1688980957
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_557
timestamp 1688980957
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_569
timestamp 1688980957
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_581
timestamp 1688980957
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_587
timestamp 1688980957
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_589
timestamp 1688980957
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_601
timestamp 1688980957
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_613
timestamp 1688980957
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_625
timestamp 1688980957
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_637
timestamp 1688980957
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_643
timestamp 1688980957
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_645
timestamp 1688980957
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_657
timestamp 1688980957
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_669
timestamp 1688980957
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_681
timestamp 1688980957
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_693
timestamp 1688980957
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_699
timestamp 1688980957
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_701
timestamp 1688980957
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_713
timestamp 1688980957
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_725
timestamp 1688980957
transform 1 0 67804 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_73
timestamp 1688980957
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_77
timestamp 1688980957
transform 1 0 8188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_83
timestamp 1688980957
transform 1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_91
timestamp 1688980957
transform 1 0 9476 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_98
timestamp 1688980957
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1688980957
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_123
timestamp 1688980957
transform 1 0 12420 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_131
timestamp 1688980957
transform 1 0 13156 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_139
timestamp 1688980957
transform 1 0 13892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_269
timestamp 1688980957
transform 1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_291
timestamp 1688980957
transform 1 0 27876 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_309
timestamp 1688980957
transform 1 0 29532 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_364
timestamp 1688980957
transform 1 0 34592 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_379
timestamp 1688980957
transform 1 0 35972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1688980957
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_405
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_417
timestamp 1688980957
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_429
timestamp 1688980957
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_441
timestamp 1688980957
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 1688980957
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_449
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_461
timestamp 1688980957
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_473
timestamp 1688980957
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_485
timestamp 1688980957
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_497
timestamp 1688980957
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_503
timestamp 1688980957
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_505
timestamp 1688980957
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_517
timestamp 1688980957
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_529
timestamp 1688980957
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_541
timestamp 1688980957
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_553
timestamp 1688980957
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_559
timestamp 1688980957
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_561
timestamp 1688980957
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_573
timestamp 1688980957
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_585
timestamp 1688980957
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_597
timestamp 1688980957
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_609
timestamp 1688980957
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_615
timestamp 1688980957
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_617
timestamp 1688980957
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_629
timestamp 1688980957
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_641
timestamp 1688980957
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_653
timestamp 1688980957
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_665
timestamp 1688980957
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_671
timestamp 1688980957
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_673
timestamp 1688980957
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_685
timestamp 1688980957
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_697
timestamp 1688980957
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_709
timestamp 1688980957
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_721
timestamp 1688980957
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_727
timestamp 1688980957
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_729
timestamp 1688980957
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_61
timestamp 1688980957
transform 1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_95
timestamp 1688980957
transform 1 0 9844 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_99
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_105
timestamp 1688980957
transform 1 0 10764 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_112
timestamp 1688980957
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_119
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_131
timestamp 1688980957
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_157
timestamp 1688980957
transform 1 0 15548 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_161
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_236
timestamp 1688980957
transform 1 0 22816 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_270
timestamp 1688980957
transform 1 0 25944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_289
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_298
timestamp 1688980957
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_316
timestamp 1688980957
transform 1 0 30176 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_331
timestamp 1688980957
transform 1 0 31556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_395
timestamp 1688980957
transform 1 0 37444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_407
timestamp 1688980957
transform 1 0 38548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1688980957
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_433
timestamp 1688980957
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_445
timestamp 1688980957
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_457
timestamp 1688980957
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_469
timestamp 1688980957
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_475
timestamp 1688980957
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_477
timestamp 1688980957
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_489
timestamp 1688980957
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_501
timestamp 1688980957
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_513
timestamp 1688980957
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_525
timestamp 1688980957
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_531
timestamp 1688980957
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_533
timestamp 1688980957
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_545
timestamp 1688980957
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_557
timestamp 1688980957
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_569
timestamp 1688980957
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_581
timestamp 1688980957
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_587
timestamp 1688980957
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_589
timestamp 1688980957
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_601
timestamp 1688980957
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_613
timestamp 1688980957
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_625
timestamp 1688980957
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_637
timestamp 1688980957
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_643
timestamp 1688980957
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_645
timestamp 1688980957
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_657
timestamp 1688980957
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_669
timestamp 1688980957
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_681
timestamp 1688980957
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_693
timestamp 1688980957
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_699
timestamp 1688980957
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_701
timestamp 1688980957
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_713
timestamp 1688980957
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_725
timestamp 1688980957
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_98
timestamp 1688980957
transform 1 0 10120 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_140
timestamp 1688980957
transform 1 0 13984 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_148
timestamp 1688980957
transform 1 0 14720 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_185
timestamp 1688980957
transform 1 0 18124 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_241
timestamp 1688980957
transform 1 0 23276 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_250
timestamp 1688980957
transform 1 0 24104 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_274
timestamp 1688980957
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_300
timestamp 1688980957
transform 1 0 28704 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_308
timestamp 1688980957
transform 1 0 29440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_325
timestamp 1688980957
transform 1 0 31004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_333
timestamp 1688980957
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_375
timestamp 1688980957
transform 1 0 35604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_387
timestamp 1688980957
transform 1 0 36708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1688980957
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1688980957
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1688980957
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_429
timestamp 1688980957
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_441
timestamp 1688980957
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 1688980957
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_449
timestamp 1688980957
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_461
timestamp 1688980957
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_473
timestamp 1688980957
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_485
timestamp 1688980957
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_497
timestamp 1688980957
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_503
timestamp 1688980957
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_505
timestamp 1688980957
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_517
timestamp 1688980957
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_529
timestamp 1688980957
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_541
timestamp 1688980957
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_553
timestamp 1688980957
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_559
timestamp 1688980957
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_561
timestamp 1688980957
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_573
timestamp 1688980957
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_585
timestamp 1688980957
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_597
timestamp 1688980957
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_609
timestamp 1688980957
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_615
timestamp 1688980957
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_617
timestamp 1688980957
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_629
timestamp 1688980957
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_641
timestamp 1688980957
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_653
timestamp 1688980957
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_665
timestamp 1688980957
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_671
timestamp 1688980957
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_673
timestamp 1688980957
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_685
timestamp 1688980957
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_697
timestamp 1688980957
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_709
timestamp 1688980957
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_721
timestamp 1688980957
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_727
timestamp 1688980957
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_729
timestamp 1688980957
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_104
timestamp 1688980957
transform 1 0 10672 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_118
timestamp 1688980957
transform 1 0 11960 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_144
timestamp 1688980957
transform 1 0 14352 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_186
timestamp 1688980957
transform 1 0 18216 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_192
timestamp 1688980957
transform 1 0 18768 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_219
timestamp 1688980957
transform 1 0 21252 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_283
timestamp 1688980957
transform 1 0 27140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_330
timestamp 1688980957
transform 1 0 31464 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_349
timestamp 1688980957
transform 1 0 33212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_361
timestamp 1688980957
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_377
timestamp 1688980957
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_397
timestamp 1688980957
transform 1 0 37628 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_409
timestamp 1688980957
transform 1 0 38732 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_417
timestamp 1688980957
transform 1 0 39468 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_433
timestamp 1688980957
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_445
timestamp 1688980957
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_457
timestamp 1688980957
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_469
timestamp 1688980957
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_475
timestamp 1688980957
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_477
timestamp 1688980957
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_489
timestamp 1688980957
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_501
timestamp 1688980957
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_513
timestamp 1688980957
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_525
timestamp 1688980957
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_531
timestamp 1688980957
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_533
timestamp 1688980957
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_545
timestamp 1688980957
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_557
timestamp 1688980957
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_569
timestamp 1688980957
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_581
timestamp 1688980957
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_587
timestamp 1688980957
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_589
timestamp 1688980957
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_601
timestamp 1688980957
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_613
timestamp 1688980957
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_625
timestamp 1688980957
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_637
timestamp 1688980957
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_643
timestamp 1688980957
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_645
timestamp 1688980957
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_657
timestamp 1688980957
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_669
timestamp 1688980957
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_681
timestamp 1688980957
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_693
timestamp 1688980957
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_699
timestamp 1688980957
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_701
timestamp 1688980957
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_713
timestamp 1688980957
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_725
timestamp 1688980957
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_89
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_107
timestamp 1688980957
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_121
timestamp 1688980957
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_177
timestamp 1688980957
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_203
timestamp 1688980957
transform 1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_221
timestamp 1688980957
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_229
timestamp 1688980957
transform 1 0 22172 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_259
timestamp 1688980957
transform 1 0 24932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_269
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_289
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_299
timestamp 1688980957
transform 1 0 28612 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_307
timestamp 1688980957
transform 1 0 29348 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_314
timestamp 1688980957
transform 1 0 29992 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_326
timestamp 1688980957
transform 1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_334
timestamp 1688980957
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_360
timestamp 1688980957
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_364
timestamp 1688980957
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_373
timestamp 1688980957
transform 1 0 35420 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_389
timestamp 1688980957
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 1688980957
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_417
timestamp 1688980957
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_429
timestamp 1688980957
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_441
timestamp 1688980957
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_447
timestamp 1688980957
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_449
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_461
timestamp 1688980957
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_473
timestamp 1688980957
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_485
timestamp 1688980957
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_497
timestamp 1688980957
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_503
timestamp 1688980957
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_505
timestamp 1688980957
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_517
timestamp 1688980957
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_529
timestamp 1688980957
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_541
timestamp 1688980957
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_553
timestamp 1688980957
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_559
timestamp 1688980957
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_561
timestamp 1688980957
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_573
timestamp 1688980957
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_585
timestamp 1688980957
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_597
timestamp 1688980957
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_609
timestamp 1688980957
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_615
timestamp 1688980957
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_617
timestamp 1688980957
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_629
timestamp 1688980957
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_641
timestamp 1688980957
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_653
timestamp 1688980957
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_665
timestamp 1688980957
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_671
timestamp 1688980957
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_673
timestamp 1688980957
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_685
timestamp 1688980957
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_697
timestamp 1688980957
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_709
timestamp 1688980957
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_721
timestamp 1688980957
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_727
timestamp 1688980957
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_729
timestamp 1688980957
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_88
timestamp 1688980957
transform 1 0 9200 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_100
timestamp 1688980957
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_132
timestamp 1688980957
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_149
timestamp 1688980957
transform 1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_187
timestamp 1688980957
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_206
timestamp 1688980957
transform 1 0 20056 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_212
timestamp 1688980957
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_222
timestamp 1688980957
transform 1 0 21528 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_256
timestamp 1688980957
transform 1 0 24656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_260
timestamp 1688980957
transform 1 0 25024 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_296
timestamp 1688980957
transform 1 0 28336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_324
timestamp 1688980957
transform 1 0 30912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_358
timestamp 1688980957
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_381
timestamp 1688980957
transform 1 0 36156 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_405
timestamp 1688980957
transform 1 0 38364 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_417
timestamp 1688980957
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 1688980957
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_445
timestamp 1688980957
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_457
timestamp 1688980957
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_469
timestamp 1688980957
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_475
timestamp 1688980957
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_477
timestamp 1688980957
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_489
timestamp 1688980957
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_501
timestamp 1688980957
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_513
timestamp 1688980957
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_525
timestamp 1688980957
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_531
timestamp 1688980957
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_533
timestamp 1688980957
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_545
timestamp 1688980957
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_557
timestamp 1688980957
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_569
timestamp 1688980957
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_581
timestamp 1688980957
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_587
timestamp 1688980957
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_589
timestamp 1688980957
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_601
timestamp 1688980957
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_613
timestamp 1688980957
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_625
timestamp 1688980957
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_637
timestamp 1688980957
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_643
timestamp 1688980957
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_645
timestamp 1688980957
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_657
timestamp 1688980957
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_669
timestamp 1688980957
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_681
timestamp 1688980957
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_693
timestamp 1688980957
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_699
timestamp 1688980957
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_701
timestamp 1688980957
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_713
timestamp 1688980957
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_725
timestamp 1688980957
transform 1 0 67804 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_116
timestamp 1688980957
transform 1 0 11776 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_128
timestamp 1688980957
transform 1 0 12880 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_154
timestamp 1688980957
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1688980957
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_177
timestamp 1688980957
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_231
timestamp 1688980957
transform 1 0 22356 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_266
timestamp 1688980957
transform 1 0 25576 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_272
timestamp 1688980957
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_289
timestamp 1688980957
transform 1 0 27692 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_306
timestamp 1688980957
transform 1 0 29256 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_333
timestamp 1688980957
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_374
timestamp 1688980957
transform 1 0 35512 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_382
timestamp 1688980957
transform 1 0 36248 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 1688980957
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_409
timestamp 1688980957
transform 1 0 38732 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_421
timestamp 1688980957
transform 1 0 39836 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_433
timestamp 1688980957
transform 1 0 40940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_445
timestamp 1688980957
transform 1 0 42044 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 1688980957
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_461
timestamp 1688980957
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_473
timestamp 1688980957
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_485
timestamp 1688980957
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_497
timestamp 1688980957
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_503
timestamp 1688980957
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_505
timestamp 1688980957
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_517
timestamp 1688980957
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_529
timestamp 1688980957
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_541
timestamp 1688980957
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_553
timestamp 1688980957
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_559
timestamp 1688980957
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_561
timestamp 1688980957
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_573
timestamp 1688980957
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_585
timestamp 1688980957
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_597
timestamp 1688980957
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_609
timestamp 1688980957
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_615
timestamp 1688980957
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_617
timestamp 1688980957
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_629
timestamp 1688980957
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_641
timestamp 1688980957
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_653
timestamp 1688980957
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_665
timestamp 1688980957
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_671
timestamp 1688980957
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_673
timestamp 1688980957
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_685
timestamp 1688980957
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_697
timestamp 1688980957
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_709
timestamp 1688980957
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_721
timestamp 1688980957
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_727
timestamp 1688980957
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_729
timestamp 1688980957
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_89
timestamp 1688980957
transform 1 0 9292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_104
timestamp 1688980957
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_125
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_149
timestamp 1688980957
transform 1 0 14812 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_159
timestamp 1688980957
transform 1 0 15732 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_186
timestamp 1688980957
transform 1 0 18216 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_216
timestamp 1688980957
transform 1 0 20976 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_222
timestamp 1688980957
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_232
timestamp 1688980957
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_236
timestamp 1688980957
transform 1 0 22816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_285
timestamp 1688980957
transform 1 0 27324 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_293
timestamp 1688980957
transform 1 0 28060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_304
timestamp 1688980957
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_336
timestamp 1688980957
transform 1 0 32016 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_362
timestamp 1688980957
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_369
timestamp 1688980957
transform 1 0 35052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_381
timestamp 1688980957
transform 1 0 36156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_389
timestamp 1688980957
transform 1 0 36892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_398
timestamp 1688980957
transform 1 0 37720 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_408
timestamp 1688980957
transform 1 0 38640 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_433
timestamp 1688980957
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_445
timestamp 1688980957
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_457
timestamp 1688980957
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_469
timestamp 1688980957
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 1688980957
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_477
timestamp 1688980957
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_489
timestamp 1688980957
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_501
timestamp 1688980957
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_513
timestamp 1688980957
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_525
timestamp 1688980957
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_531
timestamp 1688980957
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_533
timestamp 1688980957
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_545
timestamp 1688980957
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_557
timestamp 1688980957
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_569
timestamp 1688980957
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_581
timestamp 1688980957
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_587
timestamp 1688980957
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 1688980957
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_601
timestamp 1688980957
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_613
timestamp 1688980957
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_625
timestamp 1688980957
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_637
timestamp 1688980957
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_643
timestamp 1688980957
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_645
timestamp 1688980957
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_657
timestamp 1688980957
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_669
timestamp 1688980957
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_681
timestamp 1688980957
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_693
timestamp 1688980957
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_699
timestamp 1688980957
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_701
timestamp 1688980957
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_713
timestamp 1688980957
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_725
timestamp 1688980957
transform 1 0 67804 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_117
timestamp 1688980957
transform 1 0 11868 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_129
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_139
timestamp 1688980957
transform 1 0 13892 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_146
timestamp 1688980957
transform 1 0 14536 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_152
timestamp 1688980957
transform 1 0 15088 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_159
timestamp 1688980957
transform 1 0 15732 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_212
timestamp 1688980957
transform 1 0 20608 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_241
timestamp 1688980957
transform 1 0 23276 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_305
timestamp 1688980957
transform 1 0 29164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_309
timestamp 1688980957
transform 1 0 29532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_341
timestamp 1688980957
transform 1 0 32476 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 1688980957
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 1688980957
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_429
timestamp 1688980957
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_441
timestamp 1688980957
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 1688980957
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_449
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_461
timestamp 1688980957
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_473
timestamp 1688980957
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_485
timestamp 1688980957
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_497
timestamp 1688980957
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_503
timestamp 1688980957
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_505
timestamp 1688980957
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_517
timestamp 1688980957
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_529
timestamp 1688980957
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_541
timestamp 1688980957
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_553
timestamp 1688980957
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_559
timestamp 1688980957
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_561
timestamp 1688980957
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_573
timestamp 1688980957
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_585
timestamp 1688980957
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_597
timestamp 1688980957
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_609
timestamp 1688980957
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_615
timestamp 1688980957
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_617
timestamp 1688980957
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_629
timestamp 1688980957
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_641
timestamp 1688980957
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_653
timestamp 1688980957
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_665
timestamp 1688980957
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_671
timestamp 1688980957
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_673
timestamp 1688980957
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_685
timestamp 1688980957
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_697
timestamp 1688980957
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_709
timestamp 1688980957
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_721
timestamp 1688980957
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_727
timestamp 1688980957
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_729
timestamp 1688980957
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_94
timestamp 1688980957
transform 1 0 9752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_102
timestamp 1688980957
transform 1 0 10488 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_126
timestamp 1688980957
transform 1 0 12696 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_131
timestamp 1688980957
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_175
timestamp 1688980957
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_187
timestamp 1688980957
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_214
timestamp 1688980957
transform 1 0 20792 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_222
timestamp 1688980957
transform 1 0 21528 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_240
timestamp 1688980957
transform 1 0 23184 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_264
timestamp 1688980957
transform 1 0 25392 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_276
timestamp 1688980957
transform 1 0 26496 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_284
timestamp 1688980957
transform 1 0 27232 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_303
timestamp 1688980957
transform 1 0 28980 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_324
timestamp 1688980957
transform 1 0 30912 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_352
timestamp 1688980957
transform 1 0 33488 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_362
timestamp 1688980957
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_377
timestamp 1688980957
transform 1 0 35788 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_394
timestamp 1688980957
transform 1 0 37352 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_406
timestamp 1688980957
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_418
timestamp 1688980957
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_433
timestamp 1688980957
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_445
timestamp 1688980957
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_457
timestamp 1688980957
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_469
timestamp 1688980957
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_475
timestamp 1688980957
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_477
timestamp 1688980957
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_489
timestamp 1688980957
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_501
timestamp 1688980957
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_513
timestamp 1688980957
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_525
timestamp 1688980957
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_531
timestamp 1688980957
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_533
timestamp 1688980957
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_545
timestamp 1688980957
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_557
timestamp 1688980957
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_569
timestamp 1688980957
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_581
timestamp 1688980957
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_587
timestamp 1688980957
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_589
timestamp 1688980957
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_601
timestamp 1688980957
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_613
timestamp 1688980957
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_625
timestamp 1688980957
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_637
timestamp 1688980957
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_643
timestamp 1688980957
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_645
timestamp 1688980957
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_657
timestamp 1688980957
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_669
timestamp 1688980957
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_681
timestamp 1688980957
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_693
timestamp 1688980957
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_699
timestamp 1688980957
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_701
timestamp 1688980957
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_713
timestamp 1688980957
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_725
timestamp 1688980957
transform 1 0 67804 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_73
timestamp 1688980957
transform 1 0 7820 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_97
timestamp 1688980957
transform 1 0 10028 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_130
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_143
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_150
timestamp 1688980957
transform 1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_177
timestamp 1688980957
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_191
timestamp 1688980957
transform 1 0 18676 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_203
timestamp 1688980957
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_229
timestamp 1688980957
transform 1 0 22172 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_233
timestamp 1688980957
transform 1 0 22540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_245
timestamp 1688980957
transform 1 0 23644 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_301
timestamp 1688980957
transform 1 0 28796 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_316
timestamp 1688980957
transform 1 0 30176 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_322
timestamp 1688980957
transform 1 0 30728 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_326
timestamp 1688980957
transform 1 0 31096 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1688980957
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_345
timestamp 1688980957
transform 1 0 32844 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_351
timestamp 1688980957
transform 1 0 33396 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_358
timestamp 1688980957
transform 1 0 34040 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_366
timestamp 1688980957
transform 1 0 34776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_372
timestamp 1688980957
transform 1 0 35328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_389
timestamp 1688980957
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_409
timestamp 1688980957
transform 1 0 38732 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_421
timestamp 1688980957
transform 1 0 39836 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_433
timestamp 1688980957
transform 1 0 40940 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_445
timestamp 1688980957
transform 1 0 42044 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_461
timestamp 1688980957
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_473
timestamp 1688980957
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_485
timestamp 1688980957
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_497
timestamp 1688980957
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_503
timestamp 1688980957
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_505
timestamp 1688980957
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_517
timestamp 1688980957
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_529
timestamp 1688980957
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_541
timestamp 1688980957
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_553
timestamp 1688980957
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_559
timestamp 1688980957
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_561
timestamp 1688980957
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_573
timestamp 1688980957
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_585
timestamp 1688980957
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_597
timestamp 1688980957
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_609
timestamp 1688980957
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_615
timestamp 1688980957
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_617
timestamp 1688980957
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_629
timestamp 1688980957
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_641
timestamp 1688980957
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_653
timestamp 1688980957
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_665
timestamp 1688980957
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_671
timestamp 1688980957
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_673
timestamp 1688980957
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_685
timestamp 1688980957
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_697
timestamp 1688980957
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_709
timestamp 1688980957
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_721
timestamp 1688980957
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_727
timestamp 1688980957
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_729
timestamp 1688980957
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_116
timestamp 1688980957
transform 1 0 11776 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_134
timestamp 1688980957
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_162
timestamp 1688980957
transform 1 0 16008 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_232
timestamp 1688980957
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_258
timestamp 1688980957
transform 1 0 24840 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_303
timestamp 1688980957
transform 1 0 28980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_313
timestamp 1688980957
transform 1 0 29900 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_322
timestamp 1688980957
transform 1 0 30728 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_328
timestamp 1688980957
transform 1 0 31280 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_353
timestamp 1688980957
transform 1 0 33580 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_375
timestamp 1688980957
transform 1 0 35604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_387
timestamp 1688980957
transform 1 0 36708 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_391
timestamp 1688980957
transform 1 0 37076 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_408
timestamp 1688980957
transform 1 0 38640 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_433
timestamp 1688980957
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_445
timestamp 1688980957
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_457
timestamp 1688980957
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_469
timestamp 1688980957
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 1688980957
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_477
timestamp 1688980957
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_489
timestamp 1688980957
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_501
timestamp 1688980957
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_513
timestamp 1688980957
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_525
timestamp 1688980957
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_531
timestamp 1688980957
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_533
timestamp 1688980957
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_545
timestamp 1688980957
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_557
timestamp 1688980957
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_569
timestamp 1688980957
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_581
timestamp 1688980957
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_587
timestamp 1688980957
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_589
timestamp 1688980957
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_601
timestamp 1688980957
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_613
timestamp 1688980957
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_625
timestamp 1688980957
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_637
timestamp 1688980957
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_643
timestamp 1688980957
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_645
timestamp 1688980957
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_657
timestamp 1688980957
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_669
timestamp 1688980957
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_681
timestamp 1688980957
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_693
timestamp 1688980957
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_699
timestamp 1688980957
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_701
timestamp 1688980957
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_713
timestamp 1688980957
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_725
timestamp 1688980957
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_77
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_83
timestamp 1688980957
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_87
timestamp 1688980957
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_97
timestamp 1688980957
transform 1 0 10028 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_134
timestamp 1688980957
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_141
timestamp 1688980957
transform 1 0 14076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_153
timestamp 1688980957
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1688980957
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_175
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_203
timestamp 1688980957
transform 1 0 19780 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_220
timestamp 1688980957
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_246
timestamp 1688980957
transform 1 0 23736 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_258
timestamp 1688980957
transform 1 0 24840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_262
timestamp 1688980957
transform 1 0 25208 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_277
timestamp 1688980957
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_311
timestamp 1688980957
transform 1 0 29716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_328
timestamp 1688980957
transform 1 0 31280 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_367
timestamp 1688980957
transform 1 0 34868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_378
timestamp 1688980957
transform 1 0 35880 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_390
timestamp 1688980957
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1688980957
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 1688980957
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_429
timestamp 1688980957
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_441
timestamp 1688980957
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_447
timestamp 1688980957
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_461
timestamp 1688980957
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_473
timestamp 1688980957
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_485
timestamp 1688980957
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_497
timestamp 1688980957
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_503
timestamp 1688980957
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_505
timestamp 1688980957
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_517
timestamp 1688980957
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_529
timestamp 1688980957
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_541
timestamp 1688980957
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_553
timestamp 1688980957
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_559
timestamp 1688980957
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_561
timestamp 1688980957
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_573
timestamp 1688980957
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_585
timestamp 1688980957
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_597
timestamp 1688980957
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_609
timestamp 1688980957
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_615
timestamp 1688980957
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_617
timestamp 1688980957
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_629
timestamp 1688980957
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_641
timestamp 1688980957
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_653
timestamp 1688980957
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_665
timestamp 1688980957
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_671
timestamp 1688980957
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_673
timestamp 1688980957
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_685
timestamp 1688980957
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_697
timestamp 1688980957
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_709
timestamp 1688980957
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_721
timestamp 1688980957
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_727
timestamp 1688980957
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_729
timestamp 1688980957
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_88
timestamp 1688980957
transform 1 0 9200 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_96
timestamp 1688980957
transform 1 0 9936 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_106
timestamp 1688980957
transform 1 0 10856 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_118
timestamp 1688980957
transform 1 0 11960 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_124
timestamp 1688980957
transform 1 0 12512 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_187
timestamp 1688980957
transform 1 0 18308 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_208
timestamp 1688980957
transform 1 0 20240 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_230
timestamp 1688980957
transform 1 0 22264 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_242
timestamp 1688980957
transform 1 0 23368 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_329
timestamp 1688980957
transform 1 0 31372 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_376
timestamp 1688980957
transform 1 0 35696 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_410
timestamp 1688980957
transform 1 0 38824 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_418
timestamp 1688980957
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_433
timestamp 1688980957
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_445
timestamp 1688980957
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_457
timestamp 1688980957
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_469
timestamp 1688980957
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_475
timestamp 1688980957
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_477
timestamp 1688980957
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_489
timestamp 1688980957
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_501
timestamp 1688980957
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_513
timestamp 1688980957
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_525
timestamp 1688980957
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_531
timestamp 1688980957
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_533
timestamp 1688980957
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_545
timestamp 1688980957
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_557
timestamp 1688980957
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_569
timestamp 1688980957
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_581
timestamp 1688980957
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_587
timestamp 1688980957
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_589
timestamp 1688980957
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_601
timestamp 1688980957
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_613
timestamp 1688980957
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_625
timestamp 1688980957
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_637
timestamp 1688980957
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_643
timestamp 1688980957
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_645
timestamp 1688980957
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_657
timestamp 1688980957
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_669
timestamp 1688980957
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_681
timestamp 1688980957
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_693
timestamp 1688980957
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_699
timestamp 1688980957
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_701
timestamp 1688980957
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_713
timestamp 1688980957
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_725
timestamp 1688980957
transform 1 0 67804 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_73
timestamp 1688980957
transform 1 0 7820 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_131
timestamp 1688980957
transform 1 0 13156 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_148
timestamp 1688980957
transform 1 0 14720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_185
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_198
timestamp 1688980957
transform 1 0 19320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_214
timestamp 1688980957
transform 1 0 20792 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_218
timestamp 1688980957
transform 1 0 21160 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1688980957
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_250
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_268
timestamp 1688980957
transform 1 0 25760 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_292
timestamp 1688980957
transform 1 0 27968 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_303
timestamp 1688980957
transform 1 0 28980 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_314
timestamp 1688980957
transform 1 0 29992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_334
timestamp 1688980957
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_343
timestamp 1688980957
transform 1 0 32660 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_379
timestamp 1688980957
transform 1 0 35972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_387
timestamp 1688980957
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_401
timestamp 1688980957
transform 1 0 37996 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_413
timestamp 1688980957
transform 1 0 39100 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_425
timestamp 1688980957
transform 1 0 40204 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_437
timestamp 1688980957
transform 1 0 41308 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_445
timestamp 1688980957
transform 1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 1688980957
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_461
timestamp 1688980957
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_473
timestamp 1688980957
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_485
timestamp 1688980957
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_497
timestamp 1688980957
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_503
timestamp 1688980957
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_505
timestamp 1688980957
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_517
timestamp 1688980957
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_529
timestamp 1688980957
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_541
timestamp 1688980957
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_553
timestamp 1688980957
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_559
timestamp 1688980957
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_561
timestamp 1688980957
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_573
timestamp 1688980957
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_585
timestamp 1688980957
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_597
timestamp 1688980957
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_609
timestamp 1688980957
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_615
timestamp 1688980957
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_617
timestamp 1688980957
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_629
timestamp 1688980957
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_641
timestamp 1688980957
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_653
timestamp 1688980957
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_665
timestamp 1688980957
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_671
timestamp 1688980957
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_673
timestamp 1688980957
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_685
timestamp 1688980957
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_697
timestamp 1688980957
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_709
timestamp 1688980957
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_721
timestamp 1688980957
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_727
timestamp 1688980957
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_729
timestamp 1688980957
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_88
timestamp 1688980957
transform 1 0 9200 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_96
timestamp 1688980957
transform 1 0 9936 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_105
timestamp 1688980957
transform 1 0 10764 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_117
timestamp 1688980957
transform 1 0 11868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_132
timestamp 1688980957
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_162
timestamp 1688980957
transform 1 0 16008 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_175
timestamp 1688980957
transform 1 0 17204 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_205
timestamp 1688980957
transform 1 0 19964 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_210
timestamp 1688980957
transform 1 0 20424 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_222
timestamp 1688980957
transform 1 0 21528 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_234
timestamp 1688980957
transform 1 0 22632 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_243
timestamp 1688980957
transform 1 0 23460 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_287
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_300
timestamp 1688980957
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_331
timestamp 1688980957
transform 1 0 31556 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_362
timestamp 1688980957
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_388
timestamp 1688980957
transform 1 0 36800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_406
timestamp 1688980957
transform 1 0 38456 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_418
timestamp 1688980957
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_421
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_433
timestamp 1688980957
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_445
timestamp 1688980957
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_457
timestamp 1688980957
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_469
timestamp 1688980957
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_475
timestamp 1688980957
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_477
timestamp 1688980957
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_489
timestamp 1688980957
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_501
timestamp 1688980957
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_513
timestamp 1688980957
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_525
timestamp 1688980957
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_531
timestamp 1688980957
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_533
timestamp 1688980957
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_545
timestamp 1688980957
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_557
timestamp 1688980957
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_569
timestamp 1688980957
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_581
timestamp 1688980957
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_587
timestamp 1688980957
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_589
timestamp 1688980957
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_601
timestamp 1688980957
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_613
timestamp 1688980957
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_625
timestamp 1688980957
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_637
timestamp 1688980957
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_643
timestamp 1688980957
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_645
timestamp 1688980957
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_657
timestamp 1688980957
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_669
timestamp 1688980957
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_681
timestamp 1688980957
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_693
timestamp 1688980957
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_699
timestamp 1688980957
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_701
timestamp 1688980957
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_713
timestamp 1688980957
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_725
timestamp 1688980957
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_73
timestamp 1688980957
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_94
timestamp 1688980957
transform 1 0 9752 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_118
timestamp 1688980957
transform 1 0 11960 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_129
timestamp 1688980957
transform 1 0 12972 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_151
timestamp 1688980957
transform 1 0 14996 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_163
timestamp 1688980957
transform 1 0 16100 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_177
timestamp 1688980957
transform 1 0 17388 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_190
timestamp 1688980957
transform 1 0 18584 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_198
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_238
timestamp 1688980957
transform 1 0 23000 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_250
timestamp 1688980957
transform 1 0 24104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_254
timestamp 1688980957
transform 1 0 24472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_275
timestamp 1688980957
transform 1 0 26404 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_327
timestamp 1688980957
transform 1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_345
timestamp 1688980957
transform 1 0 32844 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_360
timestamp 1688980957
transform 1 0 34224 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_372
timestamp 1688980957
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_376
timestamp 1688980957
transform 1 0 35696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_384
timestamp 1688980957
transform 1 0 36432 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_389
timestamp 1688980957
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 1688980957
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 1688980957
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_429
timestamp 1688980957
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_441
timestamp 1688980957
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 1688980957
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_449
timestamp 1688980957
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_461
timestamp 1688980957
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_473
timestamp 1688980957
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_485
timestamp 1688980957
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_497
timestamp 1688980957
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_503
timestamp 1688980957
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_505
timestamp 1688980957
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_517
timestamp 1688980957
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_529
timestamp 1688980957
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_541
timestamp 1688980957
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_553
timestamp 1688980957
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_559
timestamp 1688980957
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_561
timestamp 1688980957
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_573
timestamp 1688980957
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_585
timestamp 1688980957
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_597
timestamp 1688980957
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_609
timestamp 1688980957
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 1688980957
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_617
timestamp 1688980957
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_629
timestamp 1688980957
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_641
timestamp 1688980957
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_653
timestamp 1688980957
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_665
timestamp 1688980957
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_671
timestamp 1688980957
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_673
timestamp 1688980957
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_685
timestamp 1688980957
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_697
timestamp 1688980957
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_709
timestamp 1688980957
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_721
timestamp 1688980957
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_727
timestamp 1688980957
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_729
timestamp 1688980957
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_92
timestamp 1688980957
transform 1 0 9568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_114
timestamp 1688980957
transform 1 0 11592 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_164
timestamp 1688980957
transform 1 0 16192 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_238
timestamp 1688980957
transform 1 0 23000 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 1688980957
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_258
timestamp 1688980957
transform 1 0 24840 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_288
timestamp 1688980957
transform 1 0 27600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_299
timestamp 1688980957
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_323
timestamp 1688980957
transform 1 0 30820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_331
timestamp 1688980957
transform 1 0 31556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_341
timestamp 1688980957
transform 1 0 32476 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_396
timestamp 1688980957
transform 1 0 37536 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_408
timestamp 1688980957
transform 1 0 38640 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_433
timestamp 1688980957
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_445
timestamp 1688980957
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_457
timestamp 1688980957
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_469
timestamp 1688980957
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_475
timestamp 1688980957
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_477
timestamp 1688980957
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_489
timestamp 1688980957
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_501
timestamp 1688980957
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_513
timestamp 1688980957
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_525
timestamp 1688980957
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_531
timestamp 1688980957
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_533
timestamp 1688980957
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_545
timestamp 1688980957
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_557
timestamp 1688980957
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_569
timestamp 1688980957
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_581
timestamp 1688980957
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_587
timestamp 1688980957
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_589
timestamp 1688980957
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_601
timestamp 1688980957
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_613
timestamp 1688980957
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_625
timestamp 1688980957
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_637
timestamp 1688980957
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_643
timestamp 1688980957
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_645
timestamp 1688980957
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_657
timestamp 1688980957
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_669
timestamp 1688980957
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_681
timestamp 1688980957
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_693
timestamp 1688980957
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_699
timestamp 1688980957
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_701
timestamp 1688980957
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_713
timestamp 1688980957
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_725
timestamp 1688980957
transform 1 0 67804 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_77
timestamp 1688980957
transform 1 0 8188 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_98
timestamp 1688980957
transform 1 0 10120 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_124
timestamp 1688980957
transform 1 0 12512 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_133
timestamp 1688980957
transform 1 0 13340 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_139
timestamp 1688980957
transform 1 0 13892 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_156
timestamp 1688980957
transform 1 0 15456 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_164
timestamp 1688980957
transform 1 0 16192 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_203
timestamp 1688980957
transform 1 0 19780 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_212
timestamp 1688980957
transform 1 0 20608 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_228
timestamp 1688980957
transform 1 0 22080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_269
timestamp 1688980957
transform 1 0 25852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 1688980957
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_299
timestamp 1688980957
transform 1 0 28612 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_312
timestamp 1688980957
transform 1 0 29808 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_320
timestamp 1688980957
transform 1 0 30544 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_326
timestamp 1688980957
transform 1 0 31096 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_348
timestamp 1688980957
transform 1 0 33120 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_401
timestamp 1688980957
transform 1 0 37996 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_413
timestamp 1688980957
transform 1 0 39100 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_425
timestamp 1688980957
transform 1 0 40204 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_437
timestamp 1688980957
transform 1 0 41308 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_445
timestamp 1688980957
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_461
timestamp 1688980957
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_473
timestamp 1688980957
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_485
timestamp 1688980957
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_497
timestamp 1688980957
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 1688980957
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_505
timestamp 1688980957
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_517
timestamp 1688980957
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_529
timestamp 1688980957
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_541
timestamp 1688980957
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_553
timestamp 1688980957
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_559
timestamp 1688980957
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_561
timestamp 1688980957
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_573
timestamp 1688980957
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_585
timestamp 1688980957
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_597
timestamp 1688980957
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_609
timestamp 1688980957
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_615
timestamp 1688980957
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_617
timestamp 1688980957
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_629
timestamp 1688980957
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_641
timestamp 1688980957
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_653
timestamp 1688980957
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_665
timestamp 1688980957
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_671
timestamp 1688980957
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_673
timestamp 1688980957
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_685
timestamp 1688980957
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_697
timestamp 1688980957
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_709
timestamp 1688980957
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_721
timestamp 1688980957
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_727
timestamp 1688980957
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_729
timestamp 1688980957
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_118
timestamp 1688980957
transform 1 0 11960 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_167
timestamp 1688980957
transform 1 0 16468 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_193
timestamp 1688980957
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_217
timestamp 1688980957
transform 1 0 21068 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_225
timestamp 1688980957
transform 1 0 21804 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_237
timestamp 1688980957
transform 1 0 22908 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 1688980957
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_269
timestamp 1688980957
transform 1 0 25852 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_294
timestamp 1688980957
transform 1 0 28152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_298
timestamp 1688980957
transform 1 0 28520 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_340
timestamp 1688980957
transform 1 0 32384 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1688980957
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_383
timestamp 1688980957
transform 1 0 36340 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_395
timestamp 1688980957
transform 1 0 37444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_407
timestamp 1688980957
transform 1 0 38548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1688980957
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 1688980957
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 1688980957
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_457
timestamp 1688980957
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_469
timestamp 1688980957
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_475
timestamp 1688980957
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_477
timestamp 1688980957
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_489
timestamp 1688980957
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_501
timestamp 1688980957
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_513
timestamp 1688980957
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 1688980957
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 1688980957
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 1688980957
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_545
timestamp 1688980957
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_557
timestamp 1688980957
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_569
timestamp 1688980957
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_581
timestamp 1688980957
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_587
timestamp 1688980957
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_589
timestamp 1688980957
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_601
timestamp 1688980957
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_613
timestamp 1688980957
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_625
timestamp 1688980957
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_637
timestamp 1688980957
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_643
timestamp 1688980957
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_645
timestamp 1688980957
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_657
timestamp 1688980957
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_669
timestamp 1688980957
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_681
timestamp 1688980957
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_693
timestamp 1688980957
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_699
timestamp 1688980957
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_701
timestamp 1688980957
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_713
timestamp 1688980957
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_725
timestamp 1688980957
transform 1 0 67804 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_117
timestamp 1688980957
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_121
timestamp 1688980957
transform 1 0 12236 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_131
timestamp 1688980957
transform 1 0 13156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_139
timestamp 1688980957
transform 1 0 13892 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_160
timestamp 1688980957
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_211
timestamp 1688980957
transform 1 0 20516 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_228
timestamp 1688980957
transform 1 0 22080 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_232
timestamp 1688980957
transform 1 0 22448 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_236
timestamp 1688980957
transform 1 0 22816 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_242
timestamp 1688980957
transform 1 0 23368 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_254
timestamp 1688980957
transform 1 0 24472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_268
timestamp 1688980957
transform 1 0 25760 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_276
timestamp 1688980957
transform 1 0 26496 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_296
timestamp 1688980957
transform 1 0 28336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_304
timestamp 1688980957
transform 1 0 29072 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_308
timestamp 1688980957
transform 1 0 29440 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_312
timestamp 1688980957
transform 1 0 29808 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_318
timestamp 1688980957
transform 1 0 30360 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_330
timestamp 1688980957
transform 1 0 31464 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1688980957
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1688980957
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 1688980957
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 1688980957
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 1688980957
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 1688980957
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_461
timestamp 1688980957
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_473
timestamp 1688980957
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_485
timestamp 1688980957
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_497
timestamp 1688980957
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 1688980957
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_505
timestamp 1688980957
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_517
timestamp 1688980957
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_529
timestamp 1688980957
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_541
timestamp 1688980957
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_553
timestamp 1688980957
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_559
timestamp 1688980957
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_561
timestamp 1688980957
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_573
timestamp 1688980957
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_585
timestamp 1688980957
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_597
timestamp 1688980957
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_609
timestamp 1688980957
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_615
timestamp 1688980957
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_617
timestamp 1688980957
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_629
timestamp 1688980957
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_641
timestamp 1688980957
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_653
timestamp 1688980957
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_665
timestamp 1688980957
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_671
timestamp 1688980957
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_673
timestamp 1688980957
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_685
timestamp 1688980957
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_697
timestamp 1688980957
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_709
timestamp 1688980957
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_721
timestamp 1688980957
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_727
timestamp 1688980957
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_729
timestamp 1688980957
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_117
timestamp 1688980957
transform 1 0 11868 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_144
timestamp 1688980957
transform 1 0 14352 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_156
timestamp 1688980957
transform 1 0 15456 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_168
timestamp 1688980957
transform 1 0 16560 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_180
timestamp 1688980957
transform 1 0 17664 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_188
timestamp 1688980957
transform 1 0 18400 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1688980957
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_218
timestamp 1688980957
transform 1 0 21160 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_228
timestamp 1688980957
transform 1 0 22080 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_240
timestamp 1688980957
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_285
timestamp 1688980957
transform 1 0 27324 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_293
timestamp 1688980957
transform 1 0 28060 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_316
timestamp 1688980957
transform 1 0 30176 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_326
timestamp 1688980957
transform 1 0 31096 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_338
timestamp 1688980957
transform 1 0 32200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_353
timestamp 1688980957
transform 1 0 33580 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_361
timestamp 1688980957
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1688980957
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 1688980957
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 1688980957
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 1688980957
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 1688980957
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_457
timestamp 1688980957
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_469
timestamp 1688980957
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_475
timestamp 1688980957
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_477
timestamp 1688980957
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_489
timestamp 1688980957
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_501
timestamp 1688980957
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_513
timestamp 1688980957
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_525
timestamp 1688980957
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_531
timestamp 1688980957
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_533
timestamp 1688980957
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_545
timestamp 1688980957
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_557
timestamp 1688980957
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_569
timestamp 1688980957
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_581
timestamp 1688980957
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_587
timestamp 1688980957
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 1688980957
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 1688980957
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_613
timestamp 1688980957
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_625
timestamp 1688980957
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_637
timestamp 1688980957
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_643
timestamp 1688980957
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_645
timestamp 1688980957
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_657
timestamp 1688980957
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_669
timestamp 1688980957
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_681
timestamp 1688980957
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_693
timestamp 1688980957
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_699
timestamp 1688980957
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_701
timestamp 1688980957
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_713
timestamp 1688980957
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_725
timestamp 1688980957
transform 1 0 67804 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_229
timestamp 1688980957
transform 1 0 22172 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_248
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_270
timestamp 1688980957
transform 1 0 25944 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_276
timestamp 1688980957
transform 1 0 26496 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_307
timestamp 1688980957
transform 1 0 29348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_341
timestamp 1688980957
transform 1 0 32476 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_366
timestamp 1688980957
transform 1 0 34776 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_378
timestamp 1688980957
transform 1 0 35880 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_390
timestamp 1688980957
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1688980957
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 1688980957
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 1688980957
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 1688980957
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 1688980957
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_461
timestamp 1688980957
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_473
timestamp 1688980957
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_485
timestamp 1688980957
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_497
timestamp 1688980957
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 1688980957
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_505
timestamp 1688980957
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_517
timestamp 1688980957
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_529
timestamp 1688980957
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_541
timestamp 1688980957
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_553
timestamp 1688980957
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 1688980957
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_561
timestamp 1688980957
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_573
timestamp 1688980957
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_585
timestamp 1688980957
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_597
timestamp 1688980957
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_609
timestamp 1688980957
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_615
timestamp 1688980957
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_617
timestamp 1688980957
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_629
timestamp 1688980957
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_641
timestamp 1688980957
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_653
timestamp 1688980957
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_665
timestamp 1688980957
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_671
timestamp 1688980957
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_673
timestamp 1688980957
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_685
timestamp 1688980957
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_697
timestamp 1688980957
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_709
timestamp 1688980957
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_721
timestamp 1688980957
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_727
timestamp 1688980957
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_729
timestamp 1688980957
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_213
timestamp 1688980957
transform 1 0 20700 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_217
timestamp 1688980957
transform 1 0 21068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_229
timestamp 1688980957
transform 1 0 22172 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_244
timestamp 1688980957
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_267
timestamp 1688980957
transform 1 0 25668 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_271
timestamp 1688980957
transform 1 0 26036 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_288
timestamp 1688980957
transform 1 0 27600 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_320
timestamp 1688980957
transform 1 0 30544 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_332
timestamp 1688980957
transform 1 0 31648 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_344
timestamp 1688980957
transform 1 0 32752 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_356
timestamp 1688980957
transform 1 0 33856 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_401
timestamp 1688980957
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_413
timestamp 1688980957
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 1688980957
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 1688980957
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_445
timestamp 1688980957
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_457
timestamp 1688980957
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_469
timestamp 1688980957
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_475
timestamp 1688980957
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 1688980957
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 1688980957
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_501
timestamp 1688980957
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_513
timestamp 1688980957
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_525
timestamp 1688980957
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_531
timestamp 1688980957
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 1688980957
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_545
timestamp 1688980957
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_557
timestamp 1688980957
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_569
timestamp 1688980957
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_581
timestamp 1688980957
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_587
timestamp 1688980957
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 1688980957
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 1688980957
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_613
timestamp 1688980957
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_625
timestamp 1688980957
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_637
timestamp 1688980957
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_643
timestamp 1688980957
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_645
timestamp 1688980957
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_657
timestamp 1688980957
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_669
timestamp 1688980957
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_681
timestamp 1688980957
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_693
timestamp 1688980957
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_699
timestamp 1688980957
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_701
timestamp 1688980957
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_713
timestamp 1688980957
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_725
timestamp 1688980957
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_209
timestamp 1688980957
transform 1 0 20332 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_268
timestamp 1688980957
transform 1 0 25760 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 1688980957
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 1688980957
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1688980957
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 1688980957
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 1688980957
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_429
timestamp 1688980957
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_441
timestamp 1688980957
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_447
timestamp 1688980957
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_449
timestamp 1688980957
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_461
timestamp 1688980957
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_473
timestamp 1688980957
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_485
timestamp 1688980957
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_497
timestamp 1688980957
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_503
timestamp 1688980957
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_505
timestamp 1688980957
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_517
timestamp 1688980957
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_529
timestamp 1688980957
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_541
timestamp 1688980957
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_553
timestamp 1688980957
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_559
timestamp 1688980957
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_561
timestamp 1688980957
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_573
timestamp 1688980957
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_585
timestamp 1688980957
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_597
timestamp 1688980957
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_609
timestamp 1688980957
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_615
timestamp 1688980957
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_617
timestamp 1688980957
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_629
timestamp 1688980957
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_641
timestamp 1688980957
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_653
timestamp 1688980957
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_665
timestamp 1688980957
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_671
timestamp 1688980957
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_673
timestamp 1688980957
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_685
timestamp 1688980957
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_697
timestamp 1688980957
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_709
timestamp 1688980957
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_721
timestamp 1688980957
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_727
timestamp 1688980957
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_205
timestamp 1688980957
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_250
timestamp 1688980957
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_276
timestamp 1688980957
transform 1 0 26496 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_288
timestamp 1688980957
transform 1 0 27600 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_300
timestamp 1688980957
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1688980957
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 1688980957
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 1688980957
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_401
timestamp 1688980957
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_413
timestamp 1688980957
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 1688980957
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 1688980957
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_433
timestamp 1688980957
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_445
timestamp 1688980957
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_457
timestamp 1688980957
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_469
timestamp 1688980957
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_475
timestamp 1688980957
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_477
timestamp 1688980957
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_489
timestamp 1688980957
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_501
timestamp 1688980957
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_513
timestamp 1688980957
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_525
timestamp 1688980957
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_531
timestamp 1688980957
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_533
timestamp 1688980957
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_545
timestamp 1688980957
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_557
timestamp 1688980957
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_569
timestamp 1688980957
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_581
timestamp 1688980957
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_587
timestamp 1688980957
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_589
timestamp 1688980957
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_601
timestamp 1688980957
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_613
timestamp 1688980957
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_625
timestamp 1688980957
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_637
timestamp 1688980957
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_643
timestamp 1688980957
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_645
timestamp 1688980957
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_657
timestamp 1688980957
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_669
timestamp 1688980957
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_681
timestamp 1688980957
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_693
timestamp 1688980957
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_699
timestamp 1688980957
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_701
timestamp 1688980957
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_713
timestamp 1688980957
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_725
timestamp 1688980957
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_213
timestamp 1688980957
transform 1 0 20700 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_219
timestamp 1688980957
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_233
timestamp 1688980957
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_252
timestamp 1688980957
transform 1 0 24288 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_256
timestamp 1688980957
transform 1 0 24656 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_260
timestamp 1688980957
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_272
timestamp 1688980957
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1688980957
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 1688980957
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 1688980957
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1688980957
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_405
timestamp 1688980957
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_417
timestamp 1688980957
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_429
timestamp 1688980957
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_441
timestamp 1688980957
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_447
timestamp 1688980957
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_449
timestamp 1688980957
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_461
timestamp 1688980957
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_473
timestamp 1688980957
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_485
timestamp 1688980957
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_497
timestamp 1688980957
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_503
timestamp 1688980957
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_505
timestamp 1688980957
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_517
timestamp 1688980957
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_529
timestamp 1688980957
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_541
timestamp 1688980957
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_553
timestamp 1688980957
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_559
timestamp 1688980957
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_561
timestamp 1688980957
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_573
timestamp 1688980957
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_585
timestamp 1688980957
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_597
timestamp 1688980957
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_609
timestamp 1688980957
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_615
timestamp 1688980957
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_617
timestamp 1688980957
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_629
timestamp 1688980957
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_641
timestamp 1688980957
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_653
timestamp 1688980957
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_665
timestamp 1688980957
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_671
timestamp 1688980957
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_673
timestamp 1688980957
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_685
timestamp 1688980957
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_697
timestamp 1688980957
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_709
timestamp 1688980957
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_721
timestamp 1688980957
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_727
timestamp 1688980957
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_729
timestamp 1688980957
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1688980957
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 1688980957
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 1688980957
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_401
timestamp 1688980957
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_413
timestamp 1688980957
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_419
timestamp 1688980957
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 1688980957
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 1688980957
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_445
timestamp 1688980957
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_457
timestamp 1688980957
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_469
timestamp 1688980957
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_475
timestamp 1688980957
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_477
timestamp 1688980957
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_489
timestamp 1688980957
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_501
timestamp 1688980957
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_513
timestamp 1688980957
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_525
timestamp 1688980957
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_531
timestamp 1688980957
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_533
timestamp 1688980957
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_545
timestamp 1688980957
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_557
timestamp 1688980957
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_569
timestamp 1688980957
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_581
timestamp 1688980957
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_587
timestamp 1688980957
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_589
timestamp 1688980957
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_601
timestamp 1688980957
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_613
timestamp 1688980957
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_625
timestamp 1688980957
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_637
timestamp 1688980957
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_643
timestamp 1688980957
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_645
timestamp 1688980957
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_657
timestamp 1688980957
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_669
timestamp 1688980957
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_681
timestamp 1688980957
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_693
timestamp 1688980957
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_699
timestamp 1688980957
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_701
timestamp 1688980957
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_713
timestamp 1688980957
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_725
timestamp 1688980957
transform 1 0 67804 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1688980957
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1688980957
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1688980957
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 1688980957
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_429
timestamp 1688980957
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_441
timestamp 1688980957
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_447
timestamp 1688980957
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_449
timestamp 1688980957
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_461
timestamp 1688980957
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_473
timestamp 1688980957
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_485
timestamp 1688980957
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_497
timestamp 1688980957
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_503
timestamp 1688980957
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_505
timestamp 1688980957
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_517
timestamp 1688980957
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_529
timestamp 1688980957
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_541
timestamp 1688980957
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_553
timestamp 1688980957
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_559
timestamp 1688980957
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_561
timestamp 1688980957
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_573
timestamp 1688980957
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_585
timestamp 1688980957
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_597
timestamp 1688980957
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_609
timestamp 1688980957
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_615
timestamp 1688980957
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_617
timestamp 1688980957
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_629
timestamp 1688980957
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_641
timestamp 1688980957
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_653
timestamp 1688980957
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_665
timestamp 1688980957
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_671
timestamp 1688980957
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_673
timestamp 1688980957
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_685
timestamp 1688980957
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_697
timestamp 1688980957
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_709
timestamp 1688980957
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_721
timestamp 1688980957
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_727
timestamp 1688980957
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_729
timestamp 1688980957
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1688980957
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1688980957
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_401
timestamp 1688980957
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_413
timestamp 1688980957
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 1688980957
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 1688980957
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_433
timestamp 1688980957
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_445
timestamp 1688980957
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_457
timestamp 1688980957
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_469
timestamp 1688980957
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_475
timestamp 1688980957
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_477
timestamp 1688980957
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_489
timestamp 1688980957
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_501
timestamp 1688980957
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_513
timestamp 1688980957
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_525
timestamp 1688980957
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_531
timestamp 1688980957
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_533
timestamp 1688980957
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_545
timestamp 1688980957
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_557
timestamp 1688980957
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_569
timestamp 1688980957
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_581
timestamp 1688980957
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_587
timestamp 1688980957
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_589
timestamp 1688980957
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_601
timestamp 1688980957
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_613
timestamp 1688980957
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_625
timestamp 1688980957
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_637
timestamp 1688980957
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_643
timestamp 1688980957
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_645
timestamp 1688980957
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_657
timestamp 1688980957
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_669
timestamp 1688980957
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_681
timestamp 1688980957
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_693
timestamp 1688980957
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_699
timestamp 1688980957
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_701
timestamp 1688980957
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_713
timestamp 1688980957
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_725
timestamp 1688980957
transform 1 0 67804 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1688980957
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 1688980957
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1688980957
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 1688980957
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 1688980957
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_429
timestamp 1688980957
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_441
timestamp 1688980957
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_447
timestamp 1688980957
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 1688980957
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_461
timestamp 1688980957
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_473
timestamp 1688980957
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_485
timestamp 1688980957
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_497
timestamp 1688980957
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_503
timestamp 1688980957
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_505
timestamp 1688980957
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_517
timestamp 1688980957
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_529
timestamp 1688980957
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_541
timestamp 1688980957
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_553
timestamp 1688980957
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_559
timestamp 1688980957
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_561
timestamp 1688980957
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_573
timestamp 1688980957
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_585
timestamp 1688980957
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_597
timestamp 1688980957
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_609
timestamp 1688980957
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_615
timestamp 1688980957
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_617
timestamp 1688980957
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_629
timestamp 1688980957
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_641
timestamp 1688980957
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_653
timestamp 1688980957
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_665
timestamp 1688980957
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_671
timestamp 1688980957
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_673
timestamp 1688980957
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_685
timestamp 1688980957
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_697
timestamp 1688980957
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_709
timestamp 1688980957
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_721
timestamp 1688980957
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_727
timestamp 1688980957
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_729
timestamp 1688980957
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 1688980957
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1688980957
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_401
timestamp 1688980957
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_413
timestamp 1688980957
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 1688980957
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1688980957
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 1688980957
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 1688980957
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_457
timestamp 1688980957
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_469
timestamp 1688980957
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_475
timestamp 1688980957
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_477
timestamp 1688980957
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_489
timestamp 1688980957
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_501
timestamp 1688980957
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_513
timestamp 1688980957
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_525
timestamp 1688980957
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_531
timestamp 1688980957
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_533
timestamp 1688980957
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_545
timestamp 1688980957
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_557
timestamp 1688980957
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_569
timestamp 1688980957
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_581
timestamp 1688980957
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_587
timestamp 1688980957
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_589
timestamp 1688980957
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_601
timestamp 1688980957
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_613
timestamp 1688980957
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_625
timestamp 1688980957
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_637
timestamp 1688980957
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_643
timestamp 1688980957
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_645
timestamp 1688980957
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_657
timestamp 1688980957
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_669
timestamp 1688980957
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_681
timestamp 1688980957
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_693
timestamp 1688980957
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_699
timestamp 1688980957
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_701
timestamp 1688980957
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_713
timestamp 1688980957
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_725
timestamp 1688980957
transform 1 0 67804 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1688980957
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 1688980957
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1688980957
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1688980957
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1688980957
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 1688980957
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_441
timestamp 1688980957
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_447
timestamp 1688980957
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 1688980957
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_461
timestamp 1688980957
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_473
timestamp 1688980957
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_485
timestamp 1688980957
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_497
timestamp 1688980957
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_503
timestamp 1688980957
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_505
timestamp 1688980957
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_517
timestamp 1688980957
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_529
timestamp 1688980957
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_541
timestamp 1688980957
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_553
timestamp 1688980957
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_559
timestamp 1688980957
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_561
timestamp 1688980957
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_573
timestamp 1688980957
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_585
timestamp 1688980957
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_597
timestamp 1688980957
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_609
timestamp 1688980957
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_615
timestamp 1688980957
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_617
timestamp 1688980957
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_629
timestamp 1688980957
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_641
timestamp 1688980957
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_653
timestamp 1688980957
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_665
timestamp 1688980957
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_671
timestamp 1688980957
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_673
timestamp 1688980957
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_685
timestamp 1688980957
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_697
timestamp 1688980957
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_709
timestamp 1688980957
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_721
timestamp 1688980957
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_727
timestamp 1688980957
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_729
timestamp 1688980957
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1688980957
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1688980957
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 1688980957
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 1688980957
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 1688980957
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_421
timestamp 1688980957
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_433
timestamp 1688980957
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_445
timestamp 1688980957
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_457
timestamp 1688980957
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_469
timestamp 1688980957
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_475
timestamp 1688980957
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_477
timestamp 1688980957
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_489
timestamp 1688980957
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_501
timestamp 1688980957
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_513
timestamp 1688980957
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_525
timestamp 1688980957
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_531
timestamp 1688980957
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_533
timestamp 1688980957
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_545
timestamp 1688980957
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_557
timestamp 1688980957
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_569
timestamp 1688980957
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_581
timestamp 1688980957
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_587
timestamp 1688980957
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_589
timestamp 1688980957
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_601
timestamp 1688980957
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_613
timestamp 1688980957
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_625
timestamp 1688980957
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_637
timestamp 1688980957
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_643
timestamp 1688980957
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_645
timestamp 1688980957
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_657
timestamp 1688980957
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_669
timestamp 1688980957
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_681
timestamp 1688980957
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_693
timestamp 1688980957
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_699
timestamp 1688980957
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_701
timestamp 1688980957
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_713
timestamp 1688980957
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_725
timestamp 1688980957
transform 1 0 67804 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1688980957
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1688980957
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1688980957
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1688980957
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1688980957
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_429
timestamp 1688980957
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_441
timestamp 1688980957
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 1688980957
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_449
timestamp 1688980957
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_461
timestamp 1688980957
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_473
timestamp 1688980957
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_485
timestamp 1688980957
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_497
timestamp 1688980957
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_503
timestamp 1688980957
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_505
timestamp 1688980957
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_517
timestamp 1688980957
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_529
timestamp 1688980957
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_541
timestamp 1688980957
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_553
timestamp 1688980957
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_559
timestamp 1688980957
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_561
timestamp 1688980957
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_573
timestamp 1688980957
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_585
timestamp 1688980957
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_597
timestamp 1688980957
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_609
timestamp 1688980957
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_615
timestamp 1688980957
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_617
timestamp 1688980957
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_629
timestamp 1688980957
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_641
timestamp 1688980957
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_653
timestamp 1688980957
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_665
timestamp 1688980957
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_671
timestamp 1688980957
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_673
timestamp 1688980957
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_685
timestamp 1688980957
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_697
timestamp 1688980957
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_709
timestamp 1688980957
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_721
timestamp 1688980957
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_727
timestamp 1688980957
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_729
timestamp 1688980957
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1688980957
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1688980957
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 1688980957
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1688980957
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1688980957
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_433
timestamp 1688980957
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_445
timestamp 1688980957
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_457
timestamp 1688980957
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_469
timestamp 1688980957
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_475
timestamp 1688980957
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_477
timestamp 1688980957
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_489
timestamp 1688980957
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_501
timestamp 1688980957
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_513
timestamp 1688980957
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_525
timestamp 1688980957
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_531
timestamp 1688980957
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_533
timestamp 1688980957
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_545
timestamp 1688980957
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_557
timestamp 1688980957
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_569
timestamp 1688980957
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_581
timestamp 1688980957
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_587
timestamp 1688980957
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_589
timestamp 1688980957
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_601
timestamp 1688980957
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_613
timestamp 1688980957
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_625
timestamp 1688980957
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_637
timestamp 1688980957
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_643
timestamp 1688980957
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_645
timestamp 1688980957
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_657
timestamp 1688980957
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_669
timestamp 1688980957
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_681
timestamp 1688980957
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_693
timestamp 1688980957
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_699
timestamp 1688980957
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_701
timestamp 1688980957
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_713
timestamp 1688980957
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_725
timestamp 1688980957
transform 1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1688980957
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1688980957
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1688980957
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 1688980957
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 1688980957
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 1688980957
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 1688980957
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_461
timestamp 1688980957
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_473
timestamp 1688980957
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_485
timestamp 1688980957
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_497
timestamp 1688980957
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_503
timestamp 1688980957
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_505
timestamp 1688980957
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_517
timestamp 1688980957
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_529
timestamp 1688980957
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_541
timestamp 1688980957
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_553
timestamp 1688980957
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_559
timestamp 1688980957
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_561
timestamp 1688980957
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_573
timestamp 1688980957
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_585
timestamp 1688980957
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_597
timestamp 1688980957
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_609
timestamp 1688980957
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_615
timestamp 1688980957
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_617
timestamp 1688980957
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_629
timestamp 1688980957
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_641
timestamp 1688980957
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_653
timestamp 1688980957
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_665
timestamp 1688980957
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_671
timestamp 1688980957
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_673
timestamp 1688980957
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_685
timestamp 1688980957
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_697
timestamp 1688980957
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_709
timestamp 1688980957
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_721
timestamp 1688980957
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_727
timestamp 1688980957
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_729
timestamp 1688980957
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1688980957
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 1688980957
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 1688980957
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1688980957
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 1688980957
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 1688980957
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_457
timestamp 1688980957
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_469
timestamp 1688980957
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_475
timestamp 1688980957
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_477
timestamp 1688980957
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_489
timestamp 1688980957
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_501
timestamp 1688980957
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_513
timestamp 1688980957
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_525
timestamp 1688980957
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_531
timestamp 1688980957
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_533
timestamp 1688980957
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_545
timestamp 1688980957
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_557
timestamp 1688980957
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_569
timestamp 1688980957
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_581
timestamp 1688980957
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_587
timestamp 1688980957
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_589
timestamp 1688980957
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_601
timestamp 1688980957
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_613
timestamp 1688980957
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_625
timestamp 1688980957
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_637
timestamp 1688980957
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_643
timestamp 1688980957
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_645
timestamp 1688980957
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_657
timestamp 1688980957
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_669
timestamp 1688980957
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_681
timestamp 1688980957
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_693
timestamp 1688980957
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_699
timestamp 1688980957
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_701
timestamp 1688980957
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_713
timestamp 1688980957
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_725
timestamp 1688980957
transform 1 0 67804 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1688980957
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1688980957
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1688980957
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 1688980957
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 1688980957
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 1688980957
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1688980957
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 1688980957
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_473
timestamp 1688980957
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_485
timestamp 1688980957
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_497
timestamp 1688980957
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_503
timestamp 1688980957
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_505
timestamp 1688980957
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_517
timestamp 1688980957
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_529
timestamp 1688980957
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_541
timestamp 1688980957
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_553
timestamp 1688980957
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_559
timestamp 1688980957
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_561
timestamp 1688980957
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_573
timestamp 1688980957
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_585
timestamp 1688980957
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_597
timestamp 1688980957
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_609
timestamp 1688980957
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_615
timestamp 1688980957
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_617
timestamp 1688980957
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_629
timestamp 1688980957
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_641
timestamp 1688980957
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_653
timestamp 1688980957
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_665
timestamp 1688980957
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_671
timestamp 1688980957
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_673
timestamp 1688980957
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_685
timestamp 1688980957
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_697
timestamp 1688980957
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_709
timestamp 1688980957
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_721
timestamp 1688980957
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_727
timestamp 1688980957
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_729
timestamp 1688980957
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1688980957
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1688980957
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1688980957
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1688980957
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1688980957
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1688980957
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1688980957
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1688980957
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1688980957
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 1688980957
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_445
timestamp 1688980957
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_457
timestamp 1688980957
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_469
timestamp 1688980957
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_475
timestamp 1688980957
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_477
timestamp 1688980957
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_489
timestamp 1688980957
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_501
timestamp 1688980957
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_513
timestamp 1688980957
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_525
timestamp 1688980957
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_531
timestamp 1688980957
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_533
timestamp 1688980957
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_545
timestamp 1688980957
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_557
timestamp 1688980957
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_569
timestamp 1688980957
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_581
timestamp 1688980957
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_587
timestamp 1688980957
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_589
timestamp 1688980957
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_601
timestamp 1688980957
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_613
timestamp 1688980957
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_625
timestamp 1688980957
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_637
timestamp 1688980957
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_643
timestamp 1688980957
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_645
timestamp 1688980957
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_657
timestamp 1688980957
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_669
timestamp 1688980957
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_681
timestamp 1688980957
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_693
timestamp 1688980957
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_699
timestamp 1688980957
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_701
timestamp 1688980957
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_713
timestamp 1688980957
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_725
timestamp 1688980957
transform 1 0 67804 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1688980957
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1688980957
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1688980957
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1688980957
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1688980957
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1688980957
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1688980957
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1688980957
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1688980957
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1688980957
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1688980957
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_429
timestamp 1688980957
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_441
timestamp 1688980957
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_447
timestamp 1688980957
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_449
timestamp 1688980957
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_461
timestamp 1688980957
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_473
timestamp 1688980957
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_485
timestamp 1688980957
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_497
timestamp 1688980957
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_503
timestamp 1688980957
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_505
timestamp 1688980957
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_517
timestamp 1688980957
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_529
timestamp 1688980957
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_541
timestamp 1688980957
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_553
timestamp 1688980957
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_559
timestamp 1688980957
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_561
timestamp 1688980957
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_573
timestamp 1688980957
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_585
timestamp 1688980957
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_597
timestamp 1688980957
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_609
timestamp 1688980957
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_615
timestamp 1688980957
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_617
timestamp 1688980957
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_629
timestamp 1688980957
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_641
timestamp 1688980957
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_653
timestamp 1688980957
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_665
timestamp 1688980957
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_671
timestamp 1688980957
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_673
timestamp 1688980957
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_685
timestamp 1688980957
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_697
timestamp 1688980957
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_709
timestamp 1688980957
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_721
timestamp 1688980957
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_727
timestamp 1688980957
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_729
timestamp 1688980957
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_9
timestamp 1688980957
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_21
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1688980957
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1688980957
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 1688980957
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 1688980957
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1688980957
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 1688980957
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 1688980957
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 1688980957
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1688980957
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1688980957
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 1688980957
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1688980957
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 1688980957
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 1688980957
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 1688980957
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 1688980957
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_445
timestamp 1688980957
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_457
timestamp 1688980957
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_469
timestamp 1688980957
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_475
timestamp 1688980957
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_477
timestamp 1688980957
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_489
timestamp 1688980957
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_501
timestamp 1688980957
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_513
timestamp 1688980957
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_525
timestamp 1688980957
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_531
timestamp 1688980957
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_533
timestamp 1688980957
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_545
timestamp 1688980957
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_557
timestamp 1688980957
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_569
timestamp 1688980957
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_581
timestamp 1688980957
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_587
timestamp 1688980957
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_589
timestamp 1688980957
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_601
timestamp 1688980957
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_613
timestamp 1688980957
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_625
timestamp 1688980957
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_637
timestamp 1688980957
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_643
timestamp 1688980957
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_645
timestamp 1688980957
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_657
timestamp 1688980957
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_669
timestamp 1688980957
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_681
timestamp 1688980957
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_693
timestamp 1688980957
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_699
timestamp 1688980957
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_701
timestamp 1688980957
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_713
timestamp 1688980957
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_725
timestamp 1688980957
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1688980957
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 1688980957
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 1688980957
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 1688980957
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_261
timestamp 1688980957
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_273
timestamp 1688980957
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 1688980957
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 1688980957
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 1688980957
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 1688980957
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 1688980957
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 1688980957
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1688980957
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1688980957
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1688980957
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1688980957
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 1688980957
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_429
timestamp 1688980957
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_441
timestamp 1688980957
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_447
timestamp 1688980957
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_449
timestamp 1688980957
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_461
timestamp 1688980957
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_473
timestamp 1688980957
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_485
timestamp 1688980957
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_497
timestamp 1688980957
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_503
timestamp 1688980957
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_505
timestamp 1688980957
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_517
timestamp 1688980957
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_529
timestamp 1688980957
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_541
timestamp 1688980957
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_553
timestamp 1688980957
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_559
timestamp 1688980957
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_561
timestamp 1688980957
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_573
timestamp 1688980957
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_585
timestamp 1688980957
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_597
timestamp 1688980957
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_609
timestamp 1688980957
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_615
timestamp 1688980957
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_617
timestamp 1688980957
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_629
timestamp 1688980957
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_641
timestamp 1688980957
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_653
timestamp 1688980957
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_665
timestamp 1688980957
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_671
timestamp 1688980957
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_673
timestamp 1688980957
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_685
timestamp 1688980957
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_697
timestamp 1688980957
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_709
timestamp 1688980957
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_721
timestamp 1688980957
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_727
timestamp 1688980957
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_729
timestamp 1688980957
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_209
timestamp 1688980957
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_221
timestamp 1688980957
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_233
timestamp 1688980957
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 1688980957
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 1688980957
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 1688980957
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 1688980957
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1688980957
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1688980957
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1688980957
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1688980957
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1688980957
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1688980957
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1688980957
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 1688980957
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 1688980957
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 1688980957
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_433
timestamp 1688980957
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_445
timestamp 1688980957
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_457
timestamp 1688980957
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_469
timestamp 1688980957
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_475
timestamp 1688980957
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_477
timestamp 1688980957
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_489
timestamp 1688980957
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_501
timestamp 1688980957
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_513
timestamp 1688980957
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_525
timestamp 1688980957
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_531
timestamp 1688980957
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_533
timestamp 1688980957
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_545
timestamp 1688980957
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_557
timestamp 1688980957
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_569
timestamp 1688980957
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_581
timestamp 1688980957
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_587
timestamp 1688980957
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_589
timestamp 1688980957
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_601
timestamp 1688980957
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_613
timestamp 1688980957
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_625
timestamp 1688980957
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_637
timestamp 1688980957
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_643
timestamp 1688980957
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_645
timestamp 1688980957
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_657
timestamp 1688980957
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_669
timestamp 1688980957
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_681
timestamp 1688980957
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_693
timestamp 1688980957
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_699
timestamp 1688980957
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_701
timestamp 1688980957
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_713
timestamp 1688980957
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_725
timestamp 1688980957
transform 1 0 67804 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1688980957
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 1688980957
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_237
timestamp 1688980957
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_249
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 1688980957
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 1688980957
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 1688980957
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 1688980957
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 1688980957
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1688980957
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 1688980957
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 1688980957
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 1688980957
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1688980957
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1688980957
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_429
timestamp 1688980957
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_441
timestamp 1688980957
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_447
timestamp 1688980957
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_449
timestamp 1688980957
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_461
timestamp 1688980957
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_473
timestamp 1688980957
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_485
timestamp 1688980957
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_497
timestamp 1688980957
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_503
timestamp 1688980957
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_505
timestamp 1688980957
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_517
timestamp 1688980957
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_529
timestamp 1688980957
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_541
timestamp 1688980957
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_553
timestamp 1688980957
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_559
timestamp 1688980957
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_561
timestamp 1688980957
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_573
timestamp 1688980957
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_585
timestamp 1688980957
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_597
timestamp 1688980957
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_609
timestamp 1688980957
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_615
timestamp 1688980957
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_617
timestamp 1688980957
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_629
timestamp 1688980957
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_641
timestamp 1688980957
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_653
timestamp 1688980957
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_665
timestamp 1688980957
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_671
timestamp 1688980957
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_673
timestamp 1688980957
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_685
timestamp 1688980957
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_697
timestamp 1688980957
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_709
timestamp 1688980957
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_721
timestamp 1688980957
transform 1 0 67436 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_727
timestamp 1688980957
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_729
timestamp 1688980957
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1688980957
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 1688980957
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 1688980957
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 1688980957
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_233
timestamp 1688980957
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_245
timestamp 1688980957
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 1688980957
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 1688980957
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_277
timestamp 1688980957
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 1688980957
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 1688980957
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 1688980957
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 1688980957
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_333
timestamp 1688980957
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 1688980957
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 1688980957
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 1688980957
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1688980957
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1688980957
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1688980957
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1688980957
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 1688980957
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 1688980957
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 1688980957
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_433
timestamp 1688980957
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_445
timestamp 1688980957
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_457
timestamp 1688980957
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_469
timestamp 1688980957
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_475
timestamp 1688980957
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_477
timestamp 1688980957
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_489
timestamp 1688980957
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_501
timestamp 1688980957
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_513
timestamp 1688980957
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_525
timestamp 1688980957
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_531
timestamp 1688980957
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_533
timestamp 1688980957
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_545
timestamp 1688980957
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_557
timestamp 1688980957
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_569
timestamp 1688980957
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_581
timestamp 1688980957
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_587
timestamp 1688980957
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_589
timestamp 1688980957
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_601
timestamp 1688980957
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_613
timestamp 1688980957
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_625
timestamp 1688980957
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_637
timestamp 1688980957
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_643
timestamp 1688980957
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_645
timestamp 1688980957
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_657
timestamp 1688980957
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_669
timestamp 1688980957
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_681
timestamp 1688980957
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_693
timestamp 1688980957
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_699
timestamp 1688980957
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_701
timestamp 1688980957
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_713
timestamp 1688980957
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_725
timestamp 1688980957
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1688980957
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1688980957
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 1688980957
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_205
timestamp 1688980957
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_217
timestamp 1688980957
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 1688980957
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 1688980957
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 1688980957
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 1688980957
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 1688980957
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1688980957
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 1688980957
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 1688980957
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 1688980957
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 1688980957
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 1688980957
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 1688980957
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1688980957
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 1688980957
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 1688980957
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 1688980957
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 1688980957
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 1688980957
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1688980957
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1688980957
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 1688980957
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_429
timestamp 1688980957
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_441
timestamp 1688980957
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_447
timestamp 1688980957
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_449
timestamp 1688980957
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_461
timestamp 1688980957
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_473
timestamp 1688980957
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_485
timestamp 1688980957
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_497
timestamp 1688980957
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_503
timestamp 1688980957
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_505
timestamp 1688980957
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_517
timestamp 1688980957
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_529
timestamp 1688980957
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_541
timestamp 1688980957
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_553
timestamp 1688980957
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_559
timestamp 1688980957
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_561
timestamp 1688980957
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_573
timestamp 1688980957
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_585
timestamp 1688980957
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_597
timestamp 1688980957
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_609
timestamp 1688980957
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_615
timestamp 1688980957
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_617
timestamp 1688980957
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_629
timestamp 1688980957
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_641
timestamp 1688980957
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_653
timestamp 1688980957
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_665
timestamp 1688980957
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_671
timestamp 1688980957
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_673
timestamp 1688980957
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_685
timestamp 1688980957
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_697
timestamp 1688980957
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_709
timestamp 1688980957
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_721
timestamp 1688980957
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_727
timestamp 1688980957
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_729
timestamp 1688980957
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1688980957
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 1688980957
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1688980957
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 1688980957
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 1688980957
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 1688980957
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 1688980957
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 1688980957
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 1688980957
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 1688980957
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 1688980957
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 1688980957
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 1688980957
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1688980957
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1688980957
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1688980957
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1688980957
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 1688980957
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 1688980957
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1688980957
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1688980957
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1688980957
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 1688980957
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 1688980957
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 1688980957
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 1688980957
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_433
timestamp 1688980957
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_445
timestamp 1688980957
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_457
timestamp 1688980957
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_469
timestamp 1688980957
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_475
timestamp 1688980957
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_477
timestamp 1688980957
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_489
timestamp 1688980957
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_501
timestamp 1688980957
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_513
timestamp 1688980957
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_525
timestamp 1688980957
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_531
timestamp 1688980957
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_533
timestamp 1688980957
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_545
timestamp 1688980957
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_557
timestamp 1688980957
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_569
timestamp 1688980957
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_581
timestamp 1688980957
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_587
timestamp 1688980957
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_589
timestamp 1688980957
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_601
timestamp 1688980957
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_613
timestamp 1688980957
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_625
timestamp 1688980957
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_637
timestamp 1688980957
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_643
timestamp 1688980957
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_645
timestamp 1688980957
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_657
timestamp 1688980957
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_669
timestamp 1688980957
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_681
timestamp 1688980957
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_693
timestamp 1688980957
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_699
timestamp 1688980957
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_701
timestamp 1688980957
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_713
timestamp 1688980957
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_725
timestamp 1688980957
transform 1 0 67804 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 1688980957
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 1688980957
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 1688980957
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 1688980957
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 1688980957
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_261
timestamp 1688980957
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 1688980957
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 1688980957
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1688980957
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 1688980957
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 1688980957
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 1688980957
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 1688980957
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 1688980957
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1688980957
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1688980957
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 1688980957
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 1688980957
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 1688980957
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 1688980957
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1688980957
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1688980957
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1688980957
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 1688980957
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_441
timestamp 1688980957
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 1688980957
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_449
timestamp 1688980957
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_461
timestamp 1688980957
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_473
timestamp 1688980957
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_485
timestamp 1688980957
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_497
timestamp 1688980957
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_503
timestamp 1688980957
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_505
timestamp 1688980957
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_517
timestamp 1688980957
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_529
timestamp 1688980957
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_541
timestamp 1688980957
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_553
timestamp 1688980957
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_559
timestamp 1688980957
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_561
timestamp 1688980957
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_573
timestamp 1688980957
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_585
timestamp 1688980957
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_597
timestamp 1688980957
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_609
timestamp 1688980957
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_615
timestamp 1688980957
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_617
timestamp 1688980957
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_629
timestamp 1688980957
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_641
timestamp 1688980957
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_653
timestamp 1688980957
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_665
timestamp 1688980957
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_671
timestamp 1688980957
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_673
timestamp 1688980957
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_685
timestamp 1688980957
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_697
timestamp 1688980957
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_709
timestamp 1688980957
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_721
timestamp 1688980957
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_727
timestamp 1688980957
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_729
timestamp 1688980957
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 1688980957
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1688980957
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 1688980957
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 1688980957
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 1688980957
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 1688980957
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 1688980957
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 1688980957
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 1688980957
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 1688980957
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_301
timestamp 1688980957
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 1688980957
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1688980957
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 1688980957
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 1688980957
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 1688980957
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 1688980957
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 1688980957
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1688980957
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 1688980957
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 1688980957
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 1688980957
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 1688980957
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 1688980957
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 1688980957
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_433
timestamp 1688980957
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_445
timestamp 1688980957
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_457
timestamp 1688980957
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_469
timestamp 1688980957
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_475
timestamp 1688980957
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_477
timestamp 1688980957
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_489
timestamp 1688980957
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_501
timestamp 1688980957
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_513
timestamp 1688980957
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_525
timestamp 1688980957
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_531
timestamp 1688980957
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_533
timestamp 1688980957
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_545
timestamp 1688980957
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_557
timestamp 1688980957
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_569
timestamp 1688980957
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_581
timestamp 1688980957
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_587
timestamp 1688980957
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_589
timestamp 1688980957
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_601
timestamp 1688980957
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_613
timestamp 1688980957
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_625
timestamp 1688980957
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_637
timestamp 1688980957
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_643
timestamp 1688980957
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_645
timestamp 1688980957
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_657
timestamp 1688980957
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_669
timestamp 1688980957
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_681
timestamp 1688980957
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_693
timestamp 1688980957
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_699
timestamp 1688980957
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_701
timestamp 1688980957
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_713
timestamp 1688980957
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_725
timestamp 1688980957
transform 1 0 67804 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1688980957
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_193
timestamp 1688980957
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_205
timestamp 1688980957
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_217
timestamp 1688980957
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1688980957
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 1688980957
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_249
timestamp 1688980957
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_261
timestamp 1688980957
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_273
timestamp 1688980957
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_279
timestamp 1688980957
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 1688980957
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 1688980957
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_305
timestamp 1688980957
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_317
timestamp 1688980957
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_329
timestamp 1688980957
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 1688980957
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_337
timestamp 1688980957
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_349
timestamp 1688980957
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_361
timestamp 1688980957
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_373
timestamp 1688980957
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_385
timestamp 1688980957
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 1688980957
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1688980957
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 1688980957
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 1688980957
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_429
timestamp 1688980957
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_441
timestamp 1688980957
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_447
timestamp 1688980957
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_449
timestamp 1688980957
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_461
timestamp 1688980957
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_473
timestamp 1688980957
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_485
timestamp 1688980957
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_497
timestamp 1688980957
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_503
timestamp 1688980957
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_505
timestamp 1688980957
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_517
timestamp 1688980957
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_529
timestamp 1688980957
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_541
timestamp 1688980957
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_553
timestamp 1688980957
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_559
timestamp 1688980957
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_561
timestamp 1688980957
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_573
timestamp 1688980957
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_585
timestamp 1688980957
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_597
timestamp 1688980957
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_609
timestamp 1688980957
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_615
timestamp 1688980957
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_617
timestamp 1688980957
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_629
timestamp 1688980957
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_641
timestamp 1688980957
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_653
timestamp 1688980957
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_665
timestamp 1688980957
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_671
timestamp 1688980957
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_673
timestamp 1688980957
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_685
timestamp 1688980957
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_697
timestamp 1688980957
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_709
timestamp 1688980957
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_721
timestamp 1688980957
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_727
timestamp 1688980957
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_729
timestamp 1688980957
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1688980957
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1688980957
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1688980957
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 1688980957
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 1688980957
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1688980957
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_197
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_209
timestamp 1688980957
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_221
timestamp 1688980957
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_233
timestamp 1688980957
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_245
timestamp 1688980957
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_251
timestamp 1688980957
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_253
timestamp 1688980957
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_265
timestamp 1688980957
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_277
timestamp 1688980957
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_289
timestamp 1688980957
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_301
timestamp 1688980957
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_307
timestamp 1688980957
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 1688980957
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 1688980957
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 1688980957
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 1688980957
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 1688980957
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 1688980957
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_365
timestamp 1688980957
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_377
timestamp 1688980957
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_389
timestamp 1688980957
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_401
timestamp 1688980957
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_413
timestamp 1688980957
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_419
timestamp 1688980957
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_421
timestamp 1688980957
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_433
timestamp 1688980957
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_445
timestamp 1688980957
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_457
timestamp 1688980957
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_469
timestamp 1688980957
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_475
timestamp 1688980957
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_477
timestamp 1688980957
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_489
timestamp 1688980957
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_501
timestamp 1688980957
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_513
timestamp 1688980957
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_525
timestamp 1688980957
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_531
timestamp 1688980957
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_533
timestamp 1688980957
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_545
timestamp 1688980957
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_557
timestamp 1688980957
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_569
timestamp 1688980957
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_581
timestamp 1688980957
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_587
timestamp 1688980957
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_589
timestamp 1688980957
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_601
timestamp 1688980957
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_613
timestamp 1688980957
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_625
timestamp 1688980957
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_637
timestamp 1688980957
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_643
timestamp 1688980957
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_645
timestamp 1688980957
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_657
timestamp 1688980957
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_669
timestamp 1688980957
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_681
timestamp 1688980957
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_693
timestamp 1688980957
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_699
timestamp 1688980957
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_701
timestamp 1688980957
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_713
timestamp 1688980957
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_725
timestamp 1688980957
transform 1 0 67804 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1688980957
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1688980957
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1688980957
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 1688980957
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1688980957
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 1688980957
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_181
timestamp 1688980957
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_193
timestamp 1688980957
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_205
timestamp 1688980957
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 1688980957
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 1688980957
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 1688980957
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 1688980957
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 1688980957
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 1688980957
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 1688980957
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 1688980957
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_293
timestamp 1688980957
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_305
timestamp 1688980957
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_317
timestamp 1688980957
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 1688980957
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 1688980957
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 1688980957
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_349
timestamp 1688980957
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_361
timestamp 1688980957
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_373
timestamp 1688980957
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_385
timestamp 1688980957
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_391
timestamp 1688980957
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 1688980957
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 1688980957
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 1688980957
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_429
timestamp 1688980957
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_441
timestamp 1688980957
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_447
timestamp 1688980957
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_449
timestamp 1688980957
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_461
timestamp 1688980957
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_473
timestamp 1688980957
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_485
timestamp 1688980957
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_497
timestamp 1688980957
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_503
timestamp 1688980957
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_505
timestamp 1688980957
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_517
timestamp 1688980957
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_529
timestamp 1688980957
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_541
timestamp 1688980957
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_553
timestamp 1688980957
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_559
timestamp 1688980957
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_561
timestamp 1688980957
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_573
timestamp 1688980957
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_585
timestamp 1688980957
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_597
timestamp 1688980957
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_609
timestamp 1688980957
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_615
timestamp 1688980957
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_617
timestamp 1688980957
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_629
timestamp 1688980957
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_641
timestamp 1688980957
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_653
timestamp 1688980957
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_665
timestamp 1688980957
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_671
timestamp 1688980957
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_673
timestamp 1688980957
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_685
timestamp 1688980957
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_697
timestamp 1688980957
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_709
timestamp 1688980957
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_721
timestamp 1688980957
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_727
timestamp 1688980957
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_729
timestamp 1688980957
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1688980957
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1688980957
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1688980957
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 1688980957
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1688980957
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1688980957
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1688980957
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1688980957
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 1688980957
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1688980957
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 1688980957
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 1688980957
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 1688980957
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_189
timestamp 1688980957
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 1688980957
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_197
timestamp 1688980957
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_209
timestamp 1688980957
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_221
timestamp 1688980957
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_233
timestamp 1688980957
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_245
timestamp 1688980957
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 1688980957
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_253
timestamp 1688980957
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_265
timestamp 1688980957
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_277
timestamp 1688980957
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_289
timestamp 1688980957
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_301
timestamp 1688980957
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_307
timestamp 1688980957
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 1688980957
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_321
timestamp 1688980957
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_333
timestamp 1688980957
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_345
timestamp 1688980957
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 1688980957
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 1688980957
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 1688980957
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 1688980957
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 1688980957
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 1688980957
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 1688980957
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 1688980957
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_421
timestamp 1688980957
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_433
timestamp 1688980957
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_445
timestamp 1688980957
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_457
timestamp 1688980957
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_469
timestamp 1688980957
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_475
timestamp 1688980957
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_477
timestamp 1688980957
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_489
timestamp 1688980957
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_501
timestamp 1688980957
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_513
timestamp 1688980957
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_525
timestamp 1688980957
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_531
timestamp 1688980957
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_533
timestamp 1688980957
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_545
timestamp 1688980957
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_557
timestamp 1688980957
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_569
timestamp 1688980957
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_581
timestamp 1688980957
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_587
timestamp 1688980957
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_589
timestamp 1688980957
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_601
timestamp 1688980957
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_613
timestamp 1688980957
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_625
timestamp 1688980957
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_637
timestamp 1688980957
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_643
timestamp 1688980957
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_645
timestamp 1688980957
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_657
timestamp 1688980957
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_669
timestamp 1688980957
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_681
timestamp 1688980957
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_693
timestamp 1688980957
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_699
timestamp 1688980957
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_701
timestamp 1688980957
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_713
timestamp 1688980957
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_725
timestamp 1688980957
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1688980957
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1688980957
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1688980957
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1688980957
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1688980957
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 1688980957
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 1688980957
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1688980957
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 1688980957
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 1688980957
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 1688980957
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 1688980957
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 1688980957
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 1688980957
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_181
timestamp 1688980957
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_193
timestamp 1688980957
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_205
timestamp 1688980957
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_217
timestamp 1688980957
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 1688980957
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 1688980957
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 1688980957
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 1688980957
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 1688980957
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 1688980957
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 1688980957
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 1688980957
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 1688980957
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 1688980957
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 1688980957
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 1688980957
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 1688980957
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 1688980957
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 1688980957
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 1688980957
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 1688980957
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 1688980957
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 1688980957
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 1688980957
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 1688980957
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 1688980957
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_429
timestamp 1688980957
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_441
timestamp 1688980957
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_447
timestamp 1688980957
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_449
timestamp 1688980957
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_461
timestamp 1688980957
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_473
timestamp 1688980957
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_485
timestamp 1688980957
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_497
timestamp 1688980957
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_503
timestamp 1688980957
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_505
timestamp 1688980957
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_517
timestamp 1688980957
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_529
timestamp 1688980957
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_541
timestamp 1688980957
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_553
timestamp 1688980957
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_559
timestamp 1688980957
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_561
timestamp 1688980957
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_573
timestamp 1688980957
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_585
timestamp 1688980957
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_597
timestamp 1688980957
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_609
timestamp 1688980957
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_615
timestamp 1688980957
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_617
timestamp 1688980957
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_629
timestamp 1688980957
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_641
timestamp 1688980957
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_653
timestamp 1688980957
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_665
timestamp 1688980957
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_671
timestamp 1688980957
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_673
timestamp 1688980957
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_685
timestamp 1688980957
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_697
timestamp 1688980957
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_709
timestamp 1688980957
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_721
timestamp 1688980957
transform 1 0 67436 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_727
timestamp 1688980957
transform 1 0 67988 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_729
timestamp 1688980957
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1688980957
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1688980957
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1688980957
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1688980957
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1688980957
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1688980957
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1688980957
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 1688980957
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1688980957
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1688980957
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 1688980957
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 1688980957
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 1688980957
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 1688980957
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 1688980957
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 1688980957
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 1688980957
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 1688980957
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 1688980957
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_189
timestamp 1688980957
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 1688980957
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_197
timestamp 1688980957
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_209
timestamp 1688980957
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_221
timestamp 1688980957
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_233
timestamp 1688980957
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_245
timestamp 1688980957
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_251
timestamp 1688980957
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 1688980957
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 1688980957
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 1688980957
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 1688980957
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 1688980957
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 1688980957
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1688980957
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 1688980957
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_333
timestamp 1688980957
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_345
timestamp 1688980957
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_357
timestamp 1688980957
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_363
timestamp 1688980957
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 1688980957
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 1688980957
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 1688980957
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 1688980957
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 1688980957
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 1688980957
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_421
timestamp 1688980957
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_433
timestamp 1688980957
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_445
timestamp 1688980957
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_457
timestamp 1688980957
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_469
timestamp 1688980957
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_475
timestamp 1688980957
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_477
timestamp 1688980957
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_489
timestamp 1688980957
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_501
timestamp 1688980957
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_513
timestamp 1688980957
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_525
timestamp 1688980957
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_531
timestamp 1688980957
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_533
timestamp 1688980957
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_545
timestamp 1688980957
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_557
timestamp 1688980957
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_569
timestamp 1688980957
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_581
timestamp 1688980957
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_587
timestamp 1688980957
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_589
timestamp 1688980957
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_601
timestamp 1688980957
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_613
timestamp 1688980957
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_625
timestamp 1688980957
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_637
timestamp 1688980957
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_643
timestamp 1688980957
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_645
timestamp 1688980957
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_657
timestamp 1688980957
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_669
timestamp 1688980957
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_681
timestamp 1688980957
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_693
timestamp 1688980957
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_699
timestamp 1688980957
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_701
timestamp 1688980957
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_713
timestamp 1688980957
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_725
timestamp 1688980957
transform 1 0 67804 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1688980957
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1688980957
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 1688980957
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 1688980957
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 1688980957
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 1688980957
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 1688980957
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 1688980957
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_81
timestamp 1688980957
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_93
timestamp 1688980957
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_105
timestamp 1688980957
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_111
timestamp 1688980957
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1688980957
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1688980957
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 1688980957
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 1688980957
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 1688980957
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 1688980957
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 1688980957
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 1688980957
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_193
timestamp 1688980957
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_205
timestamp 1688980957
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_217
timestamp 1688980957
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_223
timestamp 1688980957
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 1688980957
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_237
timestamp 1688980957
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_249
timestamp 1688980957
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_261
timestamp 1688980957
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_273
timestamp 1688980957
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 1688980957
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 1688980957
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 1688980957
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_305
timestamp 1688980957
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_317
timestamp 1688980957
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_329
timestamp 1688980957
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_335
timestamp 1688980957
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 1688980957
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 1688980957
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 1688980957
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 1688980957
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 1688980957
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 1688980957
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 1688980957
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 1688980957
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 1688980957
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_429
timestamp 1688980957
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_441
timestamp 1688980957
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_447
timestamp 1688980957
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_449
timestamp 1688980957
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_461
timestamp 1688980957
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_473
timestamp 1688980957
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_485
timestamp 1688980957
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_497
timestamp 1688980957
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_503
timestamp 1688980957
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_505
timestamp 1688980957
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_517
timestamp 1688980957
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_529
timestamp 1688980957
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_541
timestamp 1688980957
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_553
timestamp 1688980957
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_559
timestamp 1688980957
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_561
timestamp 1688980957
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_573
timestamp 1688980957
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_585
timestamp 1688980957
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_597
timestamp 1688980957
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_609
timestamp 1688980957
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_615
timestamp 1688980957
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_617
timestamp 1688980957
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_629
timestamp 1688980957
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_641
timestamp 1688980957
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_653
timestamp 1688980957
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_665
timestamp 1688980957
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_671
timestamp 1688980957
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_673
timestamp 1688980957
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_685
timestamp 1688980957
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_697
timestamp 1688980957
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_709
timestamp 1688980957
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_721
timestamp 1688980957
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_727
timestamp 1688980957
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_729
timestamp 1688980957
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_3
timestamp 1688980957
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_15
timestamp 1688980957
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 1688980957
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1688980957
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1688980957
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 1688980957
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 1688980957
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 1688980957
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 1688980957
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 1688980957
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1688980957
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 1688980957
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 1688980957
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 1688980957
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 1688980957
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_141
timestamp 1688980957
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 1688980957
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_165
timestamp 1688980957
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_177
timestamp 1688980957
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_189
timestamp 1688980957
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_195
timestamp 1688980957
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 1688980957
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 1688980957
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_221
timestamp 1688980957
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_233
timestamp 1688980957
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_245
timestamp 1688980957
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 1688980957
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 1688980957
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_265
timestamp 1688980957
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_277
timestamp 1688980957
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_289
timestamp 1688980957
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_301
timestamp 1688980957
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 1688980957
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 1688980957
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 1688980957
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_333
timestamp 1688980957
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_345
timestamp 1688980957
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_357
timestamp 1688980957
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_363
timestamp 1688980957
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 1688980957
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 1688980957
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_389
timestamp 1688980957
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_401
timestamp 1688980957
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_413
timestamp 1688980957
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_419
timestamp 1688980957
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_421
timestamp 1688980957
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_433
timestamp 1688980957
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_445
timestamp 1688980957
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_457
timestamp 1688980957
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_469
timestamp 1688980957
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_475
timestamp 1688980957
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_477
timestamp 1688980957
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_489
timestamp 1688980957
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_501
timestamp 1688980957
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_513
timestamp 1688980957
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_525
timestamp 1688980957
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_531
timestamp 1688980957
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_533
timestamp 1688980957
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_545
timestamp 1688980957
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_557
timestamp 1688980957
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_569
timestamp 1688980957
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_581
timestamp 1688980957
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_587
timestamp 1688980957
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_589
timestamp 1688980957
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_601
timestamp 1688980957
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_613
timestamp 1688980957
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_625
timestamp 1688980957
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_637
timestamp 1688980957
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_643
timestamp 1688980957
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_645
timestamp 1688980957
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_657
timestamp 1688980957
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_669
timestamp 1688980957
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_681
timestamp 1688980957
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_693
timestamp 1688980957
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_699
timestamp 1688980957
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_701
timestamp 1688980957
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_713
timestamp 1688980957
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_725
timestamp 1688980957
transform 1 0 67804 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_9
timestamp 1688980957
transform 1 0 1932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_21
timestamp 1688980957
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_33
timestamp 1688980957
transform 1 0 4140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_45
timestamp 1688980957
transform 1 0 5244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81_53
timestamp 1688980957
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 1688980957
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 1688980957
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 1688980957
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 1688980957
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 1688980957
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 1688980957
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 1688980957
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 1688980957
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 1688980957
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 1688980957
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 1688980957
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 1688980957
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 1688980957
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_181
timestamp 1688980957
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_193
timestamp 1688980957
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_205
timestamp 1688980957
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_217
timestamp 1688980957
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_223
timestamp 1688980957
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_225
timestamp 1688980957
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_237
timestamp 1688980957
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_249
timestamp 1688980957
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_261
timestamp 1688980957
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_273
timestamp 1688980957
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_279
timestamp 1688980957
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_281
timestamp 1688980957
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_293
timestamp 1688980957
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_305
timestamp 1688980957
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_317
timestamp 1688980957
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_329
timestamp 1688980957
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_335
timestamp 1688980957
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_337
timestamp 1688980957
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_349
timestamp 1688980957
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_361
timestamp 1688980957
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_373
timestamp 1688980957
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_385
timestamp 1688980957
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_391
timestamp 1688980957
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_393
timestamp 1688980957
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_405
timestamp 1688980957
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_417
timestamp 1688980957
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_429
timestamp 1688980957
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_441
timestamp 1688980957
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_447
timestamp 1688980957
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_449
timestamp 1688980957
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_461
timestamp 1688980957
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_473
timestamp 1688980957
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_485
timestamp 1688980957
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_497
timestamp 1688980957
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_503
timestamp 1688980957
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_505
timestamp 1688980957
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_517
timestamp 1688980957
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_529
timestamp 1688980957
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_541
timestamp 1688980957
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_553
timestamp 1688980957
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_559
timestamp 1688980957
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_561
timestamp 1688980957
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_573
timestamp 1688980957
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_585
timestamp 1688980957
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_597
timestamp 1688980957
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_609
timestamp 1688980957
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_615
timestamp 1688980957
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_617
timestamp 1688980957
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_629
timestamp 1688980957
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_641
timestamp 1688980957
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_653
timestamp 1688980957
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_665
timestamp 1688980957
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_671
timestamp 1688980957
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_673
timestamp 1688980957
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_685
timestamp 1688980957
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_697
timestamp 1688980957
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_709
timestamp 1688980957
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_721
timestamp 1688980957
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_727
timestamp 1688980957
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_729
timestamp 1688980957
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 1688980957
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 1688980957
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 1688980957
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 1688980957
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 1688980957
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_53
timestamp 1688980957
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_65
timestamp 1688980957
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_77
timestamp 1688980957
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 1688980957
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_85
timestamp 1688980957
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_97
timestamp 1688980957
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_109
timestamp 1688980957
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_121
timestamp 1688980957
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_133
timestamp 1688980957
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_139
timestamp 1688980957
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 1688980957
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 1688980957
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_165
timestamp 1688980957
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_177
timestamp 1688980957
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_189
timestamp 1688980957
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_195
timestamp 1688980957
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_197
timestamp 1688980957
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_209
timestamp 1688980957
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_221
timestamp 1688980957
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_233
timestamp 1688980957
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_245
timestamp 1688980957
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_251
timestamp 1688980957
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_253
timestamp 1688980957
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_265
timestamp 1688980957
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_277
timestamp 1688980957
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_289
timestamp 1688980957
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_301
timestamp 1688980957
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_307
timestamp 1688980957
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_309
timestamp 1688980957
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_321
timestamp 1688980957
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_333
timestamp 1688980957
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_345
timestamp 1688980957
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_357
timestamp 1688980957
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_363
timestamp 1688980957
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_365
timestamp 1688980957
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_377
timestamp 1688980957
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_389
timestamp 1688980957
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_401
timestamp 1688980957
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_413
timestamp 1688980957
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_419
timestamp 1688980957
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_421
timestamp 1688980957
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_433
timestamp 1688980957
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_445
timestamp 1688980957
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_457
timestamp 1688980957
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_469
timestamp 1688980957
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_475
timestamp 1688980957
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_477
timestamp 1688980957
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_489
timestamp 1688980957
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_501
timestamp 1688980957
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_513
timestamp 1688980957
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_525
timestamp 1688980957
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_531
timestamp 1688980957
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_533
timestamp 1688980957
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_545
timestamp 1688980957
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_557
timestamp 1688980957
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_569
timestamp 1688980957
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_581
timestamp 1688980957
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_587
timestamp 1688980957
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_589
timestamp 1688980957
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_601
timestamp 1688980957
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_613
timestamp 1688980957
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_625
timestamp 1688980957
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_637
timestamp 1688980957
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_643
timestamp 1688980957
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_645
timestamp 1688980957
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_657
timestamp 1688980957
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_669
timestamp 1688980957
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_681
timestamp 1688980957
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_693
timestamp 1688980957
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_699
timestamp 1688980957
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_701
timestamp 1688980957
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_713
timestamp 1688980957
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_725
timestamp 1688980957
transform 1 0 67804 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_3
timestamp 1688980957
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_15
timestamp 1688980957
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_27
timestamp 1688980957
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_39
timestamp 1688980957
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_51
timestamp 1688980957
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_55
timestamp 1688980957
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_57
timestamp 1688980957
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_69
timestamp 1688980957
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_81
timestamp 1688980957
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_93
timestamp 1688980957
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_105
timestamp 1688980957
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_111
timestamp 1688980957
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_113
timestamp 1688980957
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_125
timestamp 1688980957
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_137
timestamp 1688980957
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_149
timestamp 1688980957
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_161
timestamp 1688980957
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_167
timestamp 1688980957
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_169
timestamp 1688980957
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_181
timestamp 1688980957
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_193
timestamp 1688980957
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_205
timestamp 1688980957
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_217
timestamp 1688980957
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_223
timestamp 1688980957
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_225
timestamp 1688980957
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_237
timestamp 1688980957
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_249
timestamp 1688980957
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_261
timestamp 1688980957
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_273
timestamp 1688980957
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_279
timestamp 1688980957
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_281
timestamp 1688980957
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_293
timestamp 1688980957
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_305
timestamp 1688980957
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_317
timestamp 1688980957
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_329
timestamp 1688980957
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_335
timestamp 1688980957
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_337
timestamp 1688980957
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_349
timestamp 1688980957
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_361
timestamp 1688980957
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_373
timestamp 1688980957
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_385
timestamp 1688980957
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_391
timestamp 1688980957
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_393
timestamp 1688980957
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_405
timestamp 1688980957
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_417
timestamp 1688980957
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_429
timestamp 1688980957
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_441
timestamp 1688980957
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_447
timestamp 1688980957
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_449
timestamp 1688980957
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_461
timestamp 1688980957
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_473
timestamp 1688980957
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_485
timestamp 1688980957
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_497
timestamp 1688980957
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_503
timestamp 1688980957
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_505
timestamp 1688980957
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_517
timestamp 1688980957
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_529
timestamp 1688980957
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_541
timestamp 1688980957
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_553
timestamp 1688980957
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_559
timestamp 1688980957
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_561
timestamp 1688980957
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_573
timestamp 1688980957
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_585
timestamp 1688980957
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_597
timestamp 1688980957
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_609
timestamp 1688980957
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_615
timestamp 1688980957
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_617
timestamp 1688980957
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_629
timestamp 1688980957
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_641
timestamp 1688980957
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_653
timestamp 1688980957
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_665
timestamp 1688980957
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_671
timestamp 1688980957
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_673
timestamp 1688980957
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_685
timestamp 1688980957
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_697
timestamp 1688980957
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_709
timestamp 1688980957
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_721
timestamp 1688980957
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_727
timestamp 1688980957
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_729
timestamp 1688980957
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_3
timestamp 1688980957
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_15
timestamp 1688980957
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 1688980957
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_29
timestamp 1688980957
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_41
timestamp 1688980957
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_53
timestamp 1688980957
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_65
timestamp 1688980957
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 1688980957
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 1688980957
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_85
timestamp 1688980957
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_97
timestamp 1688980957
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_109
timestamp 1688980957
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_121
timestamp 1688980957
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_133
timestamp 1688980957
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_139
timestamp 1688980957
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_141
timestamp 1688980957
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_153
timestamp 1688980957
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_165
timestamp 1688980957
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_177
timestamp 1688980957
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_189
timestamp 1688980957
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_195
timestamp 1688980957
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_197
timestamp 1688980957
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_209
timestamp 1688980957
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_221
timestamp 1688980957
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_233
timestamp 1688980957
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_245
timestamp 1688980957
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_251
timestamp 1688980957
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_253
timestamp 1688980957
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_265
timestamp 1688980957
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_277
timestamp 1688980957
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_289
timestamp 1688980957
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_301
timestamp 1688980957
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_307
timestamp 1688980957
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_309
timestamp 1688980957
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_321
timestamp 1688980957
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_333
timestamp 1688980957
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_345
timestamp 1688980957
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_357
timestamp 1688980957
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_363
timestamp 1688980957
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_365
timestamp 1688980957
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_377
timestamp 1688980957
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_389
timestamp 1688980957
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_401
timestamp 1688980957
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_413
timestamp 1688980957
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_419
timestamp 1688980957
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_421
timestamp 1688980957
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_433
timestamp 1688980957
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_445
timestamp 1688980957
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_457
timestamp 1688980957
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_469
timestamp 1688980957
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_475
timestamp 1688980957
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_477
timestamp 1688980957
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_489
timestamp 1688980957
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_501
timestamp 1688980957
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_513
timestamp 1688980957
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_525
timestamp 1688980957
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_531
timestamp 1688980957
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_533
timestamp 1688980957
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_545
timestamp 1688980957
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_557
timestamp 1688980957
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_569
timestamp 1688980957
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_581
timestamp 1688980957
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_587
timestamp 1688980957
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_589
timestamp 1688980957
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_601
timestamp 1688980957
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_613
timestamp 1688980957
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_625
timestamp 1688980957
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_637
timestamp 1688980957
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_643
timestamp 1688980957
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_645
timestamp 1688980957
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_657
timestamp 1688980957
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_669
timestamp 1688980957
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_681
timestamp 1688980957
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_693
timestamp 1688980957
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_699
timestamp 1688980957
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_701
timestamp 1688980957
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_713
timestamp 1688980957
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_725
timestamp 1688980957
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_3
timestamp 1688980957
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_15
timestamp 1688980957
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_27
timestamp 1688980957
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_39
timestamp 1688980957
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_51
timestamp 1688980957
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_55
timestamp 1688980957
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_57
timestamp 1688980957
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 1688980957
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 1688980957
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_93
timestamp 1688980957
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_105
timestamp 1688980957
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_111
timestamp 1688980957
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_113
timestamp 1688980957
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_125
timestamp 1688980957
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_137
timestamp 1688980957
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_149
timestamp 1688980957
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_161
timestamp 1688980957
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_167
timestamp 1688980957
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_169
timestamp 1688980957
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_181
timestamp 1688980957
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_193
timestamp 1688980957
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_205
timestamp 1688980957
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_217
timestamp 1688980957
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_223
timestamp 1688980957
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_225
timestamp 1688980957
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_237
timestamp 1688980957
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_249
timestamp 1688980957
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_261
timestamp 1688980957
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_273
timestamp 1688980957
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_279
timestamp 1688980957
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_281
timestamp 1688980957
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_293
timestamp 1688980957
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_305
timestamp 1688980957
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_317
timestamp 1688980957
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_329
timestamp 1688980957
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_335
timestamp 1688980957
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_337
timestamp 1688980957
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_349
timestamp 1688980957
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_361
timestamp 1688980957
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_373
timestamp 1688980957
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_385
timestamp 1688980957
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_391
timestamp 1688980957
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_393
timestamp 1688980957
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_405
timestamp 1688980957
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_417
timestamp 1688980957
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_429
timestamp 1688980957
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_441
timestamp 1688980957
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_447
timestamp 1688980957
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_449
timestamp 1688980957
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_461
timestamp 1688980957
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_473
timestamp 1688980957
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_485
timestamp 1688980957
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_497
timestamp 1688980957
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_503
timestamp 1688980957
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_505
timestamp 1688980957
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_517
timestamp 1688980957
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_529
timestamp 1688980957
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_541
timestamp 1688980957
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_553
timestamp 1688980957
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_559
timestamp 1688980957
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_561
timestamp 1688980957
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_573
timestamp 1688980957
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_585
timestamp 1688980957
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_597
timestamp 1688980957
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_609
timestamp 1688980957
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_615
timestamp 1688980957
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_617
timestamp 1688980957
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_629
timestamp 1688980957
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_641
timestamp 1688980957
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_653
timestamp 1688980957
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_665
timestamp 1688980957
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_671
timestamp 1688980957
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_673
timestamp 1688980957
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_685
timestamp 1688980957
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_697
timestamp 1688980957
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_709
timestamp 1688980957
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_721
timestamp 1688980957
transform 1 0 67436 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_727
timestamp 1688980957
transform 1 0 67988 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_729
timestamp 1688980957
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_3
timestamp 1688980957
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_15
timestamp 1688980957
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 1688980957
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 1688980957
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 1688980957
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_53
timestamp 1688980957
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_65
timestamp 1688980957
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_77
timestamp 1688980957
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_83
timestamp 1688980957
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_85
timestamp 1688980957
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_97
timestamp 1688980957
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_109
timestamp 1688980957
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_121
timestamp 1688980957
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_133
timestamp 1688980957
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_139
timestamp 1688980957
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_141
timestamp 1688980957
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_153
timestamp 1688980957
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_165
timestamp 1688980957
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_177
timestamp 1688980957
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_189
timestamp 1688980957
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_195
timestamp 1688980957
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_197
timestamp 1688980957
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_209
timestamp 1688980957
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_221
timestamp 1688980957
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_233
timestamp 1688980957
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_245
timestamp 1688980957
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_251
timestamp 1688980957
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_253
timestamp 1688980957
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_265
timestamp 1688980957
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_277
timestamp 1688980957
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_289
timestamp 1688980957
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_301
timestamp 1688980957
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_307
timestamp 1688980957
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_309
timestamp 1688980957
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_321
timestamp 1688980957
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_333
timestamp 1688980957
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_345
timestamp 1688980957
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_357
timestamp 1688980957
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_363
timestamp 1688980957
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_365
timestamp 1688980957
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_377
timestamp 1688980957
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_389
timestamp 1688980957
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_401
timestamp 1688980957
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_413
timestamp 1688980957
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_419
timestamp 1688980957
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_421
timestamp 1688980957
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_433
timestamp 1688980957
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_445
timestamp 1688980957
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_457
timestamp 1688980957
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_469
timestamp 1688980957
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_475
timestamp 1688980957
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_477
timestamp 1688980957
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_489
timestamp 1688980957
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_501
timestamp 1688980957
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_513
timestamp 1688980957
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_525
timestamp 1688980957
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_531
timestamp 1688980957
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_533
timestamp 1688980957
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_545
timestamp 1688980957
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_557
timestamp 1688980957
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_569
timestamp 1688980957
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_581
timestamp 1688980957
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_587
timestamp 1688980957
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_589
timestamp 1688980957
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_601
timestamp 1688980957
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_613
timestamp 1688980957
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_625
timestamp 1688980957
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_637
timestamp 1688980957
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_643
timestamp 1688980957
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_645
timestamp 1688980957
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_657
timestamp 1688980957
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_669
timestamp 1688980957
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_681
timestamp 1688980957
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_693
timestamp 1688980957
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_699
timestamp 1688980957
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_701
timestamp 1688980957
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_713
timestamp 1688980957
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_725
timestamp 1688980957
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_3
timestamp 1688980957
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_15
timestamp 1688980957
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_27
timestamp 1688980957
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_39
timestamp 1688980957
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_51
timestamp 1688980957
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_55
timestamp 1688980957
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_57
timestamp 1688980957
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_69
timestamp 1688980957
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_81
timestamp 1688980957
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_93
timestamp 1688980957
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_105
timestamp 1688980957
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_111
timestamp 1688980957
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_113
timestamp 1688980957
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_125
timestamp 1688980957
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_137
timestamp 1688980957
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_149
timestamp 1688980957
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_161
timestamp 1688980957
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_167
timestamp 1688980957
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_169
timestamp 1688980957
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_181
timestamp 1688980957
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_193
timestamp 1688980957
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_205
timestamp 1688980957
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_217
timestamp 1688980957
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_223
timestamp 1688980957
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_225
timestamp 1688980957
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_237
timestamp 1688980957
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_249
timestamp 1688980957
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_261
timestamp 1688980957
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_273
timestamp 1688980957
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_279
timestamp 1688980957
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_281
timestamp 1688980957
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_293
timestamp 1688980957
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_305
timestamp 1688980957
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_317
timestamp 1688980957
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_329
timestamp 1688980957
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_335
timestamp 1688980957
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_337
timestamp 1688980957
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_349
timestamp 1688980957
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_361
timestamp 1688980957
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_373
timestamp 1688980957
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_385
timestamp 1688980957
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_391
timestamp 1688980957
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_393
timestamp 1688980957
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_405
timestamp 1688980957
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_417
timestamp 1688980957
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_429
timestamp 1688980957
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_441
timestamp 1688980957
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_447
timestamp 1688980957
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_449
timestamp 1688980957
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_461
timestamp 1688980957
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_473
timestamp 1688980957
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_485
timestamp 1688980957
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_497
timestamp 1688980957
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_503
timestamp 1688980957
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_505
timestamp 1688980957
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_517
timestamp 1688980957
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_529
timestamp 1688980957
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_541
timestamp 1688980957
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_553
timestamp 1688980957
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_559
timestamp 1688980957
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_561
timestamp 1688980957
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_573
timestamp 1688980957
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_585
timestamp 1688980957
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_597
timestamp 1688980957
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_609
timestamp 1688980957
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_615
timestamp 1688980957
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_617
timestamp 1688980957
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_629
timestamp 1688980957
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_641
timestamp 1688980957
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_653
timestamp 1688980957
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_665
timestamp 1688980957
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_671
timestamp 1688980957
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_673
timestamp 1688980957
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_685
timestamp 1688980957
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_697
timestamp 1688980957
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_709
timestamp 1688980957
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_721
timestamp 1688980957
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_727
timestamp 1688980957
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_729
timestamp 1688980957
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_3
timestamp 1688980957
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_15
timestamp 1688980957
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 1688980957
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 1688980957
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 1688980957
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_53
timestamp 1688980957
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_65
timestamp 1688980957
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_77
timestamp 1688980957
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 1688980957
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_85
timestamp 1688980957
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_97
timestamp 1688980957
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_109
timestamp 1688980957
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_121
timestamp 1688980957
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_133
timestamp 1688980957
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_139
timestamp 1688980957
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_141
timestamp 1688980957
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_153
timestamp 1688980957
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_165
timestamp 1688980957
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_177
timestamp 1688980957
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_189
timestamp 1688980957
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_195
timestamp 1688980957
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_197
timestamp 1688980957
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_209
timestamp 1688980957
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_221
timestamp 1688980957
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_233
timestamp 1688980957
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_245
timestamp 1688980957
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_251
timestamp 1688980957
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_253
timestamp 1688980957
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_265
timestamp 1688980957
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_277
timestamp 1688980957
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_289
timestamp 1688980957
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_301
timestamp 1688980957
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_307
timestamp 1688980957
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_309
timestamp 1688980957
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_321
timestamp 1688980957
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_333
timestamp 1688980957
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_345
timestamp 1688980957
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_357
timestamp 1688980957
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_363
timestamp 1688980957
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_365
timestamp 1688980957
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_377
timestamp 1688980957
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_389
timestamp 1688980957
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_401
timestamp 1688980957
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_413
timestamp 1688980957
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_419
timestamp 1688980957
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_421
timestamp 1688980957
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_433
timestamp 1688980957
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_445
timestamp 1688980957
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_457
timestamp 1688980957
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_469
timestamp 1688980957
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_475
timestamp 1688980957
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_477
timestamp 1688980957
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_489
timestamp 1688980957
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_501
timestamp 1688980957
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_513
timestamp 1688980957
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_525
timestamp 1688980957
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_531
timestamp 1688980957
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_533
timestamp 1688980957
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_545
timestamp 1688980957
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_557
timestamp 1688980957
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_569
timestamp 1688980957
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_581
timestamp 1688980957
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_587
timestamp 1688980957
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_589
timestamp 1688980957
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_601
timestamp 1688980957
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_613
timestamp 1688980957
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_625
timestamp 1688980957
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_637
timestamp 1688980957
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_643
timestamp 1688980957
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_645
timestamp 1688980957
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_657
timestamp 1688980957
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_669
timestamp 1688980957
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_681
timestamp 1688980957
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_693
timestamp 1688980957
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_699
timestamp 1688980957
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_701
timestamp 1688980957
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_713
timestamp 1688980957
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_725
timestamp 1688980957
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_3
timestamp 1688980957
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_15
timestamp 1688980957
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_27
timestamp 1688980957
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_39
timestamp 1688980957
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_51
timestamp 1688980957
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 1688980957
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_57
timestamp 1688980957
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_69
timestamp 1688980957
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_81
timestamp 1688980957
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_93
timestamp 1688980957
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_105
timestamp 1688980957
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_111
timestamp 1688980957
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_113
timestamp 1688980957
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_125
timestamp 1688980957
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_137
timestamp 1688980957
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_149
timestamp 1688980957
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_161
timestamp 1688980957
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_167
timestamp 1688980957
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_169
timestamp 1688980957
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_181
timestamp 1688980957
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_193
timestamp 1688980957
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_205
timestamp 1688980957
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_217
timestamp 1688980957
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_223
timestamp 1688980957
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_225
timestamp 1688980957
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_237
timestamp 1688980957
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_249
timestamp 1688980957
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_261
timestamp 1688980957
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_273
timestamp 1688980957
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_279
timestamp 1688980957
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_281
timestamp 1688980957
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_293
timestamp 1688980957
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_305
timestamp 1688980957
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_317
timestamp 1688980957
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_329
timestamp 1688980957
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_335
timestamp 1688980957
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_337
timestamp 1688980957
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_349
timestamp 1688980957
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_361
timestamp 1688980957
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_373
timestamp 1688980957
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_385
timestamp 1688980957
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_391
timestamp 1688980957
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_393
timestamp 1688980957
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_405
timestamp 1688980957
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_417
timestamp 1688980957
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_429
timestamp 1688980957
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_441
timestamp 1688980957
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_447
timestamp 1688980957
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_449
timestamp 1688980957
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_461
timestamp 1688980957
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_473
timestamp 1688980957
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_485
timestamp 1688980957
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_497
timestamp 1688980957
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_503
timestamp 1688980957
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_505
timestamp 1688980957
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_517
timestamp 1688980957
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_529
timestamp 1688980957
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_541
timestamp 1688980957
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_553
timestamp 1688980957
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_559
timestamp 1688980957
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_561
timestamp 1688980957
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_573
timestamp 1688980957
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_585
timestamp 1688980957
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_597
timestamp 1688980957
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_609
timestamp 1688980957
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_615
timestamp 1688980957
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_617
timestamp 1688980957
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_629
timestamp 1688980957
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_641
timestamp 1688980957
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_653
timestamp 1688980957
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_665
timestamp 1688980957
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_671
timestamp 1688980957
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_673
timestamp 1688980957
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_685
timestamp 1688980957
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_697
timestamp 1688980957
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_709
timestamp 1688980957
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_721
timestamp 1688980957
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_727
timestamp 1688980957
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_729
timestamp 1688980957
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_3
timestamp 1688980957
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_15
timestamp 1688980957
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 1688980957
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 1688980957
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 1688980957
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 1688980957
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 1688980957
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 1688980957
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 1688980957
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_85
timestamp 1688980957
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_97
timestamp 1688980957
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_109
timestamp 1688980957
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_121
timestamp 1688980957
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_133
timestamp 1688980957
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_139
timestamp 1688980957
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_141
timestamp 1688980957
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_153
timestamp 1688980957
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_165
timestamp 1688980957
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_177
timestamp 1688980957
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_189
timestamp 1688980957
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_195
timestamp 1688980957
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_197
timestamp 1688980957
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_209
timestamp 1688980957
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_221
timestamp 1688980957
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_233
timestamp 1688980957
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_245
timestamp 1688980957
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_251
timestamp 1688980957
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_253
timestamp 1688980957
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_265
timestamp 1688980957
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_277
timestamp 1688980957
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_289
timestamp 1688980957
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_301
timestamp 1688980957
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_307
timestamp 1688980957
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_309
timestamp 1688980957
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_321
timestamp 1688980957
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_333
timestamp 1688980957
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_345
timestamp 1688980957
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_357
timestamp 1688980957
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_363
timestamp 1688980957
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_365
timestamp 1688980957
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_377
timestamp 1688980957
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_389
timestamp 1688980957
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_401
timestamp 1688980957
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_413
timestamp 1688980957
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_419
timestamp 1688980957
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_421
timestamp 1688980957
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_433
timestamp 1688980957
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_445
timestamp 1688980957
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_457
timestamp 1688980957
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_469
timestamp 1688980957
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_475
timestamp 1688980957
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_477
timestamp 1688980957
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_489
timestamp 1688980957
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_501
timestamp 1688980957
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_513
timestamp 1688980957
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_525
timestamp 1688980957
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_531
timestamp 1688980957
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_533
timestamp 1688980957
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_545
timestamp 1688980957
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_557
timestamp 1688980957
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_569
timestamp 1688980957
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_581
timestamp 1688980957
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_587
timestamp 1688980957
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_589
timestamp 1688980957
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_601
timestamp 1688980957
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_613
timestamp 1688980957
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_625
timestamp 1688980957
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_637
timestamp 1688980957
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_643
timestamp 1688980957
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_645
timestamp 1688980957
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_657
timestamp 1688980957
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_669
timestamp 1688980957
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_681
timestamp 1688980957
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_693
timestamp 1688980957
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_699
timestamp 1688980957
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_701
timestamp 1688980957
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_713
timestamp 1688980957
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_725
timestamp 1688980957
transform 1 0 67804 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 1688980957
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 1688980957
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_27
timestamp 1688980957
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_39
timestamp 1688980957
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_51
timestamp 1688980957
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_55
timestamp 1688980957
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_57
timestamp 1688980957
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_69
timestamp 1688980957
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_81
timestamp 1688980957
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_93
timestamp 1688980957
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_105
timestamp 1688980957
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_111
timestamp 1688980957
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_113
timestamp 1688980957
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_125
timestamp 1688980957
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_137
timestamp 1688980957
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_149
timestamp 1688980957
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_161
timestamp 1688980957
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_167
timestamp 1688980957
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_169
timestamp 1688980957
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_181
timestamp 1688980957
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_193
timestamp 1688980957
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_205
timestamp 1688980957
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_217
timestamp 1688980957
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_223
timestamp 1688980957
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_225
timestamp 1688980957
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_237
timestamp 1688980957
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_249
timestamp 1688980957
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_261
timestamp 1688980957
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_273
timestamp 1688980957
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_279
timestamp 1688980957
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_281
timestamp 1688980957
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_293
timestamp 1688980957
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_305
timestamp 1688980957
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_317
timestamp 1688980957
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_329
timestamp 1688980957
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_335
timestamp 1688980957
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_337
timestamp 1688980957
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_349
timestamp 1688980957
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_361
timestamp 1688980957
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_373
timestamp 1688980957
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_385
timestamp 1688980957
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_391
timestamp 1688980957
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_393
timestamp 1688980957
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_405
timestamp 1688980957
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_417
timestamp 1688980957
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_429
timestamp 1688980957
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_441
timestamp 1688980957
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_447
timestamp 1688980957
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_449
timestamp 1688980957
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_461
timestamp 1688980957
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_473
timestamp 1688980957
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_485
timestamp 1688980957
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_497
timestamp 1688980957
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_503
timestamp 1688980957
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_505
timestamp 1688980957
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_517
timestamp 1688980957
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_529
timestamp 1688980957
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_541
timestamp 1688980957
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_553
timestamp 1688980957
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_559
timestamp 1688980957
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_561
timestamp 1688980957
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_573
timestamp 1688980957
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_585
timestamp 1688980957
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_597
timestamp 1688980957
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_609
timestamp 1688980957
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_615
timestamp 1688980957
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_617
timestamp 1688980957
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_629
timestamp 1688980957
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_641
timestamp 1688980957
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_653
timestamp 1688980957
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_665
timestamp 1688980957
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_671
timestamp 1688980957
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_673
timestamp 1688980957
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_685
timestamp 1688980957
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_697
timestamp 1688980957
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_709
timestamp 1688980957
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_721
timestamp 1688980957
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_727
timestamp 1688980957
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_729
timestamp 1688980957
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_3
timestamp 1688980957
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_15
timestamp 1688980957
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 1688980957
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_29
timestamp 1688980957
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_41
timestamp 1688980957
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_53
timestamp 1688980957
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_65
timestamp 1688980957
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_77
timestamp 1688980957
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_83
timestamp 1688980957
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_85
timestamp 1688980957
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_97
timestamp 1688980957
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_109
timestamp 1688980957
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_121
timestamp 1688980957
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_133
timestamp 1688980957
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_139
timestamp 1688980957
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_141
timestamp 1688980957
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_153
timestamp 1688980957
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_165
timestamp 1688980957
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_177
timestamp 1688980957
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_189
timestamp 1688980957
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_195
timestamp 1688980957
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_197
timestamp 1688980957
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_209
timestamp 1688980957
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_221
timestamp 1688980957
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_233
timestamp 1688980957
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_245
timestamp 1688980957
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_251
timestamp 1688980957
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_253
timestamp 1688980957
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_265
timestamp 1688980957
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_277
timestamp 1688980957
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_289
timestamp 1688980957
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_301
timestamp 1688980957
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_307
timestamp 1688980957
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_309
timestamp 1688980957
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_321
timestamp 1688980957
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_333
timestamp 1688980957
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_345
timestamp 1688980957
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_357
timestamp 1688980957
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_363
timestamp 1688980957
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_365
timestamp 1688980957
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_377
timestamp 1688980957
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_389
timestamp 1688980957
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_401
timestamp 1688980957
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_413
timestamp 1688980957
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_419
timestamp 1688980957
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_421
timestamp 1688980957
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_433
timestamp 1688980957
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_445
timestamp 1688980957
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_457
timestamp 1688980957
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_469
timestamp 1688980957
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_475
timestamp 1688980957
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_477
timestamp 1688980957
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_489
timestamp 1688980957
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_501
timestamp 1688980957
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_513
timestamp 1688980957
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_525
timestamp 1688980957
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_531
timestamp 1688980957
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_533
timestamp 1688980957
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_545
timestamp 1688980957
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_557
timestamp 1688980957
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_569
timestamp 1688980957
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_581
timestamp 1688980957
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_587
timestamp 1688980957
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_589
timestamp 1688980957
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_601
timestamp 1688980957
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_613
timestamp 1688980957
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_625
timestamp 1688980957
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_637
timestamp 1688980957
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_643
timestamp 1688980957
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_645
timestamp 1688980957
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_657
timestamp 1688980957
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_669
timestamp 1688980957
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_681
timestamp 1688980957
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_693
timestamp 1688980957
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_699
timestamp 1688980957
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_701
timestamp 1688980957
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_713
timestamp 1688980957
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_725
timestamp 1688980957
transform 1 0 67804 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 1688980957
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 1688980957
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_27
timestamp 1688980957
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_39
timestamp 1688980957
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_51
timestamp 1688980957
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_55
timestamp 1688980957
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_57
timestamp 1688980957
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_69
timestamp 1688980957
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_81
timestamp 1688980957
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_93
timestamp 1688980957
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_105
timestamp 1688980957
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_111
timestamp 1688980957
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_113
timestamp 1688980957
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_125
timestamp 1688980957
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_137
timestamp 1688980957
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_149
timestamp 1688980957
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_161
timestamp 1688980957
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_167
timestamp 1688980957
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_169
timestamp 1688980957
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_181
timestamp 1688980957
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_193
timestamp 1688980957
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_205
timestamp 1688980957
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_217
timestamp 1688980957
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_223
timestamp 1688980957
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_225
timestamp 1688980957
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_237
timestamp 1688980957
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_249
timestamp 1688980957
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_261
timestamp 1688980957
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_273
timestamp 1688980957
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_279
timestamp 1688980957
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_281
timestamp 1688980957
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_293
timestamp 1688980957
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_305
timestamp 1688980957
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_317
timestamp 1688980957
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_329
timestamp 1688980957
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_335
timestamp 1688980957
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_337
timestamp 1688980957
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_349
timestamp 1688980957
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_361
timestamp 1688980957
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_373
timestamp 1688980957
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_385
timestamp 1688980957
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_391
timestamp 1688980957
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_393
timestamp 1688980957
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_405
timestamp 1688980957
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_417
timestamp 1688980957
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_429
timestamp 1688980957
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_441
timestamp 1688980957
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_447
timestamp 1688980957
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_449
timestamp 1688980957
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_461
timestamp 1688980957
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_473
timestamp 1688980957
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_485
timestamp 1688980957
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_497
timestamp 1688980957
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_503
timestamp 1688980957
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_505
timestamp 1688980957
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_517
timestamp 1688980957
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_529
timestamp 1688980957
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_541
timestamp 1688980957
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_553
timestamp 1688980957
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_559
timestamp 1688980957
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_561
timestamp 1688980957
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_573
timestamp 1688980957
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_585
timestamp 1688980957
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_597
timestamp 1688980957
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_609
timestamp 1688980957
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_615
timestamp 1688980957
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_617
timestamp 1688980957
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_629
timestamp 1688980957
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_641
timestamp 1688980957
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_653
timestamp 1688980957
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_665
timestamp 1688980957
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_671
timestamp 1688980957
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_673
timestamp 1688980957
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_685
timestamp 1688980957
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_697
timestamp 1688980957
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_709
timestamp 1688980957
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_721
timestamp 1688980957
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_727
timestamp 1688980957
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_729
timestamp 1688980957
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_3
timestamp 1688980957
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_15
timestamp 1688980957
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 1688980957
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_29
timestamp 1688980957
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_41
timestamp 1688980957
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_53
timestamp 1688980957
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_65
timestamp 1688980957
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_77
timestamp 1688980957
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_83
timestamp 1688980957
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_85
timestamp 1688980957
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_97
timestamp 1688980957
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_109
timestamp 1688980957
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_121
timestamp 1688980957
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_133
timestamp 1688980957
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_139
timestamp 1688980957
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_141
timestamp 1688980957
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_153
timestamp 1688980957
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_165
timestamp 1688980957
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_177
timestamp 1688980957
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_189
timestamp 1688980957
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_195
timestamp 1688980957
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_197
timestamp 1688980957
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_209
timestamp 1688980957
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_221
timestamp 1688980957
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_233
timestamp 1688980957
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_245
timestamp 1688980957
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_251
timestamp 1688980957
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_253
timestamp 1688980957
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_265
timestamp 1688980957
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_277
timestamp 1688980957
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_289
timestamp 1688980957
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_301
timestamp 1688980957
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_307
timestamp 1688980957
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_309
timestamp 1688980957
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_321
timestamp 1688980957
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_333
timestamp 1688980957
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_345
timestamp 1688980957
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_357
timestamp 1688980957
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_363
timestamp 1688980957
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_365
timestamp 1688980957
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_377
timestamp 1688980957
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_389
timestamp 1688980957
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_401
timestamp 1688980957
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_413
timestamp 1688980957
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_419
timestamp 1688980957
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_421
timestamp 1688980957
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_433
timestamp 1688980957
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_445
timestamp 1688980957
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_457
timestamp 1688980957
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_469
timestamp 1688980957
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_475
timestamp 1688980957
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_477
timestamp 1688980957
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_489
timestamp 1688980957
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_501
timestamp 1688980957
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_513
timestamp 1688980957
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_525
timestamp 1688980957
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_531
timestamp 1688980957
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_533
timestamp 1688980957
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_545
timestamp 1688980957
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_557
timestamp 1688980957
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_569
timestamp 1688980957
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_581
timestamp 1688980957
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_587
timestamp 1688980957
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_589
timestamp 1688980957
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_601
timestamp 1688980957
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_613
timestamp 1688980957
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_625
timestamp 1688980957
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_637
timestamp 1688980957
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_643
timestamp 1688980957
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_645
timestamp 1688980957
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_657
timestamp 1688980957
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_669
timestamp 1688980957
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_681
timestamp 1688980957
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_693
timestamp 1688980957
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_699
timestamp 1688980957
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_701
timestamp 1688980957
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_713
timestamp 1688980957
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_725
timestamp 1688980957
transform 1 0 67804 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_3
timestamp 1688980957
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_15
timestamp 1688980957
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_27
timestamp 1688980957
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_39
timestamp 1688980957
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_51
timestamp 1688980957
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_55
timestamp 1688980957
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_57
timestamp 1688980957
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_69
timestamp 1688980957
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_81
timestamp 1688980957
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_93
timestamp 1688980957
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_105
timestamp 1688980957
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_111
timestamp 1688980957
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_113
timestamp 1688980957
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_125
timestamp 1688980957
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_137
timestamp 1688980957
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_149
timestamp 1688980957
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_161
timestamp 1688980957
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_167
timestamp 1688980957
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_169
timestamp 1688980957
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_181
timestamp 1688980957
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_193
timestamp 1688980957
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_205
timestamp 1688980957
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_217
timestamp 1688980957
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_223
timestamp 1688980957
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_225
timestamp 1688980957
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_237
timestamp 1688980957
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_249
timestamp 1688980957
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_261
timestamp 1688980957
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_273
timestamp 1688980957
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_279
timestamp 1688980957
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_281
timestamp 1688980957
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_293
timestamp 1688980957
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_305
timestamp 1688980957
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_317
timestamp 1688980957
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_329
timestamp 1688980957
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_335
timestamp 1688980957
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_337
timestamp 1688980957
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_349
timestamp 1688980957
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_361
timestamp 1688980957
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_373
timestamp 1688980957
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_385
timestamp 1688980957
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_391
timestamp 1688980957
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_393
timestamp 1688980957
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_405
timestamp 1688980957
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_417
timestamp 1688980957
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_429
timestamp 1688980957
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_441
timestamp 1688980957
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_447
timestamp 1688980957
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_449
timestamp 1688980957
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_461
timestamp 1688980957
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_473
timestamp 1688980957
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_485
timestamp 1688980957
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_497
timestamp 1688980957
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_503
timestamp 1688980957
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_505
timestamp 1688980957
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_517
timestamp 1688980957
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_529
timestamp 1688980957
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_541
timestamp 1688980957
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_553
timestamp 1688980957
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_559
timestamp 1688980957
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_561
timestamp 1688980957
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_573
timestamp 1688980957
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_585
timestamp 1688980957
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_597
timestamp 1688980957
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_609
timestamp 1688980957
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_615
timestamp 1688980957
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_617
timestamp 1688980957
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_629
timestamp 1688980957
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_641
timestamp 1688980957
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_653
timestamp 1688980957
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_665
timestamp 1688980957
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_671
timestamp 1688980957
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_673
timestamp 1688980957
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_685
timestamp 1688980957
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_697
timestamp 1688980957
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_709
timestamp 1688980957
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_721
timestamp 1688980957
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_727
timestamp 1688980957
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_729
timestamp 1688980957
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 1688980957
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 1688980957
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 1688980957
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_29
timestamp 1688980957
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_41
timestamp 1688980957
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_53
timestamp 1688980957
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_65
timestamp 1688980957
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_77
timestamp 1688980957
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 1688980957
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_85
timestamp 1688980957
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_97
timestamp 1688980957
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_109
timestamp 1688980957
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_121
timestamp 1688980957
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_133
timestamp 1688980957
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_139
timestamp 1688980957
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_141
timestamp 1688980957
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_153
timestamp 1688980957
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_165
timestamp 1688980957
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_177
timestamp 1688980957
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_189
timestamp 1688980957
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_195
timestamp 1688980957
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_197
timestamp 1688980957
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_209
timestamp 1688980957
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_221
timestamp 1688980957
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_233
timestamp 1688980957
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_245
timestamp 1688980957
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_251
timestamp 1688980957
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_253
timestamp 1688980957
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_265
timestamp 1688980957
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_277
timestamp 1688980957
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_289
timestamp 1688980957
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_301
timestamp 1688980957
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_307
timestamp 1688980957
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_309
timestamp 1688980957
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_321
timestamp 1688980957
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_333
timestamp 1688980957
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_345
timestamp 1688980957
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_357
timestamp 1688980957
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_363
timestamp 1688980957
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_365
timestamp 1688980957
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_377
timestamp 1688980957
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_389
timestamp 1688980957
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_401
timestamp 1688980957
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_413
timestamp 1688980957
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_419
timestamp 1688980957
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_421
timestamp 1688980957
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_433
timestamp 1688980957
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_445
timestamp 1688980957
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_457
timestamp 1688980957
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_469
timestamp 1688980957
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_475
timestamp 1688980957
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_477
timestamp 1688980957
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_489
timestamp 1688980957
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_501
timestamp 1688980957
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_513
timestamp 1688980957
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_525
timestamp 1688980957
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_531
timestamp 1688980957
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_533
timestamp 1688980957
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_545
timestamp 1688980957
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_557
timestamp 1688980957
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_569
timestamp 1688980957
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_581
timestamp 1688980957
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_587
timestamp 1688980957
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_589
timestamp 1688980957
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_601
timestamp 1688980957
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_613
timestamp 1688980957
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_625
timestamp 1688980957
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_637
timestamp 1688980957
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_643
timestamp 1688980957
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_645
timestamp 1688980957
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_657
timestamp 1688980957
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_669
timestamp 1688980957
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_681
timestamp 1688980957
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_693
timestamp 1688980957
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_699
timestamp 1688980957
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_701
timestamp 1688980957
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_713
timestamp 1688980957
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_725
timestamp 1688980957
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_3
timestamp 1688980957
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_15
timestamp 1688980957
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_27
timestamp 1688980957
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_39
timestamp 1688980957
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_51
timestamp 1688980957
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_55
timestamp 1688980957
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_57
timestamp 1688980957
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_69
timestamp 1688980957
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_81
timestamp 1688980957
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_93
timestamp 1688980957
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_105
timestamp 1688980957
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_111
timestamp 1688980957
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_113
timestamp 1688980957
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_125
timestamp 1688980957
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_137
timestamp 1688980957
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_149
timestamp 1688980957
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_161
timestamp 1688980957
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_167
timestamp 1688980957
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_169
timestamp 1688980957
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_181
timestamp 1688980957
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_193
timestamp 1688980957
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_205
timestamp 1688980957
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_217
timestamp 1688980957
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_223
timestamp 1688980957
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_225
timestamp 1688980957
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_237
timestamp 1688980957
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_249
timestamp 1688980957
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_261
timestamp 1688980957
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_273
timestamp 1688980957
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_279
timestamp 1688980957
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_281
timestamp 1688980957
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_293
timestamp 1688980957
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_305
timestamp 1688980957
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_317
timestamp 1688980957
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_329
timestamp 1688980957
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_335
timestamp 1688980957
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_337
timestamp 1688980957
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_349
timestamp 1688980957
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_361
timestamp 1688980957
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_373
timestamp 1688980957
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_385
timestamp 1688980957
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_391
timestamp 1688980957
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_393
timestamp 1688980957
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_405
timestamp 1688980957
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_417
timestamp 1688980957
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_429
timestamp 1688980957
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_441
timestamp 1688980957
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_447
timestamp 1688980957
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_449
timestamp 1688980957
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_461
timestamp 1688980957
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_473
timestamp 1688980957
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_485
timestamp 1688980957
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_497
timestamp 1688980957
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_503
timestamp 1688980957
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_505
timestamp 1688980957
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_517
timestamp 1688980957
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_529
timestamp 1688980957
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_541
timestamp 1688980957
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_553
timestamp 1688980957
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_559
timestamp 1688980957
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_561
timestamp 1688980957
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_573
timestamp 1688980957
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_585
timestamp 1688980957
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_597
timestamp 1688980957
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_609
timestamp 1688980957
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_615
timestamp 1688980957
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_617
timestamp 1688980957
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_629
timestamp 1688980957
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_641
timestamp 1688980957
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_653
timestamp 1688980957
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_665
timestamp 1688980957
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_671
timestamp 1688980957
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_673
timestamp 1688980957
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_685
timestamp 1688980957
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_697
timestamp 1688980957
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_709
timestamp 1688980957
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_721
timestamp 1688980957
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_727
timestamp 1688980957
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_729
timestamp 1688980957
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_3
timestamp 1688980957
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_15
timestamp 1688980957
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 1688980957
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_29
timestamp 1688980957
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_41
timestamp 1688980957
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_53
timestamp 1688980957
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_65
timestamp 1688980957
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_77
timestamp 1688980957
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_83
timestamp 1688980957
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_85
timestamp 1688980957
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_97
timestamp 1688980957
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_109
timestamp 1688980957
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_121
timestamp 1688980957
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_133
timestamp 1688980957
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_139
timestamp 1688980957
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_141
timestamp 1688980957
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_153
timestamp 1688980957
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_165
timestamp 1688980957
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_177
timestamp 1688980957
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_189
timestamp 1688980957
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_195
timestamp 1688980957
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_197
timestamp 1688980957
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_209
timestamp 1688980957
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_221
timestamp 1688980957
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_233
timestamp 1688980957
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_245
timestamp 1688980957
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_251
timestamp 1688980957
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_253
timestamp 1688980957
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_265
timestamp 1688980957
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_277
timestamp 1688980957
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_289
timestamp 1688980957
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_301
timestamp 1688980957
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_307
timestamp 1688980957
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_309
timestamp 1688980957
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_321
timestamp 1688980957
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_333
timestamp 1688980957
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_345
timestamp 1688980957
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_357
timestamp 1688980957
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_363
timestamp 1688980957
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_365
timestamp 1688980957
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_377
timestamp 1688980957
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_389
timestamp 1688980957
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_401
timestamp 1688980957
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_413
timestamp 1688980957
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_419
timestamp 1688980957
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_421
timestamp 1688980957
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_433
timestamp 1688980957
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_445
timestamp 1688980957
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_457
timestamp 1688980957
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_469
timestamp 1688980957
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_475
timestamp 1688980957
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_477
timestamp 1688980957
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_489
timestamp 1688980957
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_501
timestamp 1688980957
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_513
timestamp 1688980957
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_525
timestamp 1688980957
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_531
timestamp 1688980957
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_533
timestamp 1688980957
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_545
timestamp 1688980957
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_557
timestamp 1688980957
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_569
timestamp 1688980957
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_581
timestamp 1688980957
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_587
timestamp 1688980957
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_589
timestamp 1688980957
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_601
timestamp 1688980957
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_613
timestamp 1688980957
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_625
timestamp 1688980957
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_637
timestamp 1688980957
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_643
timestamp 1688980957
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_645
timestamp 1688980957
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_657
timestamp 1688980957
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_669
timestamp 1688980957
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_681
timestamp 1688980957
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_693
timestamp 1688980957
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_699
timestamp 1688980957
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_701
timestamp 1688980957
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_713
timestamp 1688980957
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_725
timestamp 1688980957
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_3
timestamp 1688980957
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_15
timestamp 1688980957
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_27
timestamp 1688980957
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_39
timestamp 1688980957
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_51
timestamp 1688980957
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_55
timestamp 1688980957
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 1688980957
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 1688980957
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 1688980957
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_93
timestamp 1688980957
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_105
timestamp 1688980957
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_111
timestamp 1688980957
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_113
timestamp 1688980957
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_125
timestamp 1688980957
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_137
timestamp 1688980957
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_149
timestamp 1688980957
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_161
timestamp 1688980957
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_167
timestamp 1688980957
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_169
timestamp 1688980957
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_181
timestamp 1688980957
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_193
timestamp 1688980957
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_205
timestamp 1688980957
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_217
timestamp 1688980957
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_223
timestamp 1688980957
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_225
timestamp 1688980957
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_237
timestamp 1688980957
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_249
timestamp 1688980957
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_261
timestamp 1688980957
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_273
timestamp 1688980957
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_279
timestamp 1688980957
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_281
timestamp 1688980957
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_293
timestamp 1688980957
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_305
timestamp 1688980957
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_317
timestamp 1688980957
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_329
timestamp 1688980957
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_335
timestamp 1688980957
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_337
timestamp 1688980957
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_349
timestamp 1688980957
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_361
timestamp 1688980957
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_373
timestamp 1688980957
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_385
timestamp 1688980957
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_391
timestamp 1688980957
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_393
timestamp 1688980957
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_405
timestamp 1688980957
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_417
timestamp 1688980957
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_429
timestamp 1688980957
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_441
timestamp 1688980957
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_447
timestamp 1688980957
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_449
timestamp 1688980957
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_461
timestamp 1688980957
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_473
timestamp 1688980957
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_485
timestamp 1688980957
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_497
timestamp 1688980957
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_503
timestamp 1688980957
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_505
timestamp 1688980957
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_517
timestamp 1688980957
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_529
timestamp 1688980957
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_541
timestamp 1688980957
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_553
timestamp 1688980957
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_559
timestamp 1688980957
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_561
timestamp 1688980957
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_573
timestamp 1688980957
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_585
timestamp 1688980957
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_597
timestamp 1688980957
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_609
timestamp 1688980957
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_615
timestamp 1688980957
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_617
timestamp 1688980957
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_629
timestamp 1688980957
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_641
timestamp 1688980957
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_653
timestamp 1688980957
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_665
timestamp 1688980957
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_671
timestamp 1688980957
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_673
timestamp 1688980957
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_685
timestamp 1688980957
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_697
timestamp 1688980957
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_709
timestamp 1688980957
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_721
timestamp 1688980957
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_727
timestamp 1688980957
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_729
timestamp 1688980957
transform 1 0 68172 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_3
timestamp 1688980957
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_15
timestamp 1688980957
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 1688980957
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_29
timestamp 1688980957
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_41
timestamp 1688980957
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_53
timestamp 1688980957
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_65
timestamp 1688980957
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_77
timestamp 1688980957
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_83
timestamp 1688980957
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_85
timestamp 1688980957
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_97
timestamp 1688980957
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_109
timestamp 1688980957
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_121
timestamp 1688980957
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_133
timestamp 1688980957
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_139
timestamp 1688980957
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_141
timestamp 1688980957
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_153
timestamp 1688980957
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_165
timestamp 1688980957
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_177
timestamp 1688980957
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_189
timestamp 1688980957
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_195
timestamp 1688980957
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_197
timestamp 1688980957
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_209
timestamp 1688980957
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_221
timestamp 1688980957
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_233
timestamp 1688980957
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_245
timestamp 1688980957
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_251
timestamp 1688980957
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_253
timestamp 1688980957
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_265
timestamp 1688980957
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_277
timestamp 1688980957
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_289
timestamp 1688980957
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_301
timestamp 1688980957
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_307
timestamp 1688980957
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_309
timestamp 1688980957
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_321
timestamp 1688980957
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_333
timestamp 1688980957
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_345
timestamp 1688980957
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_357
timestamp 1688980957
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_363
timestamp 1688980957
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_365
timestamp 1688980957
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_377
timestamp 1688980957
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_389
timestamp 1688980957
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_401
timestamp 1688980957
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_413
timestamp 1688980957
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_419
timestamp 1688980957
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_421
timestamp 1688980957
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_433
timestamp 1688980957
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_445
timestamp 1688980957
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_457
timestamp 1688980957
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_469
timestamp 1688980957
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_475
timestamp 1688980957
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_477
timestamp 1688980957
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_489
timestamp 1688980957
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_501
timestamp 1688980957
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_513
timestamp 1688980957
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_525
timestamp 1688980957
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_531
timestamp 1688980957
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_533
timestamp 1688980957
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_545
timestamp 1688980957
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_557
timestamp 1688980957
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_569
timestamp 1688980957
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_581
timestamp 1688980957
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_587
timestamp 1688980957
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_589
timestamp 1688980957
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_601
timestamp 1688980957
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_613
timestamp 1688980957
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_625
timestamp 1688980957
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_637
timestamp 1688980957
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_643
timestamp 1688980957
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_645
timestamp 1688980957
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_657
timestamp 1688980957
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_669
timestamp 1688980957
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_681
timestamp 1688980957
transform 1 0 63756 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_693
timestamp 1688980957
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_699
timestamp 1688980957
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_701
timestamp 1688980957
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_713
timestamp 1688980957
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_725
timestamp 1688980957
transform 1 0 67804 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_3
timestamp 1688980957
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_15
timestamp 1688980957
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_27
timestamp 1688980957
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_39
timestamp 1688980957
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_51
timestamp 1688980957
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_55
timestamp 1688980957
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_57
timestamp 1688980957
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_69
timestamp 1688980957
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_81
timestamp 1688980957
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_93
timestamp 1688980957
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_105
timestamp 1688980957
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_111
timestamp 1688980957
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_113
timestamp 1688980957
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_125
timestamp 1688980957
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_137
timestamp 1688980957
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_149
timestamp 1688980957
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_161
timestamp 1688980957
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_167
timestamp 1688980957
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_169
timestamp 1688980957
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_181
timestamp 1688980957
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_193
timestamp 1688980957
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_205
timestamp 1688980957
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_217
timestamp 1688980957
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_223
timestamp 1688980957
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_225
timestamp 1688980957
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_237
timestamp 1688980957
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_249
timestamp 1688980957
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_261
timestamp 1688980957
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_273
timestamp 1688980957
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_279
timestamp 1688980957
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_281
timestamp 1688980957
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_293
timestamp 1688980957
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_305
timestamp 1688980957
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_317
timestamp 1688980957
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_329
timestamp 1688980957
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_335
timestamp 1688980957
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_337
timestamp 1688980957
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_349
timestamp 1688980957
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_361
timestamp 1688980957
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_373
timestamp 1688980957
transform 1 0 35420 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_385
timestamp 1688980957
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_391
timestamp 1688980957
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_393
timestamp 1688980957
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_405
timestamp 1688980957
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_417
timestamp 1688980957
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_429
timestamp 1688980957
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_441
timestamp 1688980957
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_447
timestamp 1688980957
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_449
timestamp 1688980957
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_461
timestamp 1688980957
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_473
timestamp 1688980957
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_485
timestamp 1688980957
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_497
timestamp 1688980957
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_503
timestamp 1688980957
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_505
timestamp 1688980957
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_517
timestamp 1688980957
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_529
timestamp 1688980957
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_541
timestamp 1688980957
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_553
timestamp 1688980957
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_559
timestamp 1688980957
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_561
timestamp 1688980957
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_573
timestamp 1688980957
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_585
timestamp 1688980957
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_597
timestamp 1688980957
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_609
timestamp 1688980957
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_615
timestamp 1688980957
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_617
timestamp 1688980957
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_629
timestamp 1688980957
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_641
timestamp 1688980957
transform 1 0 60076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_653
timestamp 1688980957
transform 1 0 61180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_665
timestamp 1688980957
transform 1 0 62284 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_671
timestamp 1688980957
transform 1 0 62836 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_673
timestamp 1688980957
transform 1 0 63020 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_685
timestamp 1688980957
transform 1 0 64124 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_697
timestamp 1688980957
transform 1 0 65228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_709
timestamp 1688980957
transform 1 0 66332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_721
timestamp 1688980957
transform 1 0 67436 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_727
timestamp 1688980957
transform 1 0 67988 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_729
timestamp 1688980957
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_3
timestamp 1688980957
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_15
timestamp 1688980957
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_27
timestamp 1688980957
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_29
timestamp 1688980957
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_41
timestamp 1688980957
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_53
timestamp 1688980957
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_65
timestamp 1688980957
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_77
timestamp 1688980957
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_83
timestamp 1688980957
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_85
timestamp 1688980957
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_97
timestamp 1688980957
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_109
timestamp 1688980957
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_121
timestamp 1688980957
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_133
timestamp 1688980957
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_139
timestamp 1688980957
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_141
timestamp 1688980957
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_153
timestamp 1688980957
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_165
timestamp 1688980957
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_177
timestamp 1688980957
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_189
timestamp 1688980957
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_195
timestamp 1688980957
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_197
timestamp 1688980957
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_209
timestamp 1688980957
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_221
timestamp 1688980957
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_233
timestamp 1688980957
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_245
timestamp 1688980957
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_251
timestamp 1688980957
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_253
timestamp 1688980957
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_265
timestamp 1688980957
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_277
timestamp 1688980957
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_289
timestamp 1688980957
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_301
timestamp 1688980957
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_307
timestamp 1688980957
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_309
timestamp 1688980957
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_321
timestamp 1688980957
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_333
timestamp 1688980957
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_345
timestamp 1688980957
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_357
timestamp 1688980957
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_363
timestamp 1688980957
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_365
timestamp 1688980957
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_377
timestamp 1688980957
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_389
timestamp 1688980957
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_401
timestamp 1688980957
transform 1 0 37996 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_413
timestamp 1688980957
transform 1 0 39100 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_419
timestamp 1688980957
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_421
timestamp 1688980957
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_433
timestamp 1688980957
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_445
timestamp 1688980957
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_457
timestamp 1688980957
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_469
timestamp 1688980957
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_475
timestamp 1688980957
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_477
timestamp 1688980957
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_489
timestamp 1688980957
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_501
timestamp 1688980957
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_513
timestamp 1688980957
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_525
timestamp 1688980957
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_531
timestamp 1688980957
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_533
timestamp 1688980957
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_545
timestamp 1688980957
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_557
timestamp 1688980957
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_569
timestamp 1688980957
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_581
timestamp 1688980957
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_587
timestamp 1688980957
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_589
timestamp 1688980957
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_601
timestamp 1688980957
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_613
timestamp 1688980957
transform 1 0 57500 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_625
timestamp 1688980957
transform 1 0 58604 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_637
timestamp 1688980957
transform 1 0 59708 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_643
timestamp 1688980957
transform 1 0 60260 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_645
timestamp 1688980957
transform 1 0 60444 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_657
timestamp 1688980957
transform 1 0 61548 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_669
timestamp 1688980957
transform 1 0 62652 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_681
timestamp 1688980957
transform 1 0 63756 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_693
timestamp 1688980957
transform 1 0 64860 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_699
timestamp 1688980957
transform 1 0 65412 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_701
timestamp 1688980957
transform 1 0 65596 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_713
timestamp 1688980957
transform 1 0 66700 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_725
timestamp 1688980957
transform 1 0 67804 0 1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_3
timestamp 1688980957
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_15
timestamp 1688980957
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_27
timestamp 1688980957
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_39
timestamp 1688980957
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_51
timestamp 1688980957
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_55
timestamp 1688980957
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_57
timestamp 1688980957
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_69
timestamp 1688980957
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_81
timestamp 1688980957
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_93
timestamp 1688980957
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_105
timestamp 1688980957
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_111
timestamp 1688980957
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_113
timestamp 1688980957
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_125
timestamp 1688980957
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_137
timestamp 1688980957
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_149
timestamp 1688980957
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_161
timestamp 1688980957
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_167
timestamp 1688980957
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_169
timestamp 1688980957
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_181
timestamp 1688980957
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_193
timestamp 1688980957
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_205
timestamp 1688980957
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_217
timestamp 1688980957
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_223
timestamp 1688980957
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_225
timestamp 1688980957
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_237
timestamp 1688980957
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_249
timestamp 1688980957
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_261
timestamp 1688980957
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_273
timestamp 1688980957
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_279
timestamp 1688980957
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_281
timestamp 1688980957
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_293
timestamp 1688980957
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_305
timestamp 1688980957
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_317
timestamp 1688980957
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_329
timestamp 1688980957
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_335
timestamp 1688980957
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_337
timestamp 1688980957
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_349
timestamp 1688980957
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_361
timestamp 1688980957
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_373
timestamp 1688980957
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_385
timestamp 1688980957
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_391
timestamp 1688980957
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_393
timestamp 1688980957
transform 1 0 37260 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_405
timestamp 1688980957
transform 1 0 38364 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_417
timestamp 1688980957
transform 1 0 39468 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_429
timestamp 1688980957
transform 1 0 40572 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_441
timestamp 1688980957
transform 1 0 41676 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_447
timestamp 1688980957
transform 1 0 42228 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_449
timestamp 1688980957
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_461
timestamp 1688980957
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_473
timestamp 1688980957
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_485
timestamp 1688980957
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_497
timestamp 1688980957
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_503
timestamp 1688980957
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_505
timestamp 1688980957
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_517
timestamp 1688980957
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_529
timestamp 1688980957
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_541
timestamp 1688980957
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_553
timestamp 1688980957
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_559
timestamp 1688980957
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_561
timestamp 1688980957
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_573
timestamp 1688980957
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_585
timestamp 1688980957
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_597
timestamp 1688980957
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_609
timestamp 1688980957
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_615
timestamp 1688980957
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_617
timestamp 1688980957
transform 1 0 57868 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_629
timestamp 1688980957
transform 1 0 58972 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_641
timestamp 1688980957
transform 1 0 60076 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_653
timestamp 1688980957
transform 1 0 61180 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_665
timestamp 1688980957
transform 1 0 62284 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_671
timestamp 1688980957
transform 1 0 62836 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_673
timestamp 1688980957
transform 1 0 63020 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_685
timestamp 1688980957
transform 1 0 64124 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_697
timestamp 1688980957
transform 1 0 65228 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_709
timestamp 1688980957
transform 1 0 66332 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_721
timestamp 1688980957
transform 1 0 67436 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_727
timestamp 1688980957
transform 1 0 67988 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_729
timestamp 1688980957
transform 1 0 68172 0 -1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_3
timestamp 1688980957
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_15
timestamp 1688980957
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_27
timestamp 1688980957
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_29
timestamp 1688980957
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_41
timestamp 1688980957
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_53
timestamp 1688980957
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_65
timestamp 1688980957
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_77
timestamp 1688980957
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_83
timestamp 1688980957
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_85
timestamp 1688980957
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_97
timestamp 1688980957
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_109
timestamp 1688980957
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_121
timestamp 1688980957
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_133
timestamp 1688980957
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_139
timestamp 1688980957
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_141
timestamp 1688980957
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_153
timestamp 1688980957
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_165
timestamp 1688980957
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_177
timestamp 1688980957
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_189
timestamp 1688980957
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_195
timestamp 1688980957
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_197
timestamp 1688980957
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_209
timestamp 1688980957
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_221
timestamp 1688980957
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_233
timestamp 1688980957
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_245
timestamp 1688980957
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_251
timestamp 1688980957
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_253
timestamp 1688980957
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_265
timestamp 1688980957
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_277
timestamp 1688980957
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_289
timestamp 1688980957
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_301
timestamp 1688980957
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_307
timestamp 1688980957
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_309
timestamp 1688980957
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_321
timestamp 1688980957
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_333
timestamp 1688980957
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_345
timestamp 1688980957
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_357
timestamp 1688980957
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_363
timestamp 1688980957
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_365
timestamp 1688980957
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_377
timestamp 1688980957
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_389
timestamp 1688980957
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_401
timestamp 1688980957
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_413
timestamp 1688980957
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_419
timestamp 1688980957
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_421
timestamp 1688980957
transform 1 0 39836 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_433
timestamp 1688980957
transform 1 0 40940 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_445
timestamp 1688980957
transform 1 0 42044 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_457
timestamp 1688980957
transform 1 0 43148 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_469
timestamp 1688980957
transform 1 0 44252 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_475
timestamp 1688980957
transform 1 0 44804 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_477
timestamp 1688980957
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_489
timestamp 1688980957
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_501
timestamp 1688980957
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_513
timestamp 1688980957
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_525
timestamp 1688980957
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_531
timestamp 1688980957
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_533
timestamp 1688980957
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_545
timestamp 1688980957
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_557
timestamp 1688980957
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_569
timestamp 1688980957
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_581
timestamp 1688980957
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_587
timestamp 1688980957
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_589
timestamp 1688980957
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_601
timestamp 1688980957
transform 1 0 56396 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_613
timestamp 1688980957
transform 1 0 57500 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_625
timestamp 1688980957
transform 1 0 58604 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_637
timestamp 1688980957
transform 1 0 59708 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_643
timestamp 1688980957
transform 1 0 60260 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_645
timestamp 1688980957
transform 1 0 60444 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_657
timestamp 1688980957
transform 1 0 61548 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_669
timestamp 1688980957
transform 1 0 62652 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_681
timestamp 1688980957
transform 1 0 63756 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_693
timestamp 1688980957
transform 1 0 64860 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_699
timestamp 1688980957
transform 1 0 65412 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_701
timestamp 1688980957
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_713
timestamp 1688980957
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_725
timestamp 1688980957
transform 1 0 67804 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_3
timestamp 1688980957
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_15
timestamp 1688980957
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_27
timestamp 1688980957
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_39
timestamp 1688980957
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105_51
timestamp 1688980957
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_55
timestamp 1688980957
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_57
timestamp 1688980957
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_69
timestamp 1688980957
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_81
timestamp 1688980957
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_93
timestamp 1688980957
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_105
timestamp 1688980957
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_111
timestamp 1688980957
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_113
timestamp 1688980957
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_125
timestamp 1688980957
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_137
timestamp 1688980957
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_149
timestamp 1688980957
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_161
timestamp 1688980957
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_167
timestamp 1688980957
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_169
timestamp 1688980957
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_181
timestamp 1688980957
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_193
timestamp 1688980957
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_205
timestamp 1688980957
transform 1 0 19964 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_217
timestamp 1688980957
transform 1 0 21068 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_223
timestamp 1688980957
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_225
timestamp 1688980957
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_237
timestamp 1688980957
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_249
timestamp 1688980957
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_261
timestamp 1688980957
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_273
timestamp 1688980957
transform 1 0 26220 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_279
timestamp 1688980957
transform 1 0 26772 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_281
timestamp 1688980957
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_293
timestamp 1688980957
transform 1 0 28060 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_305
timestamp 1688980957
transform 1 0 29164 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_317
timestamp 1688980957
transform 1 0 30268 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_329
timestamp 1688980957
transform 1 0 31372 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_335
timestamp 1688980957
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_337
timestamp 1688980957
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_349
timestamp 1688980957
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_361
timestamp 1688980957
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_373
timestamp 1688980957
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_385
timestamp 1688980957
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_391
timestamp 1688980957
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_393
timestamp 1688980957
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_405
timestamp 1688980957
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_417
timestamp 1688980957
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_429
timestamp 1688980957
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_441
timestamp 1688980957
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_447
timestamp 1688980957
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_449
timestamp 1688980957
transform 1 0 42412 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_461
timestamp 1688980957
transform 1 0 43516 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_473
timestamp 1688980957
transform 1 0 44620 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_485
timestamp 1688980957
transform 1 0 45724 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_497
timestamp 1688980957
transform 1 0 46828 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_503
timestamp 1688980957
transform 1 0 47380 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_505
timestamp 1688980957
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_517
timestamp 1688980957
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_529
timestamp 1688980957
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_541
timestamp 1688980957
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_553
timestamp 1688980957
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_559
timestamp 1688980957
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_561
timestamp 1688980957
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_573
timestamp 1688980957
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_585
timestamp 1688980957
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_597
timestamp 1688980957
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_609
timestamp 1688980957
transform 1 0 57132 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_615
timestamp 1688980957
transform 1 0 57684 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_617
timestamp 1688980957
transform 1 0 57868 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_629
timestamp 1688980957
transform 1 0 58972 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_641
timestamp 1688980957
transform 1 0 60076 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_653
timestamp 1688980957
transform 1 0 61180 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_665
timestamp 1688980957
transform 1 0 62284 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_671
timestamp 1688980957
transform 1 0 62836 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_673
timestamp 1688980957
transform 1 0 63020 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_685
timestamp 1688980957
transform 1 0 64124 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_697
timestamp 1688980957
transform 1 0 65228 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_709
timestamp 1688980957
transform 1 0 66332 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_721
timestamp 1688980957
transform 1 0 67436 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_727
timestamp 1688980957
transform 1 0 67988 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105_729
timestamp 1688980957
transform 1 0 68172 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_3
timestamp 1688980957
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_15
timestamp 1688980957
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_27
timestamp 1688980957
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_29
timestamp 1688980957
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_41
timestamp 1688980957
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_53
timestamp 1688980957
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_65
timestamp 1688980957
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_77
timestamp 1688980957
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_83
timestamp 1688980957
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_85
timestamp 1688980957
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_97
timestamp 1688980957
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_109
timestamp 1688980957
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_121
timestamp 1688980957
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_133
timestamp 1688980957
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_139
timestamp 1688980957
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_141
timestamp 1688980957
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_153
timestamp 1688980957
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_165
timestamp 1688980957
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_177
timestamp 1688980957
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_189
timestamp 1688980957
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_195
timestamp 1688980957
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_197
timestamp 1688980957
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_209
timestamp 1688980957
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_221
timestamp 1688980957
transform 1 0 21436 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_233
timestamp 1688980957
transform 1 0 22540 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_245
timestamp 1688980957
transform 1 0 23644 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_251
timestamp 1688980957
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_253
timestamp 1688980957
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_265
timestamp 1688980957
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_277
timestamp 1688980957
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_289
timestamp 1688980957
transform 1 0 27692 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_301
timestamp 1688980957
transform 1 0 28796 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_307
timestamp 1688980957
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_309
timestamp 1688980957
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_321
timestamp 1688980957
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_333
timestamp 1688980957
transform 1 0 31740 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_345
timestamp 1688980957
transform 1 0 32844 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_357
timestamp 1688980957
transform 1 0 33948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_363
timestamp 1688980957
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_365
timestamp 1688980957
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_377
timestamp 1688980957
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_389
timestamp 1688980957
transform 1 0 36892 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_401
timestamp 1688980957
transform 1 0 37996 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_413
timestamp 1688980957
transform 1 0 39100 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_419
timestamp 1688980957
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_421
timestamp 1688980957
transform 1 0 39836 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_433
timestamp 1688980957
transform 1 0 40940 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_445
timestamp 1688980957
transform 1 0 42044 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_457
timestamp 1688980957
transform 1 0 43148 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_469
timestamp 1688980957
transform 1 0 44252 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_475
timestamp 1688980957
transform 1 0 44804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_477
timestamp 1688980957
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_489
timestamp 1688980957
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_501
timestamp 1688980957
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_513
timestamp 1688980957
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_525
timestamp 1688980957
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_531
timestamp 1688980957
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_533
timestamp 1688980957
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_545
timestamp 1688980957
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_557
timestamp 1688980957
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_569
timestamp 1688980957
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_581
timestamp 1688980957
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_587
timestamp 1688980957
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_589
timestamp 1688980957
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_601
timestamp 1688980957
transform 1 0 56396 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_613
timestamp 1688980957
transform 1 0 57500 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_625
timestamp 1688980957
transform 1 0 58604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_637
timestamp 1688980957
transform 1 0 59708 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_643
timestamp 1688980957
transform 1 0 60260 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_645
timestamp 1688980957
transform 1 0 60444 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_657
timestamp 1688980957
transform 1 0 61548 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_669
timestamp 1688980957
transform 1 0 62652 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_681
timestamp 1688980957
transform 1 0 63756 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_693
timestamp 1688980957
transform 1 0 64860 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_699
timestamp 1688980957
transform 1 0 65412 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_701
timestamp 1688980957
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_713
timestamp 1688980957
transform 1 0 66700 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_725
timestamp 1688980957
transform 1 0 67804 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_3
timestamp 1688980957
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_15
timestamp 1688980957
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_27
timestamp 1688980957
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_39
timestamp 1688980957
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_51
timestamp 1688980957
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_55
timestamp 1688980957
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_57
timestamp 1688980957
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_69
timestamp 1688980957
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_81
timestamp 1688980957
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_93
timestamp 1688980957
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_105
timestamp 1688980957
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_111
timestamp 1688980957
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_113
timestamp 1688980957
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_125
timestamp 1688980957
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_137
timestamp 1688980957
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_149
timestamp 1688980957
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_161
timestamp 1688980957
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_167
timestamp 1688980957
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_169
timestamp 1688980957
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_181
timestamp 1688980957
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_193
timestamp 1688980957
transform 1 0 18860 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_205
timestamp 1688980957
transform 1 0 19964 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_217
timestamp 1688980957
transform 1 0 21068 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_223
timestamp 1688980957
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_225
timestamp 1688980957
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_237
timestamp 1688980957
transform 1 0 22908 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_249
timestamp 1688980957
transform 1 0 24012 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_261
timestamp 1688980957
transform 1 0 25116 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_273
timestamp 1688980957
transform 1 0 26220 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_279
timestamp 1688980957
transform 1 0 26772 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_281
timestamp 1688980957
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_293
timestamp 1688980957
transform 1 0 28060 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_305
timestamp 1688980957
transform 1 0 29164 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_317
timestamp 1688980957
transform 1 0 30268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_329
timestamp 1688980957
transform 1 0 31372 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_335
timestamp 1688980957
transform 1 0 31924 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_337
timestamp 1688980957
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_349
timestamp 1688980957
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_361
timestamp 1688980957
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_373
timestamp 1688980957
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_385
timestamp 1688980957
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_391
timestamp 1688980957
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_393
timestamp 1688980957
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_405
timestamp 1688980957
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_417
timestamp 1688980957
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_429
timestamp 1688980957
transform 1 0 40572 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_441
timestamp 1688980957
transform 1 0 41676 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_447
timestamp 1688980957
transform 1 0 42228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_449
timestamp 1688980957
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_461
timestamp 1688980957
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_473
timestamp 1688980957
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_485
timestamp 1688980957
transform 1 0 45724 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_497
timestamp 1688980957
transform 1 0 46828 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_503
timestamp 1688980957
transform 1 0 47380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_505
timestamp 1688980957
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_517
timestamp 1688980957
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_529
timestamp 1688980957
transform 1 0 49772 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_541
timestamp 1688980957
transform 1 0 50876 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_553
timestamp 1688980957
transform 1 0 51980 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_559
timestamp 1688980957
transform 1 0 52532 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_561
timestamp 1688980957
transform 1 0 52716 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_573
timestamp 1688980957
transform 1 0 53820 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_585
timestamp 1688980957
transform 1 0 54924 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_597
timestamp 1688980957
transform 1 0 56028 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_609
timestamp 1688980957
transform 1 0 57132 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_615
timestamp 1688980957
transform 1 0 57684 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_617
timestamp 1688980957
transform 1 0 57868 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_629
timestamp 1688980957
transform 1 0 58972 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_641
timestamp 1688980957
transform 1 0 60076 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_653
timestamp 1688980957
transform 1 0 61180 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_665
timestamp 1688980957
transform 1 0 62284 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_671
timestamp 1688980957
transform 1 0 62836 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_673
timestamp 1688980957
transform 1 0 63020 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_685
timestamp 1688980957
transform 1 0 64124 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_697
timestamp 1688980957
transform 1 0 65228 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_709
timestamp 1688980957
transform 1 0 66332 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_721
timestamp 1688980957
transform 1 0 67436 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_727
timestamp 1688980957
transform 1 0 67988 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_729
timestamp 1688980957
transform 1 0 68172 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_3
timestamp 1688980957
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_15
timestamp 1688980957
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_27
timestamp 1688980957
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_29
timestamp 1688980957
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_41
timestamp 1688980957
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_53
timestamp 1688980957
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_65
timestamp 1688980957
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_77
timestamp 1688980957
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_83
timestamp 1688980957
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_85
timestamp 1688980957
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_97
timestamp 1688980957
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_109
timestamp 1688980957
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_121
timestamp 1688980957
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_133
timestamp 1688980957
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_139
timestamp 1688980957
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_141
timestamp 1688980957
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_153
timestamp 1688980957
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_165
timestamp 1688980957
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_177
timestamp 1688980957
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_189
timestamp 1688980957
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_195
timestamp 1688980957
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_197
timestamp 1688980957
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_209
timestamp 1688980957
transform 1 0 20332 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_221
timestamp 1688980957
transform 1 0 21436 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_233
timestamp 1688980957
transform 1 0 22540 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_245
timestamp 1688980957
transform 1 0 23644 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_251
timestamp 1688980957
transform 1 0 24196 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_253
timestamp 1688980957
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_265
timestamp 1688980957
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_277
timestamp 1688980957
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_289
timestamp 1688980957
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_301
timestamp 1688980957
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_307
timestamp 1688980957
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_309
timestamp 1688980957
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_321
timestamp 1688980957
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_333
timestamp 1688980957
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_345
timestamp 1688980957
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_357
timestamp 1688980957
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_363
timestamp 1688980957
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_365
timestamp 1688980957
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_377
timestamp 1688980957
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_389
timestamp 1688980957
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_401
timestamp 1688980957
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_413
timestamp 1688980957
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_419
timestamp 1688980957
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_421
timestamp 1688980957
transform 1 0 39836 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_433
timestamp 1688980957
transform 1 0 40940 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_445
timestamp 1688980957
transform 1 0 42044 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_457
timestamp 1688980957
transform 1 0 43148 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_469
timestamp 1688980957
transform 1 0 44252 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_475
timestamp 1688980957
transform 1 0 44804 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_477
timestamp 1688980957
transform 1 0 44988 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_489
timestamp 1688980957
transform 1 0 46092 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_501
timestamp 1688980957
transform 1 0 47196 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_513
timestamp 1688980957
transform 1 0 48300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_525
timestamp 1688980957
transform 1 0 49404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_531
timestamp 1688980957
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_533
timestamp 1688980957
transform 1 0 50140 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_545
timestamp 1688980957
transform 1 0 51244 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_557
timestamp 1688980957
transform 1 0 52348 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_569
timestamp 1688980957
transform 1 0 53452 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_581
timestamp 1688980957
transform 1 0 54556 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_587
timestamp 1688980957
transform 1 0 55108 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_589
timestamp 1688980957
transform 1 0 55292 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_601
timestamp 1688980957
transform 1 0 56396 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_613
timestamp 1688980957
transform 1 0 57500 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_625
timestamp 1688980957
transform 1 0 58604 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_637
timestamp 1688980957
transform 1 0 59708 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_643
timestamp 1688980957
transform 1 0 60260 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_645
timestamp 1688980957
transform 1 0 60444 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_657
timestamp 1688980957
transform 1 0 61548 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_669
timestamp 1688980957
transform 1 0 62652 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_681
timestamp 1688980957
transform 1 0 63756 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_693
timestamp 1688980957
transform 1 0 64860 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_699
timestamp 1688980957
transform 1 0 65412 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_701
timestamp 1688980957
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_713
timestamp 1688980957
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_725
timestamp 1688980957
transform 1 0 67804 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_3
timestamp 1688980957
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_15
timestamp 1688980957
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_27
timestamp 1688980957
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_39
timestamp 1688980957
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_51
timestamp 1688980957
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_55
timestamp 1688980957
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_57
timestamp 1688980957
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_69
timestamp 1688980957
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_81
timestamp 1688980957
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_93
timestamp 1688980957
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_105
timestamp 1688980957
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_111
timestamp 1688980957
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_113
timestamp 1688980957
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_125
timestamp 1688980957
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_137
timestamp 1688980957
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_149
timestamp 1688980957
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_161
timestamp 1688980957
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_167
timestamp 1688980957
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_169
timestamp 1688980957
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_181
timestamp 1688980957
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_193
timestamp 1688980957
transform 1 0 18860 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_205
timestamp 1688980957
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_217
timestamp 1688980957
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_223
timestamp 1688980957
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_225
timestamp 1688980957
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_237
timestamp 1688980957
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_249
timestamp 1688980957
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_261
timestamp 1688980957
transform 1 0 25116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_273
timestamp 1688980957
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_279
timestamp 1688980957
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_281
timestamp 1688980957
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_293
timestamp 1688980957
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_305
timestamp 1688980957
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_317
timestamp 1688980957
transform 1 0 30268 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_329
timestamp 1688980957
transform 1 0 31372 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_335
timestamp 1688980957
transform 1 0 31924 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_337
timestamp 1688980957
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_349
timestamp 1688980957
transform 1 0 33212 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_361
timestamp 1688980957
transform 1 0 34316 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_373
timestamp 1688980957
transform 1 0 35420 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_385
timestamp 1688980957
transform 1 0 36524 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_391
timestamp 1688980957
transform 1 0 37076 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_393
timestamp 1688980957
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_405
timestamp 1688980957
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_417
timestamp 1688980957
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_429
timestamp 1688980957
transform 1 0 40572 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_441
timestamp 1688980957
transform 1 0 41676 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_447
timestamp 1688980957
transform 1 0 42228 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_449
timestamp 1688980957
transform 1 0 42412 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_461
timestamp 1688980957
transform 1 0 43516 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_473
timestamp 1688980957
transform 1 0 44620 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_485
timestamp 1688980957
transform 1 0 45724 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_497
timestamp 1688980957
transform 1 0 46828 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_503
timestamp 1688980957
transform 1 0 47380 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_505
timestamp 1688980957
transform 1 0 47564 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_517
timestamp 1688980957
transform 1 0 48668 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_529
timestamp 1688980957
transform 1 0 49772 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_541
timestamp 1688980957
transform 1 0 50876 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_553
timestamp 1688980957
transform 1 0 51980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_559
timestamp 1688980957
transform 1 0 52532 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_561
timestamp 1688980957
transform 1 0 52716 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_573
timestamp 1688980957
transform 1 0 53820 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_585
timestamp 1688980957
transform 1 0 54924 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_597
timestamp 1688980957
transform 1 0 56028 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_609
timestamp 1688980957
transform 1 0 57132 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_615
timestamp 1688980957
transform 1 0 57684 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_617
timestamp 1688980957
transform 1 0 57868 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_629
timestamp 1688980957
transform 1 0 58972 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_641
timestamp 1688980957
transform 1 0 60076 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_653
timestamp 1688980957
transform 1 0 61180 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_665
timestamp 1688980957
transform 1 0 62284 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_671
timestamp 1688980957
transform 1 0 62836 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_673
timestamp 1688980957
transform 1 0 63020 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_685
timestamp 1688980957
transform 1 0 64124 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_697
timestamp 1688980957
transform 1 0 65228 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_709
timestamp 1688980957
transform 1 0 66332 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_721
timestamp 1688980957
transform 1 0 67436 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_727
timestamp 1688980957
transform 1 0 67988 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_729
timestamp 1688980957
transform 1 0 68172 0 -1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_3
timestamp 1688980957
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_15
timestamp 1688980957
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_27
timestamp 1688980957
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_29
timestamp 1688980957
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_41
timestamp 1688980957
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_53
timestamp 1688980957
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_65
timestamp 1688980957
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_77
timestamp 1688980957
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_83
timestamp 1688980957
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_85
timestamp 1688980957
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_97
timestamp 1688980957
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_109
timestamp 1688980957
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_121
timestamp 1688980957
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_133
timestamp 1688980957
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_139
timestamp 1688980957
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_141
timestamp 1688980957
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_153
timestamp 1688980957
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_165
timestamp 1688980957
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_177
timestamp 1688980957
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_189
timestamp 1688980957
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_195
timestamp 1688980957
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_197
timestamp 1688980957
transform 1 0 19228 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_209
timestamp 1688980957
transform 1 0 20332 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_221
timestamp 1688980957
transform 1 0 21436 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_233
timestamp 1688980957
transform 1 0 22540 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_245
timestamp 1688980957
transform 1 0 23644 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_251
timestamp 1688980957
transform 1 0 24196 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_253
timestamp 1688980957
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_265
timestamp 1688980957
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_277
timestamp 1688980957
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_289
timestamp 1688980957
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_301
timestamp 1688980957
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_307
timestamp 1688980957
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_309
timestamp 1688980957
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_321
timestamp 1688980957
transform 1 0 30636 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_333
timestamp 1688980957
transform 1 0 31740 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_345
timestamp 1688980957
transform 1 0 32844 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_357
timestamp 1688980957
transform 1 0 33948 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_363
timestamp 1688980957
transform 1 0 34500 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_365
timestamp 1688980957
transform 1 0 34684 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_377
timestamp 1688980957
transform 1 0 35788 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_389
timestamp 1688980957
transform 1 0 36892 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_401
timestamp 1688980957
transform 1 0 37996 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_413
timestamp 1688980957
transform 1 0 39100 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_419
timestamp 1688980957
transform 1 0 39652 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_421
timestamp 1688980957
transform 1 0 39836 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_433
timestamp 1688980957
transform 1 0 40940 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_445
timestamp 1688980957
transform 1 0 42044 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_457
timestamp 1688980957
transform 1 0 43148 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_469
timestamp 1688980957
transform 1 0 44252 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_475
timestamp 1688980957
transform 1 0 44804 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_477
timestamp 1688980957
transform 1 0 44988 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_489
timestamp 1688980957
transform 1 0 46092 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_501
timestamp 1688980957
transform 1 0 47196 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_513
timestamp 1688980957
transform 1 0 48300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_525
timestamp 1688980957
transform 1 0 49404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_531
timestamp 1688980957
transform 1 0 49956 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_533
timestamp 1688980957
transform 1 0 50140 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_545
timestamp 1688980957
transform 1 0 51244 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_557
timestamp 1688980957
transform 1 0 52348 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_569
timestamp 1688980957
transform 1 0 53452 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_581
timestamp 1688980957
transform 1 0 54556 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_587
timestamp 1688980957
transform 1 0 55108 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_589
timestamp 1688980957
transform 1 0 55292 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_601
timestamp 1688980957
transform 1 0 56396 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_613
timestamp 1688980957
transform 1 0 57500 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_625
timestamp 1688980957
transform 1 0 58604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_637
timestamp 1688980957
transform 1 0 59708 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_643
timestamp 1688980957
transform 1 0 60260 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_645
timestamp 1688980957
transform 1 0 60444 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_657
timestamp 1688980957
transform 1 0 61548 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_669
timestamp 1688980957
transform 1 0 62652 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_681
timestamp 1688980957
transform 1 0 63756 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_693
timestamp 1688980957
transform 1 0 64860 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_699
timestamp 1688980957
transform 1 0 65412 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_701
timestamp 1688980957
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_713
timestamp 1688980957
transform 1 0 66700 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_725
timestamp 1688980957
transform 1 0 67804 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_3
timestamp 1688980957
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_15
timestamp 1688980957
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_27
timestamp 1688980957
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_39
timestamp 1688980957
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_51
timestamp 1688980957
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_55
timestamp 1688980957
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_57
timestamp 1688980957
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_69
timestamp 1688980957
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_81
timestamp 1688980957
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_93
timestamp 1688980957
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_105
timestamp 1688980957
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_111
timestamp 1688980957
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_113
timestamp 1688980957
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_125
timestamp 1688980957
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_137
timestamp 1688980957
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_149
timestamp 1688980957
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_161
timestamp 1688980957
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_167
timestamp 1688980957
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_169
timestamp 1688980957
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_181
timestamp 1688980957
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_193
timestamp 1688980957
transform 1 0 18860 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_205
timestamp 1688980957
transform 1 0 19964 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_217
timestamp 1688980957
transform 1 0 21068 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_223
timestamp 1688980957
transform 1 0 21620 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_225
timestamp 1688980957
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_237
timestamp 1688980957
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_249
timestamp 1688980957
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_261
timestamp 1688980957
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_273
timestamp 1688980957
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_279
timestamp 1688980957
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_281
timestamp 1688980957
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_293
timestamp 1688980957
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_305
timestamp 1688980957
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_317
timestamp 1688980957
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_329
timestamp 1688980957
transform 1 0 31372 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_335
timestamp 1688980957
transform 1 0 31924 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_337
timestamp 1688980957
transform 1 0 32108 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_349
timestamp 1688980957
transform 1 0 33212 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_361
timestamp 1688980957
transform 1 0 34316 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_373
timestamp 1688980957
transform 1 0 35420 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_385
timestamp 1688980957
transform 1 0 36524 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_391
timestamp 1688980957
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_393
timestamp 1688980957
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_405
timestamp 1688980957
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_417
timestamp 1688980957
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_429
timestamp 1688980957
transform 1 0 40572 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_441
timestamp 1688980957
transform 1 0 41676 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_447
timestamp 1688980957
transform 1 0 42228 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_449
timestamp 1688980957
transform 1 0 42412 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_461
timestamp 1688980957
transform 1 0 43516 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_473
timestamp 1688980957
transform 1 0 44620 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_485
timestamp 1688980957
transform 1 0 45724 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_497
timestamp 1688980957
transform 1 0 46828 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_503
timestamp 1688980957
transform 1 0 47380 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_505
timestamp 1688980957
transform 1 0 47564 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_517
timestamp 1688980957
transform 1 0 48668 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_529
timestamp 1688980957
transform 1 0 49772 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_541
timestamp 1688980957
transform 1 0 50876 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_553
timestamp 1688980957
transform 1 0 51980 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_559
timestamp 1688980957
transform 1 0 52532 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_561
timestamp 1688980957
transform 1 0 52716 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_573
timestamp 1688980957
transform 1 0 53820 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_585
timestamp 1688980957
transform 1 0 54924 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_597
timestamp 1688980957
transform 1 0 56028 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_609
timestamp 1688980957
transform 1 0 57132 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_615
timestamp 1688980957
transform 1 0 57684 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_617
timestamp 1688980957
transform 1 0 57868 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_629
timestamp 1688980957
transform 1 0 58972 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_641
timestamp 1688980957
transform 1 0 60076 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_653
timestamp 1688980957
transform 1 0 61180 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_665
timestamp 1688980957
transform 1 0 62284 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_671
timestamp 1688980957
transform 1 0 62836 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_673
timestamp 1688980957
transform 1 0 63020 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_685
timestamp 1688980957
transform 1 0 64124 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_697
timestamp 1688980957
transform 1 0 65228 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_709
timestamp 1688980957
transform 1 0 66332 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_721
timestamp 1688980957
transform 1 0 67436 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_727
timestamp 1688980957
transform 1 0 67988 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_729
timestamp 1688980957
transform 1 0 68172 0 -1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_3
timestamp 1688980957
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_15
timestamp 1688980957
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_27
timestamp 1688980957
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_29
timestamp 1688980957
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_41
timestamp 1688980957
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_53
timestamp 1688980957
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_65
timestamp 1688980957
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_77
timestamp 1688980957
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_83
timestamp 1688980957
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_85
timestamp 1688980957
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_97
timestamp 1688980957
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_109
timestamp 1688980957
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_121
timestamp 1688980957
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_133
timestamp 1688980957
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_139
timestamp 1688980957
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_141
timestamp 1688980957
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_153
timestamp 1688980957
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_165
timestamp 1688980957
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_177
timestamp 1688980957
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_189
timestamp 1688980957
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_195
timestamp 1688980957
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_197
timestamp 1688980957
transform 1 0 19228 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_209
timestamp 1688980957
transform 1 0 20332 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_221
timestamp 1688980957
transform 1 0 21436 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_233
timestamp 1688980957
transform 1 0 22540 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_245
timestamp 1688980957
transform 1 0 23644 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_251
timestamp 1688980957
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_253
timestamp 1688980957
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_265
timestamp 1688980957
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_277
timestamp 1688980957
transform 1 0 26588 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_289
timestamp 1688980957
transform 1 0 27692 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_301
timestamp 1688980957
transform 1 0 28796 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_307
timestamp 1688980957
transform 1 0 29348 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_309
timestamp 1688980957
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_321
timestamp 1688980957
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_333
timestamp 1688980957
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_345
timestamp 1688980957
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_357
timestamp 1688980957
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_363
timestamp 1688980957
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_365
timestamp 1688980957
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_377
timestamp 1688980957
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_389
timestamp 1688980957
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_401
timestamp 1688980957
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_413
timestamp 1688980957
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_419
timestamp 1688980957
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_421
timestamp 1688980957
transform 1 0 39836 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_433
timestamp 1688980957
transform 1 0 40940 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_445
timestamp 1688980957
transform 1 0 42044 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_457
timestamp 1688980957
transform 1 0 43148 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_469
timestamp 1688980957
transform 1 0 44252 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_475
timestamp 1688980957
transform 1 0 44804 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_477
timestamp 1688980957
transform 1 0 44988 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_489
timestamp 1688980957
transform 1 0 46092 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_501
timestamp 1688980957
transform 1 0 47196 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_513
timestamp 1688980957
transform 1 0 48300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_525
timestamp 1688980957
transform 1 0 49404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_531
timestamp 1688980957
transform 1 0 49956 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_533
timestamp 1688980957
transform 1 0 50140 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_545
timestamp 1688980957
transform 1 0 51244 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_557
timestamp 1688980957
transform 1 0 52348 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_569
timestamp 1688980957
transform 1 0 53452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_581
timestamp 1688980957
transform 1 0 54556 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_587
timestamp 1688980957
transform 1 0 55108 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_589
timestamp 1688980957
transform 1 0 55292 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_601
timestamp 1688980957
transform 1 0 56396 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_613
timestamp 1688980957
transform 1 0 57500 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_625
timestamp 1688980957
transform 1 0 58604 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_637
timestamp 1688980957
transform 1 0 59708 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_643
timestamp 1688980957
transform 1 0 60260 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_645
timestamp 1688980957
transform 1 0 60444 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_657
timestamp 1688980957
transform 1 0 61548 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_669
timestamp 1688980957
transform 1 0 62652 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_681
timestamp 1688980957
transform 1 0 63756 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_693
timestamp 1688980957
transform 1 0 64860 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_699
timestamp 1688980957
transform 1 0 65412 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_701
timestamp 1688980957
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_713
timestamp 1688980957
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_112_725
timestamp 1688980957
transform 1 0 67804 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_3
timestamp 1688980957
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_15
timestamp 1688980957
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_27
timestamp 1688980957
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_39
timestamp 1688980957
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_51
timestamp 1688980957
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_55
timestamp 1688980957
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_57
timestamp 1688980957
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_69
timestamp 1688980957
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_81
timestamp 1688980957
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_93
timestamp 1688980957
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_105
timestamp 1688980957
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_111
timestamp 1688980957
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_113
timestamp 1688980957
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_125
timestamp 1688980957
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_137
timestamp 1688980957
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_149
timestamp 1688980957
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_161
timestamp 1688980957
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_167
timestamp 1688980957
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_169
timestamp 1688980957
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_181
timestamp 1688980957
transform 1 0 17756 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_193
timestamp 1688980957
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_205
timestamp 1688980957
transform 1 0 19964 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_217
timestamp 1688980957
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_223
timestamp 1688980957
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_225
timestamp 1688980957
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_237
timestamp 1688980957
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_249
timestamp 1688980957
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_261
timestamp 1688980957
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_273
timestamp 1688980957
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_279
timestamp 1688980957
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_281
timestamp 1688980957
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_293
timestamp 1688980957
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_305
timestamp 1688980957
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_317
timestamp 1688980957
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_329
timestamp 1688980957
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_335
timestamp 1688980957
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_337
timestamp 1688980957
transform 1 0 32108 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_349
timestamp 1688980957
transform 1 0 33212 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_361
timestamp 1688980957
transform 1 0 34316 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_373
timestamp 1688980957
transform 1 0 35420 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_385
timestamp 1688980957
transform 1 0 36524 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_391
timestamp 1688980957
transform 1 0 37076 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_393
timestamp 1688980957
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_405
timestamp 1688980957
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_417
timestamp 1688980957
transform 1 0 39468 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_429
timestamp 1688980957
transform 1 0 40572 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_441
timestamp 1688980957
transform 1 0 41676 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_447
timestamp 1688980957
transform 1 0 42228 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_449
timestamp 1688980957
transform 1 0 42412 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_461
timestamp 1688980957
transform 1 0 43516 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_473
timestamp 1688980957
transform 1 0 44620 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_485
timestamp 1688980957
transform 1 0 45724 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_497
timestamp 1688980957
transform 1 0 46828 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_503
timestamp 1688980957
transform 1 0 47380 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_505
timestamp 1688980957
transform 1 0 47564 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_517
timestamp 1688980957
transform 1 0 48668 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_529
timestamp 1688980957
transform 1 0 49772 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_541
timestamp 1688980957
transform 1 0 50876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_553
timestamp 1688980957
transform 1 0 51980 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_559
timestamp 1688980957
transform 1 0 52532 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_561
timestamp 1688980957
transform 1 0 52716 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_573
timestamp 1688980957
transform 1 0 53820 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_585
timestamp 1688980957
transform 1 0 54924 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_597
timestamp 1688980957
transform 1 0 56028 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_609
timestamp 1688980957
transform 1 0 57132 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_615
timestamp 1688980957
transform 1 0 57684 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_617
timestamp 1688980957
transform 1 0 57868 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_629
timestamp 1688980957
transform 1 0 58972 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_641
timestamp 1688980957
transform 1 0 60076 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_653
timestamp 1688980957
transform 1 0 61180 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_665
timestamp 1688980957
transform 1 0 62284 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_671
timestamp 1688980957
transform 1 0 62836 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_673
timestamp 1688980957
transform 1 0 63020 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_685
timestamp 1688980957
transform 1 0 64124 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_697
timestamp 1688980957
transform 1 0 65228 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_709
timestamp 1688980957
transform 1 0 66332 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_721
timestamp 1688980957
transform 1 0 67436 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_727
timestamp 1688980957
transform 1 0 67988 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_729
timestamp 1688980957
transform 1 0 68172 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_3
timestamp 1688980957
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_15
timestamp 1688980957
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_27
timestamp 1688980957
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_29
timestamp 1688980957
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_41
timestamp 1688980957
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_53
timestamp 1688980957
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_65
timestamp 1688980957
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_77
timestamp 1688980957
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_83
timestamp 1688980957
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_85
timestamp 1688980957
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_97
timestamp 1688980957
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_109
timestamp 1688980957
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_121
timestamp 1688980957
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_133
timestamp 1688980957
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_139
timestamp 1688980957
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_141
timestamp 1688980957
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_153
timestamp 1688980957
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_165
timestamp 1688980957
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_177
timestamp 1688980957
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_189
timestamp 1688980957
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_195
timestamp 1688980957
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_197
timestamp 1688980957
transform 1 0 19228 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_209
timestamp 1688980957
transform 1 0 20332 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_221
timestamp 1688980957
transform 1 0 21436 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_233
timestamp 1688980957
transform 1 0 22540 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_245
timestamp 1688980957
transform 1 0 23644 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_251
timestamp 1688980957
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_253
timestamp 1688980957
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_265
timestamp 1688980957
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_277
timestamp 1688980957
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_289
timestamp 1688980957
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_301
timestamp 1688980957
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_307
timestamp 1688980957
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_309
timestamp 1688980957
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_321
timestamp 1688980957
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_333
timestamp 1688980957
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_345
timestamp 1688980957
transform 1 0 32844 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_357
timestamp 1688980957
transform 1 0 33948 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_363
timestamp 1688980957
transform 1 0 34500 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_365
timestamp 1688980957
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_377
timestamp 1688980957
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_389
timestamp 1688980957
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_401
timestamp 1688980957
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_413
timestamp 1688980957
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_419
timestamp 1688980957
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_421
timestamp 1688980957
transform 1 0 39836 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_433
timestamp 1688980957
transform 1 0 40940 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_445
timestamp 1688980957
transform 1 0 42044 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_457
timestamp 1688980957
transform 1 0 43148 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_469
timestamp 1688980957
transform 1 0 44252 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_475
timestamp 1688980957
transform 1 0 44804 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_477
timestamp 1688980957
transform 1 0 44988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_489
timestamp 1688980957
transform 1 0 46092 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_501
timestamp 1688980957
transform 1 0 47196 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_513
timestamp 1688980957
transform 1 0 48300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_525
timestamp 1688980957
transform 1 0 49404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_531
timestamp 1688980957
transform 1 0 49956 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_533
timestamp 1688980957
transform 1 0 50140 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_545
timestamp 1688980957
transform 1 0 51244 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_557
timestamp 1688980957
transform 1 0 52348 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_569
timestamp 1688980957
transform 1 0 53452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_581
timestamp 1688980957
transform 1 0 54556 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_587
timestamp 1688980957
transform 1 0 55108 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_589
timestamp 1688980957
transform 1 0 55292 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_601
timestamp 1688980957
transform 1 0 56396 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_613
timestamp 1688980957
transform 1 0 57500 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_625
timestamp 1688980957
transform 1 0 58604 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_637
timestamp 1688980957
transform 1 0 59708 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_643
timestamp 1688980957
transform 1 0 60260 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_645
timestamp 1688980957
transform 1 0 60444 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_657
timestamp 1688980957
transform 1 0 61548 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_669
timestamp 1688980957
transform 1 0 62652 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_681
timestamp 1688980957
transform 1 0 63756 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_693
timestamp 1688980957
transform 1 0 64860 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_699
timestamp 1688980957
transform 1 0 65412 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_701
timestamp 1688980957
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_713
timestamp 1688980957
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_725
timestamp 1688980957
transform 1 0 67804 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_6
timestamp 1688980957
transform 1 0 1656 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_18
timestamp 1688980957
transform 1 0 2760 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_30
timestamp 1688980957
transform 1 0 3864 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_42
timestamp 1688980957
transform 1 0 4968 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115_54
timestamp 1688980957
transform 1 0 6072 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_57
timestamp 1688980957
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_69
timestamp 1688980957
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_81
timestamp 1688980957
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_93
timestamp 1688980957
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_105
timestamp 1688980957
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_111
timestamp 1688980957
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_113
timestamp 1688980957
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_125
timestamp 1688980957
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_137
timestamp 1688980957
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_149
timestamp 1688980957
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_161
timestamp 1688980957
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_167
timestamp 1688980957
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_169
timestamp 1688980957
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_181
timestamp 1688980957
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_193
timestamp 1688980957
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_205
timestamp 1688980957
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_217
timestamp 1688980957
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_223
timestamp 1688980957
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_225
timestamp 1688980957
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_237
timestamp 1688980957
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_249
timestamp 1688980957
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_261
timestamp 1688980957
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_273
timestamp 1688980957
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_279
timestamp 1688980957
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_281
timestamp 1688980957
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_293
timestamp 1688980957
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_305
timestamp 1688980957
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_317
timestamp 1688980957
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_329
timestamp 1688980957
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_335
timestamp 1688980957
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_337
timestamp 1688980957
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_349
timestamp 1688980957
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_361
timestamp 1688980957
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_373
timestamp 1688980957
transform 1 0 35420 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_385
timestamp 1688980957
transform 1 0 36524 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_391
timestamp 1688980957
transform 1 0 37076 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_393
timestamp 1688980957
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_405
timestamp 1688980957
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_417
timestamp 1688980957
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_429
timestamp 1688980957
transform 1 0 40572 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_441
timestamp 1688980957
transform 1 0 41676 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_447
timestamp 1688980957
transform 1 0 42228 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_449
timestamp 1688980957
transform 1 0 42412 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_461
timestamp 1688980957
transform 1 0 43516 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_473
timestamp 1688980957
transform 1 0 44620 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_485
timestamp 1688980957
transform 1 0 45724 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_497
timestamp 1688980957
transform 1 0 46828 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_503
timestamp 1688980957
transform 1 0 47380 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_505
timestamp 1688980957
transform 1 0 47564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_517
timestamp 1688980957
transform 1 0 48668 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_529
timestamp 1688980957
transform 1 0 49772 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_541
timestamp 1688980957
transform 1 0 50876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_553
timestamp 1688980957
transform 1 0 51980 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_559
timestamp 1688980957
transform 1 0 52532 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_561
timestamp 1688980957
transform 1 0 52716 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_573
timestamp 1688980957
transform 1 0 53820 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_585
timestamp 1688980957
transform 1 0 54924 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_597
timestamp 1688980957
transform 1 0 56028 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_609
timestamp 1688980957
transform 1 0 57132 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_615
timestamp 1688980957
transform 1 0 57684 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_617
timestamp 1688980957
transform 1 0 57868 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_629
timestamp 1688980957
transform 1 0 58972 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_641
timestamp 1688980957
transform 1 0 60076 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_653
timestamp 1688980957
transform 1 0 61180 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_665
timestamp 1688980957
transform 1 0 62284 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_671
timestamp 1688980957
transform 1 0 62836 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_673
timestamp 1688980957
transform 1 0 63020 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_685
timestamp 1688980957
transform 1 0 64124 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_697
timestamp 1688980957
transform 1 0 65228 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_709
timestamp 1688980957
transform 1 0 66332 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_721
timestamp 1688980957
transform 1 0 67436 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_727
timestamp 1688980957
transform 1 0 67988 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_729
timestamp 1688980957
transform 1 0 68172 0 -1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_3
timestamp 1688980957
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_15
timestamp 1688980957
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_27
timestamp 1688980957
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_29
timestamp 1688980957
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_41
timestamp 1688980957
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_53
timestamp 1688980957
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_65
timestamp 1688980957
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_77
timestamp 1688980957
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_83
timestamp 1688980957
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_85
timestamp 1688980957
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_97
timestamp 1688980957
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_109
timestamp 1688980957
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_121
timestamp 1688980957
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_133
timestamp 1688980957
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_139
timestamp 1688980957
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_141
timestamp 1688980957
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_153
timestamp 1688980957
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_165
timestamp 1688980957
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_177
timestamp 1688980957
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_189
timestamp 1688980957
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_195
timestamp 1688980957
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_197
timestamp 1688980957
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_209
timestamp 1688980957
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_221
timestamp 1688980957
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_233
timestamp 1688980957
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_245
timestamp 1688980957
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_251
timestamp 1688980957
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_253
timestamp 1688980957
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_265
timestamp 1688980957
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_277
timestamp 1688980957
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_289
timestamp 1688980957
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_301
timestamp 1688980957
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_307
timestamp 1688980957
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_309
timestamp 1688980957
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_321
timestamp 1688980957
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_333
timestamp 1688980957
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_345
timestamp 1688980957
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_357
timestamp 1688980957
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_363
timestamp 1688980957
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_365
timestamp 1688980957
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_377
timestamp 1688980957
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_389
timestamp 1688980957
transform 1 0 36892 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_401
timestamp 1688980957
transform 1 0 37996 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_413
timestamp 1688980957
transform 1 0 39100 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_419
timestamp 1688980957
transform 1 0 39652 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_421
timestamp 1688980957
transform 1 0 39836 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_433
timestamp 1688980957
transform 1 0 40940 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_445
timestamp 1688980957
transform 1 0 42044 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_457
timestamp 1688980957
transform 1 0 43148 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_469
timestamp 1688980957
transform 1 0 44252 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_475
timestamp 1688980957
transform 1 0 44804 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_477
timestamp 1688980957
transform 1 0 44988 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_489
timestamp 1688980957
transform 1 0 46092 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_501
timestamp 1688980957
transform 1 0 47196 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_513
timestamp 1688980957
transform 1 0 48300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_525
timestamp 1688980957
transform 1 0 49404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_531
timestamp 1688980957
transform 1 0 49956 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_533
timestamp 1688980957
transform 1 0 50140 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_545
timestamp 1688980957
transform 1 0 51244 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_557
timestamp 1688980957
transform 1 0 52348 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_569
timestamp 1688980957
transform 1 0 53452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_581
timestamp 1688980957
transform 1 0 54556 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_587
timestamp 1688980957
transform 1 0 55108 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_589
timestamp 1688980957
transform 1 0 55292 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_601
timestamp 1688980957
transform 1 0 56396 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_613
timestamp 1688980957
transform 1 0 57500 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_625
timestamp 1688980957
transform 1 0 58604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_637
timestamp 1688980957
transform 1 0 59708 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_643
timestamp 1688980957
transform 1 0 60260 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_645
timestamp 1688980957
transform 1 0 60444 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_657
timestamp 1688980957
transform 1 0 61548 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_669
timestamp 1688980957
transform 1 0 62652 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_681
timestamp 1688980957
transform 1 0 63756 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_693
timestamp 1688980957
transform 1 0 64860 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_699
timestamp 1688980957
transform 1 0 65412 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_701
timestamp 1688980957
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_713
timestamp 1688980957
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_725
timestamp 1688980957
transform 1 0 67804 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_3
timestamp 1688980957
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_15
timestamp 1688980957
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_27
timestamp 1688980957
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_39
timestamp 1688980957
transform 1 0 4692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_51
timestamp 1688980957
transform 1 0 5796 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_55
timestamp 1688980957
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_57
timestamp 1688980957
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_69
timestamp 1688980957
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_81
timestamp 1688980957
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_93
timestamp 1688980957
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_105
timestamp 1688980957
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_111
timestamp 1688980957
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_113
timestamp 1688980957
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_125
timestamp 1688980957
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_137
timestamp 1688980957
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_149
timestamp 1688980957
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_161
timestamp 1688980957
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_167
timestamp 1688980957
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_169
timestamp 1688980957
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_181
timestamp 1688980957
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_193
timestamp 1688980957
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_205
timestamp 1688980957
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_217
timestamp 1688980957
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_223
timestamp 1688980957
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_225
timestamp 1688980957
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_237
timestamp 1688980957
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_249
timestamp 1688980957
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_261
timestamp 1688980957
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_273
timestamp 1688980957
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_279
timestamp 1688980957
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_281
timestamp 1688980957
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_293
timestamp 1688980957
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_305
timestamp 1688980957
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_317
timestamp 1688980957
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_329
timestamp 1688980957
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_335
timestamp 1688980957
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_337
timestamp 1688980957
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_349
timestamp 1688980957
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_361
timestamp 1688980957
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_373
timestamp 1688980957
transform 1 0 35420 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_385
timestamp 1688980957
transform 1 0 36524 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_391
timestamp 1688980957
transform 1 0 37076 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_393
timestamp 1688980957
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_405
timestamp 1688980957
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_417
timestamp 1688980957
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_429
timestamp 1688980957
transform 1 0 40572 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_441
timestamp 1688980957
transform 1 0 41676 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_447
timestamp 1688980957
transform 1 0 42228 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_449
timestamp 1688980957
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_461
timestamp 1688980957
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_473
timestamp 1688980957
transform 1 0 44620 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_485
timestamp 1688980957
transform 1 0 45724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_497
timestamp 1688980957
transform 1 0 46828 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_503
timestamp 1688980957
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_505
timestamp 1688980957
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_517
timestamp 1688980957
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_529
timestamp 1688980957
transform 1 0 49772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_541
timestamp 1688980957
transform 1 0 50876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_553
timestamp 1688980957
transform 1 0 51980 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_559
timestamp 1688980957
transform 1 0 52532 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_561
timestamp 1688980957
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_573
timestamp 1688980957
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_585
timestamp 1688980957
transform 1 0 54924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_597
timestamp 1688980957
transform 1 0 56028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_609
timestamp 1688980957
transform 1 0 57132 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_615
timestamp 1688980957
transform 1 0 57684 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_617
timestamp 1688980957
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_629
timestamp 1688980957
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_641
timestamp 1688980957
transform 1 0 60076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_653
timestamp 1688980957
transform 1 0 61180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_665
timestamp 1688980957
transform 1 0 62284 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_671
timestamp 1688980957
transform 1 0 62836 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_673
timestamp 1688980957
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_685
timestamp 1688980957
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_697
timestamp 1688980957
transform 1 0 65228 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_709
timestamp 1688980957
transform 1 0 66332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_721
timestamp 1688980957
transform 1 0 67436 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_727
timestamp 1688980957
transform 1 0 67988 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_729
timestamp 1688980957
transform 1 0 68172 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_3
timestamp 1688980957
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_15
timestamp 1688980957
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_27
timestamp 1688980957
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_29
timestamp 1688980957
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_41
timestamp 1688980957
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_53
timestamp 1688980957
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_65
timestamp 1688980957
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_77
timestamp 1688980957
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_83
timestamp 1688980957
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_85
timestamp 1688980957
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_97
timestamp 1688980957
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_109
timestamp 1688980957
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_121
timestamp 1688980957
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_133
timestamp 1688980957
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_139
timestamp 1688980957
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_141
timestamp 1688980957
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_153
timestamp 1688980957
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_165
timestamp 1688980957
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_177
timestamp 1688980957
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_189
timestamp 1688980957
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_195
timestamp 1688980957
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_197
timestamp 1688980957
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_209
timestamp 1688980957
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_221
timestamp 1688980957
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_233
timestamp 1688980957
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_245
timestamp 1688980957
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_251
timestamp 1688980957
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_253
timestamp 1688980957
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_265
timestamp 1688980957
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_277
timestamp 1688980957
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_289
timestamp 1688980957
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_301
timestamp 1688980957
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_307
timestamp 1688980957
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_309
timestamp 1688980957
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_321
timestamp 1688980957
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_333
timestamp 1688980957
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_345
timestamp 1688980957
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_357
timestamp 1688980957
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_363
timestamp 1688980957
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_365
timestamp 1688980957
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_377
timestamp 1688980957
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_389
timestamp 1688980957
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_401
timestamp 1688980957
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_413
timestamp 1688980957
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_419
timestamp 1688980957
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_421
timestamp 1688980957
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_433
timestamp 1688980957
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_445
timestamp 1688980957
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_457
timestamp 1688980957
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_469
timestamp 1688980957
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_475
timestamp 1688980957
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_477
timestamp 1688980957
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_489
timestamp 1688980957
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_501
timestamp 1688980957
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_513
timestamp 1688980957
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_525
timestamp 1688980957
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_531
timestamp 1688980957
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_533
timestamp 1688980957
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_545
timestamp 1688980957
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_557
timestamp 1688980957
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_569
timestamp 1688980957
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_581
timestamp 1688980957
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_587
timestamp 1688980957
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_589
timestamp 1688980957
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_601
timestamp 1688980957
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_613
timestamp 1688980957
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_625
timestamp 1688980957
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_637
timestamp 1688980957
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_643
timestamp 1688980957
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_645
timestamp 1688980957
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_657
timestamp 1688980957
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_669
timestamp 1688980957
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_681
timestamp 1688980957
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_693
timestamp 1688980957
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_699
timestamp 1688980957
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_701
timestamp 1688980957
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_713
timestamp 1688980957
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_725
timestamp 1688980957
transform 1 0 67804 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_3
timestamp 1688980957
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_15
timestamp 1688980957
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_27
timestamp 1688980957
transform 1 0 3588 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_29
timestamp 1688980957
transform 1 0 3772 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_41
timestamp 1688980957
transform 1 0 4876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_53
timestamp 1688980957
transform 1 0 5980 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_57
timestamp 1688980957
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_69
timestamp 1688980957
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_81
timestamp 1688980957
transform 1 0 8556 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_85
timestamp 1688980957
transform 1 0 8924 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_97
timestamp 1688980957
transform 1 0 10028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_109
timestamp 1688980957
transform 1 0 11132 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_113
timestamp 1688980957
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_125
timestamp 1688980957
transform 1 0 12604 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_132
timestamp 1688980957
transform 1 0 13248 0 -1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_141
timestamp 1688980957
transform 1 0 14076 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_153
timestamp 1688980957
transform 1 0 15180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_165
timestamp 1688980957
transform 1 0 16284 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_169
timestamp 1688980957
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_181
timestamp 1688980957
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_193
timestamp 1688980957
transform 1 0 18860 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_197
timestamp 1688980957
transform 1 0 19228 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_209
timestamp 1688980957
transform 1 0 20332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_221
timestamp 1688980957
transform 1 0 21436 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_225
timestamp 1688980957
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_237
timestamp 1688980957
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_249
timestamp 1688980957
transform 1 0 24012 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_253
timestamp 1688980957
transform 1 0 24380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_265
timestamp 1688980957
transform 1 0 25484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_277
timestamp 1688980957
transform 1 0 26588 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_281
timestamp 1688980957
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_293
timestamp 1688980957
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_305
timestamp 1688980957
transform 1 0 29164 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_309
timestamp 1688980957
transform 1 0 29532 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_317
timestamp 1688980957
transform 1 0 30268 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_321
timestamp 1688980957
transform 1 0 30636 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_333
timestamp 1688980957
transform 1 0 31740 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_337
timestamp 1688980957
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_349
timestamp 1688980957
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_361
timestamp 1688980957
transform 1 0 34316 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_365
timestamp 1688980957
transform 1 0 34684 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_377
timestamp 1688980957
transform 1 0 35788 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_389
timestamp 1688980957
transform 1 0 36892 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_393
timestamp 1688980957
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_405
timestamp 1688980957
transform 1 0 38364 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_413
timestamp 1688980957
transform 1 0 39100 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_419
timestamp 1688980957
transform 1 0 39652 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_421
timestamp 1688980957
transform 1 0 39836 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_433
timestamp 1688980957
transform 1 0 40940 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_445
timestamp 1688980957
transform 1 0 42044 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_449
timestamp 1688980957
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_461
timestamp 1688980957
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_473
timestamp 1688980957
transform 1 0 44620 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_477
timestamp 1688980957
transform 1 0 44988 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_489
timestamp 1688980957
transform 1 0 46092 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_501
timestamp 1688980957
transform 1 0 47196 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_505
timestamp 1688980957
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_517
timestamp 1688980957
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_529
timestamp 1688980957
transform 1 0 49772 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_533
timestamp 1688980957
transform 1 0 50140 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_545
timestamp 1688980957
transform 1 0 51244 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_557
timestamp 1688980957
transform 1 0 52348 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_561
timestamp 1688980957
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_573
timestamp 1688980957
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_585
timestamp 1688980957
transform 1 0 54924 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_589
timestamp 1688980957
transform 1 0 55292 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_601
timestamp 1688980957
transform 1 0 56396 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_613
timestamp 1688980957
transform 1 0 57500 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_617
timestamp 1688980957
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_629
timestamp 1688980957
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_641
timestamp 1688980957
transform 1 0 60076 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_645
timestamp 1688980957
transform 1 0 60444 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_657
timestamp 1688980957
transform 1 0 61548 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_669
timestamp 1688980957
transform 1 0 62652 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_673
timestamp 1688980957
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_685
timestamp 1688980957
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_697
timestamp 1688980957
transform 1 0 65228 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_701
timestamp 1688980957
transform 1 0 65596 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_713
timestamp 1688980957
transform 1 0 66700 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119_725
timestamp 1688980957
transform 1 0 67804 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_729
timestamp 1688980957
transform 1 0 68172 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32936 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 21344 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 17388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 17388 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 31740 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 27692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 26772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 21436 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 21620 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 11500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 26588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 26404 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 17664 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 28980 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 23644 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 19044 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 15456 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 38824 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 20700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 37996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 37168 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 17572 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold31 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22264 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 29440 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 28428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 30728 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 27968 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 27876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 13984 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 16928 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 26404 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 23276 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 22080 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 33396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 18676 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 38640 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 30268 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold48
timestamp 1688980957
transform -1 0 25576 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 24748 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 16100 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 16560 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 33856 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 36616 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform -1 0 37352 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 12880 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 24840 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 24288 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 22540 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform -1 0 34776 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 34040 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 35972 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 30268 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 28612 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 21252 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 27968 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 30544 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 31740 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform -1 0 28888 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 30268 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform -1 0 33948 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform -1 0 17664 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 37996 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 24564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 30268 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 20332 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 22632 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 26956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 27784 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 16744 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 15916 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 35236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 35420 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 16192 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 36892 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 37168 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 30268 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 28520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 20608 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 38640 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 37168 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 36708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform -1 0 16560 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 16008 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 21344 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 19228 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform -1 0 33672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform -1 0 34408 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold102 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform -1 0 27968 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform -1 0 27140 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform -1 0 26864 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 13064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 19136 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 29624 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 33580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 32844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform -1 0 28980 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform -1 0 37996 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform -1 0 36432 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform -1 0 31004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 34776 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 23092 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 23184 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 29900 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 32384 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform 1 0 17020 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 18860 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 16192 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 24104 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform 1 0 22356 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 35420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform -1 0 25576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform -1 0 27692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform -1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 17296 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 13984 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform 1 0 9936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 13984 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform -1 0 24288 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 25300 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform -1 0 10212 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform 1 0 16744 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform -1 0 10948 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 10304 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 21528 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform -1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 17480 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform -1 0 10856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform -1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform 1 0 16744 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 21712 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform -1 0 25392 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform -1 0 37168 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform -1 0 68540 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output3
timestamp 1688980957
transform 1 0 67528 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1688980957
transform -1 0 1932 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1688980957
transform 1 0 43884 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1688980957
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1688980957
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1688980957
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1688980957
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1688980957
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1688980957
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1688980957
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1688980957
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1688980957
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1688980957
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1688980957
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1688980957
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1688980957
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1688980957
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1688980957
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1688980957
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1688980957
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1688980957
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1688980957
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1688980957
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1688980957
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1688980957
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1688980957
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1688980957
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1688980957
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1688980957
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1688980957
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1688980957
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1688980957
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1688980957
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1688980957
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1688980957
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1688980957
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1688980957
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1688980957
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1688980957
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1688980957
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1688980957
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1688980957
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1688980957
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1688980957
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1688980957
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1688980957
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1688980957
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1688980957
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1688980957
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1688980957
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1688980957
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1688980957
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1688980957
transform -1 0 68816 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1688980957
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1688980957
transform -1 0 68816 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1688980957
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1688980957
transform -1 0 68816 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1688980957
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1688980957
transform -1 0 68816 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1688980957
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1688980957
transform -1 0 68816 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1688980957
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1688980957
transform -1 0 68816 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1688980957
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1688980957
transform -1 0 68816 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1688980957
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1688980957
transform -1 0 68816 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1688980957
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1688980957
transform -1 0 68816 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1688980957
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1688980957
transform -1 0 68816 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1688980957
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1688980957
transform -1 0 68816 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1688980957
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1688980957
transform -1 0 68816 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1688980957
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1688980957
transform -1 0 68816 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1688980957
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1688980957
transform -1 0 68816 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1688980957
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1688980957
transform -1 0 68816 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1688980957
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1688980957
transform -1 0 68816 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1688980957
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1688980957
transform -1 0 68816 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1688980957
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1688980957
transform -1 0 68816 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1688980957
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1688980957
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1688980957
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1688980957
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1688980957
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1688980957
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1688980957
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1688980957
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1688980957
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1688980957
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1688980957
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1688980957
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1688980957
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1688980957
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1688980957
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1688980957
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1688980957
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1688980957
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1688980957
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1688980957
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1688980957
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1688980957
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1688980957
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1688980957
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1688980957
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1688980957
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1688980957
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1688980957
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1688980957
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1688980957
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1688980957
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1688980957
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1688980957
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1688980957
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1688980957
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1688980957
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1688980957
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1688980957
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1688980957
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1688980957
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1688980957
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1688980957
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1688980957
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1688980957
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1688980957
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1688980957
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1688980957
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1688980957
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1688980957
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1688980957
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1688980957
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1688980957
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1688980957
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1688980957
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1688980957
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1688980957
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1688980957
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1688980957
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1688980957
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1688980957
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1688980957
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1688980957
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1688980957
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1688980957
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1688980957
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1688980957
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1688980957
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1688980957
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1688980957
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1688980957
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1688980957
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1688980957
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1688980957
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1688980957
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1688980957
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1688980957
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1688980957
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1688980957
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1688980957
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1688980957
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1688980957
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1688980957
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1688980957
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1688980957
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1688980957
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1688980957
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1688980957
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1688980957
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1688980957
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1688980957
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1688980957
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1688980957
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1688980957
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1688980957
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1688980957
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1688980957
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1688980957
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1688980957
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1688980957
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1688980957
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1688980957
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1688980957
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1688980957
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1688980957
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1688980957
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1688980957
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1688980957
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1688980957
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1688980957
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1688980957
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1688980957
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1688980957
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1688980957
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1688980957
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1688980957
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1688980957
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1688980957
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1688980957
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1688980957
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1688980957
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1688980957
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1688980957
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1688980957
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1688980957
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1688980957
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1688980957
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1688980957
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1688980957
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1688980957
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1688980957
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1688980957
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1688980957
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1688980957
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1688980957
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1688980957
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1688980957
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1688980957
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1688980957
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1688980957
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1688980957
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1688980957
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1688980957
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1688980957
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1688980957
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1688980957
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1688980957
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1688980957
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1688980957
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1688980957
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1688980957
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1688980957
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1688980957
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1688980957
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1688980957
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1688980957
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1688980957
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1688980957
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1688980957
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1688980957
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1688980957
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1688980957
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1688980957
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1688980957
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1688980957
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1688980957
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1688980957
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1688980957
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1688980957
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1688980957
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1688980957
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1688980957
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1688980957
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1688980957
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1688980957
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1688980957
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1688980957
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1688980957
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1688980957
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1688980957
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1688980957
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1688980957
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1688980957
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1688980957
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1688980957
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1688980957
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1688980957
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1688980957
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1688980957
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1688980957
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1688980957
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1688980957
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1688980957
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1688980957
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1688980957
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1688980957
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1688980957
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1688980957
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1688980957
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1688980957
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1688980957
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1688980957
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1688980957
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1688980957
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1688980957
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1688980957
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1688980957
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1688980957
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1688980957
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1688980957
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1688980957
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1688980957
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1688980957
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1688980957
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1688980957
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1688980957
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1688980957
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1688980957
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1688980957
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1688980957
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1688980957
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1688980957
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1688980957
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1688980957
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1688980957
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1688980957
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1688980957
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1688980957
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1688980957
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1688980957
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1688980957
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1688980957
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1688980957
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1688980957
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1688980957
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1688980957
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1688980957
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1688980957
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1688980957
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1688980957
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1688980957
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1688980957
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1688980957
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1688980957
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1688980957
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1688980957
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1688980957
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1688980957
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1688980957
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1688980957
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1688980957
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1688980957
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1688980957
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1688980957
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1688980957
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1688980957
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1688980957
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1688980957
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1688980957
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1688980957
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1688980957
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1688980957
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1688980957
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1688980957
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1688980957
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1688980957
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1688980957
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1688980957
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1688980957
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1688980957
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1688980957
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1688980957
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1688980957
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1688980957
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1688980957
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1688980957
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1688980957
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1688980957
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1688980957
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1688980957
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1688980957
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1688980957
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1688980957
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1688980957
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1688980957
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1688980957
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1688980957
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1688980957
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1688980957
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1688980957
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1688980957
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1688980957
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1688980957
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1688980957
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1688980957
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1688980957
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1688980957
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1688980957
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1688980957
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1688980957
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1688980957
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1688980957
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1688980957
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1688980957
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1688980957
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1688980957
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1688980957
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1688980957
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1688980957
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1688980957
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1688980957
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1688980957
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1688980957
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1688980957
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1688980957
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1688980957
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1688980957
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1688980957
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1688980957
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1688980957
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1688980957
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1688980957
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1688980957
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1688980957
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1688980957
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1688980957
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1688980957
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1688980957
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1688980957
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1688980957
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1688980957
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1688980957
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1688980957
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1688980957
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1688980957
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1688980957
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1688980957
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1688980957
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1688980957
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1688980957
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1688980957
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1688980957
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1688980957
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1688980957
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1688980957
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1688980957
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1688980957
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1688980957
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1688980957
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1688980957
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1688980957
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1688980957
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1688980957
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1688980957
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1688980957
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1688980957
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1688980957
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1688980957
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1688980957
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1688980957
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1688980957
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1688980957
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1688980957
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1688980957
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1688980957
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1688980957
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1688980957
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1688980957
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1688980957
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1688980957
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1688980957
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1688980957
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1688980957
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1688980957
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1688980957
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1688980957
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1688980957
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1688980957
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1688980957
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1688980957
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1688980957
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1688980957
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1688980957
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1688980957
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1688980957
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1688980957
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1688980957
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1688980957
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1688980957
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1688980957
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1688980957
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1688980957
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1688980957
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1688980957
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1688980957
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1688980957
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1688980957
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1688980957
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1688980957
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1688980957
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1688980957
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1688980957
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1688980957
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1688980957
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1688980957
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1688980957
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1688980957
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1688980957
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1688980957
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1688980957
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1688980957
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1688980957
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1688980957
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1688980957
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1688980957
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1688980957
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1688980957
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1688980957
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1688980957
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1688980957
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1688980957
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1688980957
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1688980957
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1688980957
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1688980957
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1688980957
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1688980957
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1688980957
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1688980957
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1688980957
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1688980957
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1688980957
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1688980957
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1688980957
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1688980957
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1688980957
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1688980957
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1688980957
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1688980957
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1688980957
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1688980957
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1688980957
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1688980957
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1688980957
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1688980957
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1688980957
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1688980957
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1688980957
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1688980957
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1688980957
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1688980957
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1688980957
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1688980957
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1688980957
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1688980957
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1688980957
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1688980957
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1688980957
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1688980957
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1688980957
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1688980957
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1688980957
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1688980957
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1688980957
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1688980957
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1688980957
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1688980957
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1688980957
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1688980957
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1688980957
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1688980957
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1688980957
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1688980957
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1688980957
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1688980957
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1688980957
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1688980957
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1688980957
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1688980957
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1688980957
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1688980957
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1688980957
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1688980957
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1688980957
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1688980957
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1688980957
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1688980957
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1688980957
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1688980957
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1688980957
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1688980957
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1688980957
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1688980957
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1688980957
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1688980957
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1688980957
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1688980957
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1688980957
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1688980957
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1688980957
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1688980957
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1688980957
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1688980957
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1688980957
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1688980957
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1688980957
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1688980957
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1688980957
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1688980957
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1688980957
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1688980957
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1688980957
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1688980957
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1688980957
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1688980957
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1688980957
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1688980957
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1688980957
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1688980957
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1688980957
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1688980957
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1688980957
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1688980957
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1688980957
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1688980957
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1688980957
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1688980957
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1688980957
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1688980957
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1688980957
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1688980957
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1688980957
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1688980957
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1688980957
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1688980957
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1688980957
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1688980957
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1688980957
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1688980957
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1688980957
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1688980957
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1688980957
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1688980957
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1688980957
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1688980957
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1688980957
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1688980957
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1688980957
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1688980957
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1688980957
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1688980957
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1688980957
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1688980957
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1688980957
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1688980957
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1688980957
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1688980957
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1688980957
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1688980957
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1688980957
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1688980957
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1688980957
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1688980957
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1688980957
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1688980957
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1688980957
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1688980957
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1688980957
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1688980957
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1688980957
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1688980957
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1688980957
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1688980957
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1688980957
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1688980957
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1688980957
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1688980957
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1688980957
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1688980957
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1688980957
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1688980957
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1688980957
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1688980957
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1688980957
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1688980957
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1688980957
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1688980957
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1688980957
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1688980957
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1688980957
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1688980957
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1688980957
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1688980957
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1688980957
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1688980957
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1688980957
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1688980957
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1688980957
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1688980957
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1688980957
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1688980957
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1688980957
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1688980957
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1688980957
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1688980957
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1688980957
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1688980957
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1688980957
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1688980957
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1688980957
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1688980957
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1688980957
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1688980957
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1688980957
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1688980957
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1688980957
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1688980957
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1688980957
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1688980957
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1688980957
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1688980957
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1688980957
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1688980957
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1688980957
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1688980957
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1688980957
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1688980957
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1688980957
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1688980957
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1688980957
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1688980957
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1688980957
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1688980957
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1688980957
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1688980957
transform 1 0 60352 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1688980957
transform 1 0 65504 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1688980957
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1688980957
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1688980957
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1688980957
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1688980957
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1688980957
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1688980957
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1688980957
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1688980957
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1688980957
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1688980957
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1688980957
transform 1 0 62928 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1688980957
transform 1 0 68080 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1688980957
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1688980957
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1688980957
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1688980957
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1688980957
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1688980957
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1688980957
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1688980957
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1688980957
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1688980957
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1688980957
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1688980957
transform 1 0 60352 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1688980957
transform 1 0 65504 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1688980957
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1688980957
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1688980957
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1688980957
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1688980957
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1688980957
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1688980957
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1688980957
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1688980957
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1688980957
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1688980957
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1688980957
transform 1 0 62928 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1688980957
transform 1 0 68080 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1688980957
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1688980957
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1688980957
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1688980957
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1688980957
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1688980957
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1688980957
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1688980957
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1688980957
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1688980957
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1688980957
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1688980957
transform 1 0 60352 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1688980957
transform 1 0 65504 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1688980957
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1688980957
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1688980957
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1688980957
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1688980957
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1688980957
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1688980957
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1688980957
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1688980957
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1688980957
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1688980957
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1688980957
transform 1 0 62928 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1688980957
transform 1 0 68080 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1688980957
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1688980957
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1688980957
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1688980957
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1688980957
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1688980957
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1688980957
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1688980957
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1688980957
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1688980957
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1688980957
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1688980957
transform 1 0 60352 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1688980957
transform 1 0 65504 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1688980957
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1688980957
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1688980957
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1688980957
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1688980957
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1688980957
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1688980957
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1688980957
transform 1 0 42320 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1688980957
transform 1 0 47472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1688980957
transform 1 0 52624 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1688980957
transform 1 0 57776 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1688980957
transform 1 0 62928 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1688980957
transform 1 0 68080 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1688980957
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1688980957
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1688980957
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1688980957
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1688980957
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1688980957
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1688980957
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1688980957
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1688980957
transform 1 0 44896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1688980957
transform 1 0 50048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1688980957
transform 1 0 55200 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1688980957
transform 1 0 60352 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1688980957
transform 1 0 65504 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1688980957
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1688980957
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1688980957
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1688980957
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1688980957
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1688980957
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1688980957
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1688980957
transform 1 0 42320 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1688980957
transform 1 0 47472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1688980957
transform 1 0 52624 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1688980957
transform 1 0 57776 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1688980957
transform 1 0 62928 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1688980957
transform 1 0 68080 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1688980957
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1688980957
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1688980957
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1688980957
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1688980957
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1688980957
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1688980957
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1688980957
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1688980957
transform 1 0 44896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1688980957
transform 1 0 50048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1688980957
transform 1 0 55200 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1688980957
transform 1 0 60352 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1688980957
transform 1 0 65504 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1688980957
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1688980957
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1688980957
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1688980957
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1688980957
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1688980957
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1688980957
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1688980957
transform 1 0 42320 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1688980957
transform 1 0 47472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1688980957
transform 1 0 52624 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1688980957
transform 1 0 57776 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1688980957
transform 1 0 62928 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1688980957
transform 1 0 68080 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1688980957
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1688980957
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1688980957
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1688980957
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1688980957
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1688980957
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1688980957
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1688980957
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1688980957
transform 1 0 44896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1688980957
transform 1 0 50048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1688980957
transform 1 0 55200 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1688980957
transform 1 0 60352 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1688980957
transform 1 0 65504 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1688980957
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1688980957
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1688980957
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1688980957
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1688980957
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1688980957
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1688980957
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1688980957
transform 1 0 42320 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1688980957
transform 1 0 47472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1688980957
transform 1 0 52624 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1688980957
transform 1 0 57776 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1688980957
transform 1 0 62928 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1688980957
transform 1 0 68080 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1688980957
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1688980957
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1688980957
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1688980957
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1688980957
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1688980957
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1688980957
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1688980957
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1688980957
transform 1 0 44896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1688980957
transform 1 0 50048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1688980957
transform 1 0 55200 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1688980957
transform 1 0 60352 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1688980957
transform 1 0 65504 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1688980957
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1688980957
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1688980957
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1688980957
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1688980957
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1688980957
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1688980957
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1688980957
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1688980957
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1688980957
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1688980957
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1688980957
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1688980957
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1688980957
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1688980957
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1688980957
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1688980957
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1688980957
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1688980957
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1688980957
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1688980957
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1688980957
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1688980957
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1688980957
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1688980957
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1688980957
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1688980957
transform 1 0 3680 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1688980957
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1688980957
transform 1 0 8832 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1688980957
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1688980957
transform 1 0 13984 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1688980957
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1688980957
transform 1 0 19136 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1688980957
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1688980957
transform 1 0 24288 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1688980957
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1688980957
transform 1 0 29440 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1688980957
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1688980957
transform 1 0 34592 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1688980957
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1688980957
transform 1 0 39744 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1688980957
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1688980957
transform 1 0 44896 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1688980957
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1688980957
transform 1 0 50048 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1688980957
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1688980957
transform 1 0 55200 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1688980957
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1688980957
transform 1 0 60352 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1688980957
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1688980957
transform 1 0 65504 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1688980957
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire6
timestamp 1688980957
transform -1 0 12512 0 1 16320
box -38 -48 314 592
<< labels >>
flabel metal3 s 69200 46248 70000 46368 0 FreeSans 480 0 0 0 audio_sample[0]
port 0 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 audio_sample[10]
port 1 nsew signal input
flabel metal3 s 0 55768 800 55888 0 FreeSans 480 0 0 0 audio_sample[11]
port 2 nsew signal input
flabel metal3 s 69200 37408 70000 37528 0 FreeSans 480 0 0 0 audio_sample[12]
port 3 nsew signal input
flabel metal2 s 47674 69200 47730 70000 0 FreeSans 224 90 0 0 audio_sample[13]
port 4 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 audio_sample[14]
port 5 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 audio_sample[15]
port 6 nsew signal input
flabel metal3 s 69200 65288 70000 65408 0 FreeSans 480 0 0 0 audio_sample[1]
port 7 nsew signal input
flabel metal2 s 56690 69200 56746 70000 0 FreeSans 224 90 0 0 audio_sample[2]
port 8 nsew signal input
flabel metal3 s 69200 18368 70000 18488 0 FreeSans 480 0 0 0 audio_sample[3]
port 9 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 audio_sample[4]
port 10 nsew signal input
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 audio_sample[5]
port 11 nsew signal input
flabel metal2 s 65706 69200 65762 70000 0 FreeSans 224 90 0 0 audio_sample[6]
port 12 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 audio_sample[7]
port 13 nsew signal input
flabel metal2 s 21270 69200 21326 70000 0 FreeSans 224 90 0 0 audio_sample[8]
port 14 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 audio_sample[9]
port 15 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 clk
port 16 nsew signal input
flabel metal3 s 69200 8 70000 128 0 FreeSans 480 0 0 0 done
port 17 nsew signal tristate
flabel metal3 s 0 46248 800 46368 0 FreeSans 480 0 0 0 psram_ce_n
port 18 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 psram_d[0]
port 19 nsew signal bidirectional
flabel metal2 s 12898 69200 12954 70000 0 FreeSans 224 90 0 0 psram_d[1]
port 20 nsew signal bidirectional
flabel metal3 s 69200 9528 70000 9648 0 FreeSans 480 0 0 0 psram_d[2]
port 21 nsew signal bidirectional
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 psram_d[3]
port 22 nsew signal bidirectional
flabel metal3 s 0 64608 800 64728 0 FreeSans 480 0 0 0 psram_douten[0]
port 23 nsew signal tristate
flabel metal3 s 69200 55768 70000 55888 0 FreeSans 480 0 0 0 psram_douten[1]
port 24 nsew signal tristate
flabel metal2 s 30286 69200 30342 70000 0 FreeSans 224 90 0 0 psram_douten[2]
port 25 nsew signal tristate
flabel metal2 s 39302 69200 39358 70000 0 FreeSans 224 90 0 0 psram_douten[3]
port 26 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 psram_sck
port 27 nsew signal tristate
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 rst
port 28 nsew signal input
flabel metal2 s 3882 69200 3938 70000 0 FreeSans 224 90 0 0 sample_valid
port 29 nsew signal input
flabel metal3 s 69200 27888 70000 28008 0 FreeSans 480 0 0 0 start
port 30 nsew signal input
flabel metal4 s 4208 2128 4528 67504 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 34928 2128 35248 67504 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 65648 2128 65968 67504 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 19568 2128 19888 67504 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 67504 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
rlabel via1 34960 66912 34960 66912 0 vccd1
rlabel metal1 34960 67456 34960 67456 0 vssd1
rlabel metal1 18078 16762 18078 16762 0 _0000_
rlabel metal1 17909 17578 17909 17578 0 _0001_
rlabel metal1 19416 21522 19416 21522 0 _0002_
rlabel metal1 16560 24922 16560 24922 0 _0003_
rlabel metal1 24844 19346 24844 19346 0 _0004_
rlabel metal1 24968 20434 24968 20434 0 _0005_
rlabel metal1 22034 15096 22034 15096 0 _0006_
rlabel metal1 18998 15130 18998 15130 0 _0007_
rlabel metal1 25054 16150 25054 16150 0 _0008_
rlabel via1 25433 17646 25433 17646 0 _0009_
rlabel metal2 29394 21284 29394 21284 0 _0010_
rlabel metal2 29486 21794 29486 21794 0 _0011_
rlabel metal1 17802 18326 17802 18326 0 _0012_
rlabel metal1 15364 17306 15364 17306 0 _0013_
rlabel metal1 16882 14586 16882 14586 0 _0014_
rlabel metal1 17802 18394 17802 18394 0 _0015_
rlabel metal2 17710 21692 17710 21692 0 _0016_
rlabel metal1 16652 24378 16652 24378 0 _0017_
rlabel metal2 18538 23970 18538 23970 0 _0018_
rlabel via1 17346 20910 17346 20910 0 _0019_
rlabel metal1 20378 20570 20378 20570 0 _0020_
rlabel metal1 25948 20910 25948 20910 0 _0021_
rlabel metal1 23092 20570 23092 20570 0 _0022_
rlabel metal2 22494 20434 22494 20434 0 _0023_
rlabel metal2 22402 16524 22402 16524 0 _0024_
rlabel metal1 19764 16490 19764 16490 0 _0025_
rlabel metal1 18921 15402 18921 15402 0 _0026_
rlabel metal1 22218 15470 22218 15470 0 _0027_
rlabel metal1 27140 16762 27140 16762 0 _0028_
rlabel metal1 27937 17578 27937 17578 0 _0029_
rlabel metal1 25852 18938 25852 18938 0 _0030_
rlabel metal1 37030 20570 37030 20570 0 _0031_
rlabel metal2 34270 21318 34270 21318 0 _0032_
rlabel metal1 28106 20434 28106 20434 0 _0033_
rlabel metal2 29394 22882 29394 22882 0 _0034_
rlabel metal1 30364 25194 30364 25194 0 _0035_
rlabel metal2 35374 15266 35374 15266 0 _0036_
rlabel metal1 21735 19482 21735 19482 0 _0037_
rlabel metal1 13999 16490 13999 16490 0 _0038_
rlabel metal1 24472 15130 24472 15130 0 _0039_
rlabel metal1 34132 15674 34132 15674 0 _0040_
rlabel metal1 22356 17170 22356 17170 0 _0041_
rlabel metal1 19918 18938 19918 18938 0 _0042_
rlabel metal2 28198 14756 28198 14756 0 _0043_
rlabel metal1 11684 17714 11684 17714 0 _0044_
rlabel metal1 14398 20978 14398 20978 0 _0045_
rlabel metal1 20700 22406 20700 22406 0 _0046_
rlabel metal2 20470 13124 20470 13124 0 _0047_
rlabel metal1 24794 11662 24794 11662 0 _0048_
rlabel metal1 28934 12818 28934 12818 0 _0049_
rlabel metal1 15594 14858 15594 14858 0 _0050_
rlabel metal1 32469 17238 32469 17238 0 _0051_
rlabel metal1 30084 11322 30084 11322 0 _0052_
rlabel metal1 12972 17306 12972 17306 0 _0053_
rlabel metal1 11677 11118 11677 11118 0 _0054_
rlabel metal1 13892 13498 13892 13498 0 _0055_
rlabel metal1 13064 11866 13064 11866 0 _0056_
rlabel metal1 9568 12410 9568 12410 0 _0057_
rlabel metal2 8602 13736 8602 13736 0 _0058_
rlabel metal2 8602 15266 8602 15266 0 _0059_
rlabel metal1 8556 16762 8556 16762 0 _0060_
rlabel metal2 9522 18462 9522 18462 0 _0061_
rlabel metal2 10994 18428 10994 18428 0 _0062_
rlabel metal1 14812 20570 14812 20570 0 _0063_
rlabel metal2 8694 20638 8694 20638 0 _0064_
rlabel metal1 11684 19482 11684 19482 0 _0065_
rlabel metal2 9614 20468 9614 20468 0 _0066_
rlabel metal1 9016 22202 9016 22202 0 _0067_
rlabel metal1 9016 23290 9016 23290 0 _0068_
rlabel metal1 9384 24378 9384 24378 0 _0069_
rlabel metal2 11178 25058 11178 25058 0 _0070_
rlabel metal1 13945 26282 13945 26282 0 _0071_
rlabel metal2 16330 25704 16330 25704 0 _0072_
rlabel metal1 14444 19142 14444 19142 0 _0073_
rlabel metal2 21298 22005 21298 22005 0 _0074_
rlabel metal2 21114 28696 21114 28696 0 _0075_
rlabel metal1 24656 29002 24656 29002 0 _0076_
rlabel metal2 24886 28526 24886 28526 0 _0077_
rlabel metal1 23138 29002 23138 29002 0 _0078_
rlabel metal1 24656 24378 24656 24378 0 _0079_
rlabel metal1 21903 24174 21903 24174 0 _0080_
rlabel metal2 18814 26792 18814 26792 0 _0081_
rlabel metal1 19412 26282 19412 26282 0 _0082_
rlabel metal1 19826 24922 19826 24922 0 _0083_
rlabel metal1 16376 19482 16376 19482 0 _0084_
rlabel metal2 21482 13090 21482 13090 0 _0085_
rlabel metal1 16836 7514 16836 7514 0 _0086_
rlabel metal1 16245 10030 16245 10030 0 _0087_
rlabel metal2 16422 11288 16422 11288 0 _0088_
rlabel metal2 15962 9384 15962 9384 0 _0089_
rlabel metal1 18400 6970 18400 6970 0 _0090_
rlabel metal1 21535 6698 21535 6698 0 _0091_
rlabel metal2 21206 7582 21206 7582 0 _0092_
rlabel metal2 22678 8738 22678 8738 0 _0093_
rlabel metal1 20891 11798 20891 11798 0 _0094_
rlabel metal1 24472 17850 24472 17850 0 _0095_
rlabel metal2 23966 11560 23966 11560 0 _0096_
rlabel metal1 23598 8602 23598 8602 0 _0097_
rlabel metal2 23690 10472 23690 10472 0 _0098_
rlabel metal2 23598 6596 23598 6596 0 _0099_
rlabel metal2 22862 7582 22862 7582 0 _0100_
rlabel metal1 26128 6426 26128 6426 0 _0101_
rlabel metal1 29309 6698 29309 6698 0 _0102_
rlabel metal1 29256 9894 29256 9894 0 _0103_
rlabel metal2 30222 8296 30222 8296 0 _0104_
rlabel metal1 28987 11050 28987 11050 0 _0105_
rlabel metal1 23559 12886 23559 12886 0 _0106_
rlabel metal2 28382 11832 28382 11832 0 _0107_
rlabel metal1 31188 9146 31188 9146 0 _0108_
rlabel metal2 30498 10472 30498 10472 0 _0109_
rlabel metal2 32062 8738 32062 8738 0 _0110_
rlabel metal1 35703 9622 35703 9622 0 _0111_
rlabel metal2 36846 10914 36846 10914 0 _0112_
rlabel metal2 33166 13464 33166 13464 0 _0113_
rlabel metal2 34362 14110 34362 14110 0 _0114_
rlabel metal2 36386 12648 36386 12648 0 _0115_
rlabel metal1 31287 13974 31287 13974 0 _0116_
rlabel metal1 35558 19244 35558 19244 0 _0117_
rlabel metal1 32609 19754 32609 19754 0 _0118_
rlabel metal1 33227 18632 33227 18632 0 _0119_
rlabel metal2 34730 17408 34730 17408 0 _0120_
rlabel metal1 37301 16558 37301 16558 0 _0121_
rlabel metal1 37290 18326 37290 18326 0 _0122_
rlabel metal1 34638 22134 34638 22134 0 _0123_
rlabel metal1 36105 24854 36105 24854 0 _0124_
rlabel metal1 34776 24378 34776 24378 0 _0125_
rlabel via1 37301 23086 37301 23086 0 _0126_
rlabel metal2 36938 21658 36938 21658 0 _0127_
rlabel metal1 31540 17578 31540 17578 0 _0128_
rlabel metal1 28193 19822 28193 19822 0 _0129_
rlabel metal1 28423 18326 28423 18326 0 _0130_
rlabel metal1 31050 17850 31050 17850 0 _0131_
rlabel metal1 31878 18938 31878 18938 0 _0132_
rlabel metal1 25146 14314 25146 14314 0 _0133_
rlabel metal1 25346 14042 25346 14042 0 _0134_
rlabel metal1 32292 20366 32292 20366 0 _0135_
rlabel via1 26721 20910 26721 20910 0 _0136_
rlabel metal1 30861 22610 30861 22610 0 _0137_
rlabel via1 32149 21930 32149 21930 0 _0138_
rlabel metal1 33994 23494 33994 23494 0 _0139_
rlabel metal1 33212 24922 33212 24922 0 _0140_
rlabel metal2 32430 26690 32430 26690 0 _0141_
rlabel metal1 30263 27030 30263 27030 0 _0142_
rlabel metal1 28708 23766 28708 23766 0 _0143_
rlabel metal1 26537 23086 26537 23086 0 _0144_
rlabel metal1 26537 25262 26537 25262 0 _0145_
rlabel metal1 26680 27098 26680 27098 0 _0146_
rlabel metal2 28658 27234 28658 27234 0 _0147_
rlabel metal2 25346 12002 25346 12002 0 _0148_
rlabel via1 32057 15470 32057 15470 0 _0149_
rlabel metal1 29992 11662 29992 11662 0 _0150_
rlabel metal1 10665 11322 10665 11322 0 _0151_
rlabel metal2 12926 14144 12926 14144 0 _0152_
rlabel metal1 12328 12274 12328 12274 0 _0153_
rlabel metal1 8832 12886 8832 12886 0 _0154_
rlabel metal1 8411 13702 8411 13702 0 _0155_
rlabel metal1 7636 15130 7636 15130 0 _0156_
rlabel metal1 9200 16762 9200 16762 0 _0157_
rlabel metal1 8740 17850 8740 17850 0 _0158_
rlabel metal1 15134 16762 15134 16762 0 _0159_
rlabel metal1 14720 14790 14720 14790 0 _0160_
rlabel metal1 8372 20502 8372 20502 0 _0161_
rlabel metal1 11040 19754 11040 19754 0 _0162_
rlabel metal1 10718 20808 10718 20808 0 _0163_
rlabel metal1 9016 22542 9016 22542 0 _0164_
rlabel metal1 9660 23630 9660 23630 0 _0165_
rlabel metal1 10304 24378 10304 24378 0 _0166_
rlabel metal2 12006 25024 12006 25024 0 _0167_
rlabel metal2 12466 26010 12466 26010 0 _0168_
rlabel metal1 14398 24378 14398 24378 0 _0169_
rlabel metal1 17388 22542 17388 22542 0 _0170_
rlabel metal1 15134 13770 15134 13770 0 _0171_
rlabel metal1 13478 18360 13478 18360 0 _0172_
rlabel metal1 20424 28186 20424 28186 0 _0173_
rlabel metal2 24702 27778 24702 27778 0 _0174_
rlabel metal2 25070 27812 25070 27812 0 _0175_
rlabel metal1 22356 28186 22356 28186 0 _0176_
rlabel metal1 23782 24854 23782 24854 0 _0177_
rlabel metal1 21114 24242 21114 24242 0 _0178_
rlabel metal2 19826 26724 19826 26724 0 _0179_
rlabel metal1 18446 25976 18446 25976 0 _0180_
rlabel metal1 20332 23290 20332 23290 0 _0181_
rlabel metal1 24104 22746 24104 22746 0 _0182_
rlabel metal1 15502 19890 15502 19890 0 _0183_
rlabel metal1 14996 22542 14996 22542 0 _0184_
rlabel metal1 14356 22678 14356 22678 0 _0185_
rlabel metal1 16008 7514 16008 7514 0 _0186_
rlabel metal1 18262 10132 18262 10132 0 _0187_
rlabel metal2 18078 11016 18078 11016 0 _0188_
rlabel metal1 15824 9486 15824 9486 0 _0189_
rlabel metal1 17618 7480 17618 7480 0 _0190_
rlabel metal1 19816 6970 19816 6970 0 _0191_
rlabel metal2 20194 7854 20194 7854 0 _0192_
rlabel metal1 20923 9146 20923 9146 0 _0193_
rlabel metal1 18344 12818 18344 12818 0 _0194_
rlabel metal1 19228 14586 19228 14586 0 _0195_
rlabel metal1 23322 18360 23322 18360 0 _0196_
rlabel metal2 26450 22338 26450 22338 0 _0197_
rlabel metal1 25249 23018 25249 23018 0 _0198_
rlabel metal1 22908 9010 22908 9010 0 _0199_
rlabel metal2 24518 10404 24518 10404 0 _0200_
rlabel metal1 23453 6970 23453 6970 0 _0201_
rlabel metal1 22954 7310 22954 7310 0 _0202_
rlabel metal2 28290 6494 28290 6494 0 _0203_
rlabel metal1 28060 6426 28060 6426 0 _0204_
rlabel metal1 28520 8942 28520 8942 0 _0205_
rlabel metal1 29026 8398 29026 8398 0 _0206_
rlabel metal1 27646 14450 27646 14450 0 _0207_
rlabel metal1 22218 12410 22218 12410 0 _0208_
rlabel metal1 17061 13294 17061 13294 0 _0209_
rlabel metal1 16560 12682 16560 12682 0 _0210_
rlabel metal2 30774 9044 30774 9044 0 _0211_
rlabel metal1 30406 10574 30406 10574 0 _0212_
rlabel metal2 32246 9180 32246 9180 0 _0213_
rlabel metal2 34270 9469 34270 9469 0 _0214_
rlabel metal1 35374 11050 35374 11050 0 _0215_
rlabel metal1 32660 12954 32660 12954 0 _0216_
rlabel metal1 35420 13294 35420 13294 0 _0217_
rlabel metal1 35788 12886 35788 12886 0 _0218_
rlabel metal2 28566 16354 28566 16354 0 _0219_
rlabel metal1 30778 16558 30778 16558 0 _0220_
rlabel metal1 32844 15130 32844 15130 0 _0221_
rlabel metal1 17618 12342 17618 12342 0 _0222_
rlabel metal1 28658 16014 28658 16014 0 _0223_
rlabel metal1 31234 15028 31234 15028 0 _0224_
rlabel metal2 33626 11798 33626 11798 0 _0225_
rlabel metal1 33718 11798 33718 11798 0 _0226_
rlabel metal1 32430 11764 32430 11764 0 _0227_
rlabel metal1 31050 12172 31050 12172 0 _0228_
rlabel metal1 36662 13362 36662 13362 0 _0229_
rlabel metal1 34914 10438 34914 10438 0 _0230_
rlabel via1 34654 13226 34654 13226 0 _0231_
rlabel metal1 35006 13430 35006 13430 0 _0232_
rlabel metal1 36386 13260 36386 13260 0 _0233_
rlabel metal1 34270 11186 34270 11186 0 _0234_
rlabel via1 36041 13226 36041 13226 0 _0235_
rlabel metal2 36708 12988 36708 12988 0 _0236_
rlabel metal2 35282 12002 35282 12002 0 _0237_
rlabel metal1 34362 12818 34362 12818 0 _0238_
rlabel metal1 31234 10030 31234 10030 0 _0239_
rlabel metal1 34454 12716 34454 12716 0 _0240_
rlabel metal1 33534 12818 33534 12818 0 _0241_
rlabel metal2 35190 10948 35190 10948 0 _0242_
rlabel metal1 33580 9554 33580 9554 0 _0243_
rlabel metal1 33396 9560 33396 9560 0 _0244_
rlabel metal1 32522 9656 32522 9656 0 _0245_
rlabel metal1 32430 9622 32430 9622 0 _0246_
rlabel metal1 31280 11322 31280 11322 0 _0247_
rlabel metal2 31786 11424 31786 11424 0 _0248_
rlabel metal1 30958 8534 30958 8534 0 _0249_
rlabel metal1 22862 12274 22862 12274 0 _0250_
rlabel metal1 22356 12274 22356 12274 0 _0251_
rlabel metal1 20562 9996 20562 9996 0 _0252_
rlabel metal1 18814 10132 18814 10132 0 _0253_
rlabel metal1 22724 10438 22724 10438 0 _0254_
rlabel metal1 20194 10030 20194 10030 0 _0255_
rlabel metal1 20792 10234 20792 10234 0 _0256_
rlabel metal1 19090 16184 19090 16184 0 _0257_
rlabel metal2 26358 9622 26358 9622 0 _0258_
rlabel metal2 26450 9316 26450 9316 0 _0259_
rlabel metal1 26450 9690 26450 9690 0 _0260_
rlabel metal1 25484 17034 25484 17034 0 _0261_
rlabel metal1 28014 10676 28014 10676 0 _0262_
rlabel metal2 25990 7854 25990 7854 0 _0263_
rlabel metal1 26634 7310 26634 7310 0 _0264_
rlabel metal1 28214 8874 28214 8874 0 _0265_
rlabel metal2 28290 8636 28290 8636 0 _0266_
rlabel metal1 29394 8058 29394 8058 0 _0267_
rlabel metal2 27830 10064 27830 10064 0 _0268_
rlabel metal1 29417 8874 29417 8874 0 _0269_
rlabel metal1 28428 8466 28428 8466 0 _0270_
rlabel metal1 25300 9622 25300 9622 0 _0271_
rlabel metal2 27370 7174 27370 7174 0 _0272_
rlabel metal1 28014 7446 28014 7446 0 _0273_
rlabel metal1 27554 7310 27554 7310 0 _0274_
rlabel metal1 28382 6290 28382 6290 0 _0275_
rlabel metal1 25438 7752 25438 7752 0 _0276_
rlabel metal1 25254 7854 25254 7854 0 _0277_
rlabel metal1 24472 7446 24472 7446 0 _0278_
rlabel metal1 24702 7378 24702 7378 0 _0279_
rlabel metal1 25576 10642 25576 10642 0 _0280_
rlabel metal1 23552 9554 23552 9554 0 _0281_
rlabel metal1 23690 18700 23690 18700 0 _0282_
rlabel metal1 23690 18802 23690 18802 0 _0283_
rlabel metal1 22494 26928 22494 26928 0 _0284_
rlabel metal2 22218 24990 22218 24990 0 _0285_
rlabel metal1 22448 23630 22448 23630 0 _0286_
rlabel metal1 23322 26554 23322 26554 0 _0287_
rlabel metal1 23598 25874 23598 25874 0 _0288_
rlabel metal1 20332 22610 20332 22610 0 _0289_
rlabel metal1 20332 11118 20332 11118 0 _0290_
rlabel metal1 18568 9622 18568 9622 0 _0291_
rlabel metal1 18906 8874 18906 8874 0 _0292_
rlabel metal1 19672 8874 19672 8874 0 _0293_
rlabel metal1 20838 8806 20838 8806 0 _0294_
rlabel metal1 20286 9078 20286 9078 0 _0295_
rlabel metal1 20332 9622 20332 9622 0 _0296_
rlabel metal2 20746 8942 20746 8942 0 _0297_
rlabel metal1 21068 8602 21068 8602 0 _0298_
rlabel metal1 19542 8602 19542 8602 0 _0299_
rlabel metal2 19642 8092 19642 8092 0 _0300_
rlabel metal2 18446 11390 18446 11390 0 _0301_
rlabel metal2 19090 8092 19090 8092 0 _0302_
rlabel metal1 19320 7378 19320 7378 0 _0303_
rlabel metal1 18078 7820 18078 7820 0 _0304_
rlabel metal1 17388 9146 17388 9146 0 _0305_
rlabel metal1 16882 9520 16882 9520 0 _0306_
rlabel metal2 18354 11390 18354 11390 0 _0307_
rlabel viali 18262 10664 18262 10664 0 _0308_
rlabel metal1 18814 9962 18814 9962 0 _0309_
rlabel metal1 16468 7378 16468 7378 0 _0310_
rlabel metal1 15686 20468 15686 20468 0 _0311_
rlabel metal1 15686 20230 15686 20230 0 _0312_
rlabel metal1 12604 22134 12604 22134 0 _0313_
rlabel metal1 13662 22542 13662 22542 0 _0314_
rlabel metal1 12581 22542 12581 22542 0 _0315_
rlabel metal1 12604 21998 12604 21998 0 _0316_
rlabel metal1 12604 22610 12604 22610 0 _0317_
rlabel metal1 13156 22746 13156 22746 0 _0318_
rlabel metal1 15410 20502 15410 20502 0 _0319_
rlabel metal1 21988 26010 21988 26010 0 _0320_
rlabel metal1 22034 25364 22034 25364 0 _0321_
rlabel metal1 22586 27098 22586 27098 0 _0322_
rlabel metal1 21436 26758 21436 26758 0 _0323_
rlabel metal1 21377 27098 21377 27098 0 _0324_
rlabel metal1 21344 26486 21344 26486 0 _0325_
rlabel metal2 22586 27676 22586 27676 0 _0326_
rlabel metal1 22704 28084 22704 28084 0 _0327_
rlabel metal2 20286 26554 20286 26554 0 _0328_
rlabel metal1 19734 26452 19734 26452 0 _0329_
rlabel metal1 20010 26452 20010 26452 0 _0330_
rlabel metal2 22356 24786 22356 24786 0 _0331_
rlabel metal2 23690 24939 23690 24939 0 _0332_
rlabel metal1 23230 25160 23230 25160 0 _0333_
rlabel metal1 22494 24854 22494 24854 0 _0334_
rlabel metal1 22678 27642 22678 27642 0 _0335_
rlabel metal1 25668 27302 25668 27302 0 _0336_
rlabel metal1 25162 26928 25162 26928 0 _0337_
rlabel metal2 24794 27234 24794 27234 0 _0338_
rlabel metal1 24886 27472 24886 27472 0 _0339_
rlabel metal1 24840 27030 24840 27030 0 _0340_
rlabel metal1 20700 28050 20700 28050 0 _0341_
rlabel metal1 13708 18802 13708 18802 0 _0342_
rlabel metal1 13340 18802 13340 18802 0 _0343_
rlabel metal1 12466 14450 12466 14450 0 _0344_
rlabel metal1 11454 15470 11454 15470 0 _0345_
rlabel metal1 11454 14994 11454 14994 0 _0346_
rlabel metal1 11454 15062 11454 15062 0 _0347_
rlabel metal1 12052 14994 12052 14994 0 _0348_
rlabel metal2 13386 18530 13386 18530 0 _0349_
rlabel metal1 13432 24786 13432 24786 0 _0350_
rlabel metal1 11500 23698 11500 23698 0 _0351_
rlabel metal2 13386 24514 13386 24514 0 _0352_
rlabel metal1 13570 25398 13570 25398 0 _0353_
rlabel metal1 13202 25466 13202 25466 0 _0354_
rlabel metal2 12926 23970 12926 23970 0 _0355_
rlabel metal1 12558 24072 12558 24072 0 _0356_
rlabel metal1 12696 24174 12696 24174 0 _0357_
rlabel metal1 12466 24820 12466 24820 0 _0358_
rlabel metal1 12190 25874 12190 25874 0 _0359_
rlabel metal1 12052 24786 12052 24786 0 _0360_
rlabel metal1 10672 23766 10672 23766 0 _0361_
rlabel metal2 10534 24004 10534 24004 0 _0362_
rlabel metal1 11270 24106 11270 24106 0 _0363_
rlabel metal1 11546 23290 11546 23290 0 _0364_
rlabel metal1 11132 23290 11132 23290 0 _0365_
rlabel metal1 10074 22576 10074 22576 0 _0366_
rlabel metal1 10120 22202 10120 22202 0 _0367_
rlabel metal1 11408 20570 11408 20570 0 _0368_
rlabel metal1 11730 20910 11730 20910 0 _0369_
rlabel metal2 11730 21046 11730 21046 0 _0370_
rlabel metal1 8970 21522 8970 21522 0 _0371_
rlabel metal1 11730 13430 11730 13430 0 _0372_
rlabel viali 10074 13905 10074 13905 0 _0373_
rlabel metal1 9782 16150 9782 16150 0 _0374_
rlabel metal2 9706 16694 9706 16694 0 _0375_
rlabel metal1 11454 16524 11454 16524 0 _0376_
rlabel metal1 11316 16422 11316 16422 0 _0377_
rlabel metal1 10166 16490 10166 16490 0 _0378_
rlabel metal2 9982 16864 9982 16864 0 _0379_
rlabel metal1 9292 17034 9292 17034 0 _0380_
rlabel metal2 10166 14756 10166 14756 0 _0381_
rlabel metal1 9752 15402 9752 15402 0 _0382_
rlabel metal1 12098 12818 12098 12818 0 _0383_
rlabel metal1 9476 14382 9476 14382 0 _0384_
rlabel metal1 8142 15028 8142 15028 0 _0385_
rlabel metal1 11684 14042 11684 14042 0 _0386_
rlabel metal1 10534 13804 10534 13804 0 _0387_
rlabel metal1 9706 13328 9706 13328 0 _0388_
rlabel metal1 11960 12886 11960 12886 0 _0389_
rlabel metal2 12558 14722 12558 14722 0 _0390_
rlabel metal1 12558 14416 12558 14416 0 _0391_
rlabel metal1 11224 12206 11224 12206 0 _0392_
rlabel metal1 30406 12886 30406 12886 0 _0393_
rlabel metal1 29716 12410 29716 12410 0 _0394_
rlabel metal1 30774 13498 30774 13498 0 _0395_
rlabel metal2 25530 11798 25530 11798 0 _0396_
rlabel metal2 25714 11900 25714 11900 0 _0397_
rlabel metal2 15594 18462 15594 18462 0 _0398_
rlabel metal1 35466 18292 35466 18292 0 _0399_
rlabel metal1 18170 21930 18170 21930 0 _0400_
rlabel metal2 21850 17952 21850 17952 0 _0401_
rlabel metal2 33902 20978 33902 20978 0 _0402_
rlabel metal1 26772 15674 26772 15674 0 _0403_
rlabel metal1 27554 17306 27554 17306 0 _0404_
rlabel metal1 18308 20434 18308 20434 0 _0405_
rlabel metal1 18170 20570 18170 20570 0 _0406_
rlabel metal1 13938 19278 13938 19278 0 _0407_
rlabel metal2 31970 13333 31970 13333 0 _0408_
rlabel metal1 16974 14348 16974 14348 0 _0409_
rlabel metal2 22218 16456 22218 16456 0 _0410_
rlabel metal1 20470 18190 20470 18190 0 _0411_
rlabel metal1 35328 14382 35328 14382 0 _0412_
rlabel metal1 28704 15062 28704 15062 0 _0413_
rlabel metal2 27830 15130 27830 15130 0 _0414_
rlabel metal1 19826 20434 19826 20434 0 _0415_
rlabel metal1 20654 18666 20654 18666 0 _0416_
rlabel metal1 22954 17578 22954 17578 0 _0417_
rlabel metal1 34730 15334 34730 15334 0 _0418_
rlabel metal1 34178 15538 34178 15538 0 _0419_
rlabel metal1 24334 14960 24334 14960 0 _0420_
rlabel metal1 14674 24140 14674 24140 0 _0421_
rlabel metal1 18998 17068 18998 17068 0 _0422_
rlabel metal2 21206 19856 21206 19856 0 _0423_
rlabel metal1 20976 19346 20976 19346 0 _0424_
rlabel metal1 35650 14892 35650 14892 0 _0425_
rlabel metal1 31050 15504 31050 15504 0 _0426_
rlabel metal1 31234 14382 31234 14382 0 _0427_
rlabel metal1 28428 26010 28428 26010 0 _0428_
rlabel metal1 28658 25296 28658 25296 0 _0429_
rlabel metal1 31326 24684 31326 24684 0 _0430_
rlabel metal1 30774 24786 30774 24786 0 _0431_
rlabel metal1 29335 24922 29335 24922 0 _0432_
rlabel metal1 29302 24650 29302 24650 0 _0433_
rlabel metal1 27738 22066 27738 22066 0 _0434_
rlabel metal1 28704 20774 28704 20774 0 _0435_
rlabel metal1 29946 20400 29946 20400 0 _0436_
rlabel metal1 30406 19754 30406 19754 0 _0437_
rlabel metal1 29624 20570 29624 20570 0 _0438_
rlabel metal2 21022 20400 21022 20400 0 _0439_
rlabel via1 36010 21930 36010 21930 0 _0440_
rlabel viali 35742 20433 35742 20433 0 _0441_
rlabel metal2 35374 18054 35374 18054 0 _0442_
rlabel metal1 35328 20026 35328 20026 0 _0443_
rlabel metal1 35282 20570 35282 20570 0 _0444_
rlabel metal1 33994 20876 33994 20876 0 _0445_
rlabel metal1 34316 20910 34316 20910 0 _0446_
rlabel metal1 32936 19346 32936 19346 0 _0447_
rlabel metal2 34822 18938 34822 18938 0 _0448_
rlabel via1 36731 20434 36731 20434 0 _0449_
rlabel metal1 36478 20400 36478 20400 0 _0450_
rlabel metal1 26358 18122 26358 18122 0 _0451_
rlabel metal1 16464 17306 16464 17306 0 _0452_
rlabel metal1 16974 16082 16974 16082 0 _0453_
rlabel metal1 17296 14450 17296 14450 0 _0454_
rlabel metal1 20562 14960 20562 14960 0 _0455_
rlabel viali 19182 14993 19182 14993 0 _0456_
rlabel metal1 17526 24276 17526 24276 0 _0457_
rlabel metal1 19136 15946 19136 15946 0 _0458_
rlabel metal1 23046 15402 23046 15402 0 _0459_
rlabel metal1 18124 23290 18124 23290 0 _0460_
rlabel metal1 18308 23698 18308 23698 0 _0461_
rlabel metal1 24288 20910 24288 20910 0 _0462_
rlabel metal2 23506 20876 23506 20876 0 _0463_
rlabel metal1 25576 21998 25576 21998 0 _0464_
rlabel metal2 26082 13192 26082 13192 0 _0465_
rlabel metal1 21482 14042 21482 14042 0 _0466_
rlabel metal2 20746 18088 20746 18088 0 _0467_
rlabel metal2 19458 17816 19458 17816 0 _0468_
rlabel metal2 20286 14620 20286 14620 0 _0469_
rlabel metal1 23736 12954 23736 12954 0 _0470_
rlabel metal1 22678 13498 22678 13498 0 _0471_
rlabel metal1 16376 18734 16376 18734 0 _0472_
rlabel metal1 14628 18938 14628 18938 0 _0473_
rlabel metal1 13064 19482 13064 19482 0 _0474_
rlabel metal1 13156 22134 13156 22134 0 _0475_
rlabel metal1 13064 20502 13064 20502 0 _0476_
rlabel metal1 13340 21862 13340 21862 0 _0477_
rlabel metal1 12512 20434 12512 20434 0 _0478_
rlabel metal1 13018 20332 13018 20332 0 _0479_
rlabel metal2 24978 26044 24978 26044 0 _0480_
rlabel metal1 25438 25738 25438 25738 0 _0481_
rlabel via1 25343 25262 25343 25262 0 _0482_
rlabel metal1 25622 24922 25622 24922 0 _0483_
rlabel metal1 24978 25466 24978 25466 0 _0484_
rlabel metal1 23598 19958 23598 19958 0 _0485_
rlabel metal2 23046 21053 23046 21053 0 _0486_
rlabel metal2 25070 8976 25070 8976 0 _0487_
rlabel metal1 26082 10642 26082 10642 0 _0488_
rlabel metal1 26036 13906 26036 13906 0 _0489_
rlabel metal1 25576 10166 25576 10166 0 _0490_
rlabel metal1 25576 9146 25576 9146 0 _0491_
rlabel metal1 24840 9146 24840 9146 0 _0492_
rlabel metal1 25622 9690 25622 9690 0 _0493_
rlabel metal2 25254 10880 25254 10880 0 _0494_
rlabel metal1 34040 15334 34040 15334 0 _0495_
rlabel metal2 32706 13090 32706 13090 0 _0496_
rlabel metal1 32430 11220 32430 11220 0 _0497_
rlabel viali 32982 11729 32982 11729 0 _0498_
rlabel metal2 32614 11628 32614 11628 0 _0499_
rlabel metal1 32982 11118 32982 11118 0 _0500_
rlabel metal1 32613 11118 32613 11118 0 _0501_
rlabel metal1 31786 11118 31786 11118 0 _0502_
rlabel viali 18613 11118 18613 11118 0 _0503_
rlabel metal1 18413 11050 18413 11050 0 _0504_
rlabel metal1 18676 9554 18676 9554 0 _0505_
rlabel metal2 18170 10370 18170 10370 0 _0506_
rlabel metal2 18722 11424 18722 11424 0 _0507_
rlabel metal2 22310 11220 22310 11220 0 _0508_
rlabel metal2 22402 15300 22402 15300 0 _0509_
rlabel via2 13938 20451 13938 20451 0 _0510_
rlabel metal2 13294 18156 13294 18156 0 _0511_
rlabel metal1 12834 14858 12834 14858 0 _0512_
rlabel metal1 12696 14790 12696 14790 0 _0513_
rlabel metal1 12098 15674 12098 15674 0 _0514_
rlabel metal1 12144 16218 12144 16218 0 _0515_
rlabel metal1 13018 15130 13018 15130 0 _0516_
rlabel metal1 10580 17850 10580 17850 0 _0517_
rlabel metal1 14628 25262 14628 25262 0 _0518_
rlabel metal1 19458 24378 19458 24378 0 _0519_
rlabel metal1 19964 11118 19964 11118 0 _0520_
rlabel metal1 26634 11696 26634 11696 0 _0521_
rlabel metal2 30406 13940 30406 13940 0 _0522_
rlabel metal1 17388 16218 17388 16218 0 _0523_
rlabel metal1 18170 16592 18170 16592 0 _0524_
rlabel metal1 25668 17306 25668 17306 0 _0525_
rlabel metal1 18032 23494 18032 23494 0 _0526_
rlabel metal1 18676 23086 18676 23086 0 _0527_
rlabel metal1 16652 23834 16652 23834 0 _0528_
rlabel metal1 18538 15028 18538 15028 0 _0529_
rlabel metal1 21298 14994 21298 14994 0 _0530_
rlabel metal1 29440 21522 29440 21522 0 _0531_
rlabel metal1 29210 20876 29210 20876 0 _0532_
rlabel metal1 24104 20434 24104 20434 0 _0533_
rlabel metal1 24334 19822 24334 19822 0 _0534_
rlabel metal1 37214 19958 37214 19958 0 _0535_
rlabel metal1 32660 19210 32660 19210 0 _0536_
rlabel metal1 33902 19244 33902 19244 0 _0537_
rlabel metal1 34868 17170 34868 17170 0 _0538_
rlabel metal1 36662 17034 36662 17034 0 _0539_
rlabel metal1 37490 18700 37490 18700 0 _0540_
rlabel metal1 37122 18122 37122 18122 0 _0541_
rlabel metal1 35274 21998 35274 21998 0 _0542_
rlabel metal1 34684 21998 34684 21998 0 _0543_
rlabel metal1 34914 21964 34914 21964 0 _0544_
rlabel metal1 35512 24174 35512 24174 0 _0545_
rlabel metal2 37306 24820 37306 24820 0 _0546_
rlabel metal1 35512 23834 35512 23834 0 _0547_
rlabel metal1 36386 23290 36386 23290 0 _0548_
rlabel metal2 36616 21828 36616 21828 0 _0549_
rlabel metal1 36938 21624 36938 21624 0 _0550_
rlabel metal1 31418 17748 31418 17748 0 _0551_
rlabel metal2 29302 20298 29302 20298 0 _0552_
rlabel metal1 28888 20298 28888 20298 0 _0553_
rlabel metal1 29026 18700 29026 18700 0 _0554_
rlabel metal1 28566 18666 28566 18666 0 _0555_
rlabel metal1 30360 17034 30360 17034 0 _0556_
rlabel metal1 31142 18870 31142 18870 0 _0557_
rlabel metal1 26312 14042 26312 14042 0 _0558_
rlabel metal1 31280 20298 31280 20298 0 _0559_
rlabel metal1 31004 24786 31004 24786 0 _0560_
rlabel metal1 30866 24922 30866 24922 0 _0561_
rlabel metal1 33271 22950 33271 22950 0 _0562_
rlabel metal1 32476 22406 32476 22406 0 _0563_
rlabel metal1 31464 22066 31464 22066 0 _0564_
rlabel metal1 32844 23290 32844 23290 0 _0565_
rlabel metal1 32338 22678 32338 22678 0 _0566_
rlabel metal1 33902 23800 33902 23800 0 _0567_
rlabel metal1 31740 24922 31740 24922 0 _0568_
rlabel metal1 31326 25296 31326 25296 0 _0569_
rlabel metal1 32016 25466 32016 25466 0 _0570_
rlabel metal1 32292 24378 32292 24378 0 _0571_
rlabel metal1 32890 24820 32890 24820 0 _0572_
rlabel metal1 32338 26418 32338 26418 0 _0573_
rlabel metal1 32522 26384 32522 26384 0 _0574_
rlabel metal1 30682 26384 30682 26384 0 _0575_
rlabel metal1 30590 26418 30590 26418 0 _0576_
rlabel metal1 30314 25874 30314 25874 0 _0577_
rlabel metal1 30452 25806 30452 25806 0 _0578_
rlabel metal1 27784 24242 27784 24242 0 _0579_
rlabel metal1 27968 23290 27968 23290 0 _0580_
rlabel metal1 28290 23290 28290 23290 0 _0581_
rlabel metal1 26864 23698 26864 23698 0 _0582_
rlabel via1 27462 26894 27462 26894 0 _0583_
rlabel metal1 27600 25466 27600 25466 0 _0584_
rlabel metal1 26910 25874 26910 25874 0 _0585_
rlabel metal1 29118 26928 29118 26928 0 _0586_
rlabel metal1 26634 26996 26634 26996 0 _0587_
rlabel metal1 29210 26554 29210 26554 0 _0588_
rlabel metal1 9476 12206 9476 12206 0 _0589_
rlabel metal2 32522 15776 32522 15776 0 _0590_
rlabel metal1 14674 20332 14674 20332 0 _0591_
rlabel metal2 15962 15844 15962 15844 0 _0592_
rlabel metal1 14858 15028 14858 15028 0 _0593_
rlabel metal1 15916 19482 15916 19482 0 _0594_
rlabel metal1 16146 23494 16146 23494 0 _0595_
rlabel metal1 17894 22576 17894 22576 0 _0596_
rlabel metal1 17986 13294 17986 13294 0 _0597_
rlabel metal1 15686 14892 15686 14892 0 _0598_
rlabel metal1 21022 18326 21022 18326 0 _0599_
rlabel metal1 22954 22134 22954 22134 0 _0600_
rlabel metal1 23598 22644 23598 22644 0 _0601_
rlabel metal1 16836 22610 16836 22610 0 _0602_
rlabel metal2 14398 23290 14398 23290 0 _0603_
rlabel metal2 21850 7310 21850 7310 0 _0604_
rlabel metal1 18216 13906 18216 13906 0 _0605_
rlabel metal1 20562 13838 20562 13838 0 _0606_
rlabel metal1 24702 22066 24702 22066 0 _0607_
rlabel metal1 25392 23834 25392 23834 0 _0608_
rlabel metal1 24380 12818 24380 12818 0 _0609_
rlabel metal1 17943 14042 17943 14042 0 _0610_
rlabel metal2 4094 17867 4094 17867 0 clk
rlabel metal1 14766 12818 14766 12818 0 clknet_0_clk
rlabel metal1 15732 7922 15732 7922 0 clknet_4_0_0_clk
rlabel metal1 35236 13906 35236 13906 0 clknet_4_10_0_clk
rlabel metal1 32982 16082 32982 16082 0 clknet_4_11_0_clk
rlabel metal1 22908 20910 22908 20910 0 clknet_4_12_0_clk
rlabel metal1 25714 28084 25714 28084 0 clknet_4_13_0_clk
rlabel metal2 37306 19312 37306 19312 0 clknet_4_14_0_clk
rlabel metal1 33672 21590 33672 21590 0 clknet_4_15_0_clk
rlabel metal1 11960 12274 11960 12274 0 clknet_4_1_0_clk
rlabel metal1 21712 12750 21712 12750 0 clknet_4_2_0_clk
rlabel metal2 17618 16320 17618 16320 0 clknet_4_3_0_clk
rlabel metal2 12558 20366 12558 20366 0 clknet_4_4_0_clk
rlabel metal1 13386 21454 13386 21454 0 clknet_4_5_0_clk
rlabel metal1 17664 18734 17664 18734 0 clknet_4_6_0_clk
rlabel metal1 18078 22066 18078 22066 0 clknet_4_7_0_clk
rlabel metal2 29118 12585 29118 12585 0 clknet_4_8_0_clk
rlabel metal1 24794 15470 24794 15470 0 clknet_4_9_0_clk
rlabel metal1 15870 15062 15870 15062 0 conv1.addr\[8\]
rlabel metal1 13156 16082 13156 16082 0 conv1.data_valid
rlabel metal2 18998 17748 18998 17748 0 conv1.done
rlabel metal1 13018 18734 13018 18734 0 conv1.psram_ce_n
rlabel metal2 12190 11934 12190 11934 0 conv1.psram_ctrl.counter\[0\]
rlabel metal1 12926 13328 12926 13328 0 conv1.psram_ctrl.counter\[1\]
rlabel metal1 13754 12750 13754 12750 0 conv1.psram_ctrl.counter\[2\]
rlabel metal2 10718 13022 10718 13022 0 conv1.psram_ctrl.counter\[3\]
rlabel metal1 10994 13974 10994 13974 0 conv1.psram_ctrl.counter\[4\]
rlabel metal1 9200 15538 9200 15538 0 conv1.psram_ctrl.counter\[5\]
rlabel metal1 10902 16014 10902 16014 0 conv1.psram_ctrl.counter\[6\]
rlabel metal1 9706 18054 9706 18054 0 conv1.psram_ctrl.counter\[7\]
rlabel metal1 14306 15028 14306 15028 0 conv1.psram_ctrl.has_wait_states
rlabel metal1 10028 18326 10028 18326 0 conv1.psram_ctrl.nstate
rlabel metal1 16146 18326 16146 18326 0 conv1.psram_ctrl.sck
rlabel metal1 13018 17068 13018 17068 0 conv1.psram_ctrl.start
rlabel metal1 11454 18394 11454 18394 0 conv1.psram_ctrl.state
rlabel metal1 18676 18802 18676 18802 0 conv1.state\[0\]
rlabel metal1 16054 17510 16054 17510 0 conv1.state\[1\]
rlabel metal1 14720 16014 14720 16014 0 conv1.state\[2\]
rlabel via1 16054 17102 16054 17102 0 conv1.state\[3\]
rlabel metal1 16928 17170 16928 17170 0 conv1.state\[5\]
rlabel metal1 14444 21998 14444 21998 0 conv2.addr\[8\]
rlabel metal1 13432 21998 13432 21998 0 conv2.addr\[9\]
rlabel metal1 18400 21658 18400 21658 0 conv2.data_out_valid
rlabel metal1 14030 20400 14030 20400 0 conv2.data_valid
rlabel metal1 15962 20400 15962 20400 0 conv2.psram_ce_n
rlabel metal1 13156 20434 13156 20434 0 conv2.psram_ctrl.counter\[0\]
rlabel metal1 12466 21522 12466 21522 0 conv2.psram_ctrl.counter\[1\]
rlabel metal1 12788 23154 12788 23154 0 conv2.psram_ctrl.counter\[2\]
rlabel metal1 12144 22610 12144 22610 0 conv2.psram_ctrl.counter\[3\]
rlabel metal1 9844 23834 9844 23834 0 conv2.psram_ctrl.counter\[4\]
rlabel metal1 12926 21964 12926 21964 0 conv2.psram_ctrl.counter\[5\]
rlabel metal1 13294 25296 13294 25296 0 conv2.psram_ctrl.counter\[6\]
rlabel metal1 13478 25806 13478 25806 0 conv2.psram_ctrl.counter\[7\]
rlabel metal1 15594 22610 15594 22610 0 conv2.psram_ctrl.has_wait_states
rlabel metal1 14352 25466 14352 25466 0 conv2.psram_ctrl.nstate
rlabel metal2 16054 20910 16054 20910 0 conv2.psram_ctrl.sck
rlabel metal1 15732 24922 15732 24922 0 conv2.psram_ctrl.start
rlabel metal1 15548 25330 15548 25330 0 conv2.psram_ctrl.state
rlabel metal1 17848 21114 17848 21114 0 conv2.state\[0\]
rlabel metal2 16698 23358 16698 23358 0 conv2.state\[1\]
rlabel metal1 16790 23630 16790 23630 0 conv2.state\[2\]
rlabel metal1 17572 20502 17572 20502 0 conv2.state\[3\]
rlabel metal1 18400 24786 18400 24786 0 conv2.state\[5\]
rlabel metal1 67988 2278 67988 2278 0 done
rlabel metal1 26036 23698 26036 23698 0 fc1.addr\[10\]
rlabel metal1 24748 22746 24748 22746 0 fc1.addr\[8\]
rlabel metal1 23782 17714 23782 17714 0 fc1.data_out_valid
rlabel metal2 22126 20332 22126 20332 0 fc1.psram_ce_n
rlabel metal2 22126 28220 22126 28220 0 fc1.psram_ctrl.counter\[0\]
rlabel metal1 25944 26962 25944 26962 0 fc1.psram_ctrl.counter\[1\]
rlabel metal2 25438 26928 25438 26928 0 fc1.psram_ctrl.counter\[2\]
rlabel metal2 22678 23902 22678 23902 0 fc1.psram_ctrl.counter\[3\]
rlabel metal1 22310 25262 22310 25262 0 fc1.psram_ctrl.counter\[4\]
rlabel metal1 22172 24786 22172 24786 0 fc1.psram_ctrl.counter\[5\]
rlabel metal1 21022 26894 21022 26894 0 fc1.psram_ctrl.counter\[6\]
rlabel via1 20378 25942 20378 25942 0 fc1.psram_ctrl.counter\[7\]
rlabel metal1 23092 23698 23092 23698 0 fc1.psram_ctrl.has_wait_states
rlabel metal2 19458 25058 19458 25058 0 fc1.psram_ctrl.nstate
rlabel metal1 24610 18802 24610 18802 0 fc1.psram_ctrl.sck
rlabel metal1 20792 23834 20792 23834 0 fc1.psram_ctrl.start
rlabel metal1 20930 25126 20930 25126 0 fc1.psram_ctrl.state
rlabel metal1 20884 20434 20884 20434 0 fc1.state\[0\]
rlabel metal1 25116 20774 25116 20774 0 fc1.state\[1\]
rlabel metal1 24840 21114 24840 21114 0 fc1.state\[2\]
rlabel metal1 22356 20434 22356 20434 0 fc1.state\[3\]
rlabel metal1 26312 20570 26312 20570 0 fc1.state\[5\]
rlabel metal2 16974 12988 16974 12988 0 fc2.addr\[10\]
rlabel metal1 18262 13498 18262 13498 0 fc2.addr\[8\]
rlabel metal1 23828 15470 23828 15470 0 fc2.done
rlabel metal2 21850 12682 21850 12682 0 fc2.psram_ce_n
rlabel metal1 17526 10710 17526 10710 0 fc2.psram_ctrl.counter\[0\]
rlabel metal1 19228 10574 19228 10574 0 fc2.psram_ctrl.counter\[1\]
rlabel metal1 17296 11118 17296 11118 0 fc2.psram_ctrl.counter\[2\]
rlabel metal1 19274 9622 19274 9622 0 fc2.psram_ctrl.counter\[3\]
rlabel metal1 19136 11050 19136 11050 0 fc2.psram_ctrl.counter\[4\]
rlabel metal1 19458 10064 19458 10064 0 fc2.psram_ctrl.counter\[5\]
rlabel metal2 21942 8976 21942 8976 0 fc2.psram_ctrl.counter\[6\]
rlabel metal1 22402 9486 22402 9486 0 fc2.psram_ctrl.counter\[7\]
rlabel metal1 19182 14042 19182 14042 0 fc2.psram_ctrl.has_wait_states
rlabel metal2 19734 11560 19734 11560 0 fc2.psram_ctrl.nstate
rlabel metal1 21666 12138 21666 12138 0 fc2.psram_ctrl.sck
rlabel metal1 20194 12716 20194 12716 0 fc2.psram_ctrl.start
rlabel metal1 21068 12750 21068 12750 0 fc2.psram_ctrl.state
rlabel metal1 22954 16082 22954 16082 0 fc2.state\[0\]
rlabel metal2 18998 16320 18998 16320 0 fc2.state\[1\]
rlabel metal2 17710 14620 17710 14620 0 fc2.state\[2\]
rlabel metal1 18814 14416 18814 14416 0 fc2.state\[3\]
rlabel metal1 20976 16218 20976 16218 0 fc2.state\[5\]
rlabel metal1 24702 14484 24702 14484 0 maxpool.addr\[11\]
rlabel metal2 26726 14076 26726 14076 0 maxpool.addr\[8\]
rlabel metal1 26634 15878 26634 15878 0 maxpool.done
rlabel metal1 25024 12750 25024 12750 0 maxpool.psram_ce_n
rlabel metal1 25898 9962 25898 9962 0 maxpool.psram_ctrl.counter\[0\]
rlabel metal1 25392 8466 25392 8466 0 maxpool.psram_ctrl.counter\[1\]
rlabel metal1 25714 8976 25714 8976 0 maxpool.psram_ctrl.counter\[2\]
rlabel metal1 24288 7854 24288 7854 0 maxpool.psram_ctrl.counter\[3\]
rlabel metal1 26496 7310 26496 7310 0 maxpool.psram_ctrl.counter\[4\]
rlabel metal2 28888 8874 28888 8874 0 maxpool.psram_ctrl.counter\[5\]
rlabel metal1 29578 9418 29578 9418 0 maxpool.psram_ctrl.counter\[6\]
rlabel metal2 30682 8772 30682 8772 0 maxpool.psram_ctrl.counter\[7\]
rlabel metal1 27462 11186 27462 11186 0 maxpool.psram_ctrl.nstate
rlabel metal1 25622 12852 25622 12852 0 maxpool.psram_ctrl.sck
rlabel metal1 28566 13362 28566 13362 0 maxpool.psram_ctrl.start
rlabel metal2 28106 11152 28106 11152 0 maxpool.psram_ctrl.state
rlabel metal1 25944 12750 25944 12750 0 maxpool.start
rlabel metal1 27416 16218 27416 16218 0 maxpool.state\[0\]
rlabel metal1 27094 17850 27094 17850 0 maxpool.state\[2\]
rlabel metal1 26496 14790 26496 14790 0 maxpool.state\[3\]
rlabel metal1 25944 18258 25944 18258 0 maxpool.state\[4\]
rlabel metal1 33120 20978 33120 20978 0 mfcc.dct.data_valid
rlabel metal1 32936 17714 32936 17714 0 mfcc.dct.dct_valid
rlabel metal1 35742 22542 35742 22542 0 mfcc.dct.input_counter\[0\]
rlabel metal1 37122 24684 37122 24684 0 mfcc.dct.input_counter\[1\]
rlabel metal1 36800 21862 36800 21862 0 mfcc.dct.input_counter\[2\]
rlabel metal1 38180 22610 38180 22610 0 mfcc.dct.input_counter\[3\]
rlabel metal1 38364 22066 38364 22066 0 mfcc.dct.input_counter\[4\]
rlabel metal1 36800 19822 36800 19822 0 mfcc.dct.output_counter\[0\]
rlabel metal2 34914 19414 34914 19414 0 mfcc.dct.output_counter\[1\]
rlabel metal2 34638 19108 34638 19108 0 mfcc.dct.output_counter\[2\]
rlabel metal1 36846 17680 36846 17680 0 mfcc.dct.output_counter\[3\]
rlabel metal1 37536 17578 37536 17578 0 mfcc.dct.output_counter\[4\]
rlabel via1 36478 18258 36478 18258 0 mfcc.dct.output_counter\[5\]
rlabel metal1 38640 20910 38640 20910 0 mfcc.dct.state\[0\]
rlabel metal1 35144 21590 35144 21590 0 mfcc.dct.state\[1\]
rlabel metal2 27830 21556 27830 21556 0 mfcc.log.data_valid
rlabel metal1 30130 19924 30130 19924 0 mfcc.log.shift_count\[0\]
rlabel metal1 29670 18734 29670 18734 0 mfcc.log.shift_count\[1\]
rlabel metal2 30314 18190 30314 18190 0 mfcc.log.shift_count\[2\]
rlabel metal1 30682 19142 30682 19142 0 mfcc.log.shift_count\[3\]
rlabel metal1 28750 21658 28750 21658 0 mfcc.log.state\[0\]
rlabel metal1 30590 19856 30590 19856 0 mfcc.log.state\[1\]
rlabel metal1 29164 21454 29164 21454 0 mfcc.log.state\[2\]
rlabel metal2 27738 26044 27738 26044 0 mfcc.mel.coeff_counter\[0\]
rlabel metal1 27692 23630 27692 23630 0 mfcc.mel.coeff_counter\[1\]
rlabel metal1 28014 25942 28014 25942 0 mfcc.mel.coeff_counter\[2\]
rlabel metal2 27738 27132 27738 27132 0 mfcc.mel.coeff_counter\[3\]
rlabel metal1 29854 26316 29854 26316 0 mfcc.mel.coeff_counter\[4\]
rlabel metal1 32614 23256 32614 23256 0 mfcc.mel.filter_counter\[0\]
rlabel metal1 33396 23086 33396 23086 0 mfcc.mel.filter_counter\[1\]
rlabel metal2 33074 23834 33074 23834 0 mfcc.mel.filter_counter\[2\]
rlabel metal1 31924 24854 31924 24854 0 mfcc.mel.filter_counter\[3\]
rlabel metal1 34316 26826 34316 26826 0 mfcc.mel.filter_counter\[4\]
rlabel metal1 31878 26384 31878 26384 0 mfcc.mel.filter_counter\[5\]
rlabel metal1 31004 23630 31004 23630 0 mfcc.mel.state\[0\]
rlabel metal1 28014 25262 28014 25262 0 mfcc.mel.state\[1\]
rlabel metal1 33534 17306 33534 17306 0 mfcc.mfcc_valid
rlabel metal1 10028 37298 10028 37298 0 net1
rlabel metal2 68494 55981 68494 55981 0 net10
rlabel metal1 15272 25194 15272 25194 0 net100
rlabel metal1 35374 17136 35374 17136 0 net101
rlabel metal1 38226 17238 38226 17238 0 net102
rlabel metal1 29394 8942 29394 8942 0 net103
rlabel metal2 27830 9316 27830 9316 0 net104
rlabel metal1 19964 24106 19964 24106 0 net105
rlabel metal1 36368 20434 36368 20434 0 net106
rlabel metal1 37715 20502 37715 20502 0 net107
rlabel metal1 35972 10778 35972 10778 0 net108
rlabel metal1 15502 16082 15502 16082 0 net109
rlabel metal2 30406 67371 30406 67371 0 net11
rlabel metal1 15272 16558 15272 16558 0 net110
rlabel metal1 20286 15028 20286 15028 0 net111
rlabel via1 20014 13974 20014 13974 0 net112
rlabel metal1 32798 22542 32798 22542 0 net113
rlabel metal1 33534 19754 33534 19754 0 net114
rlabel metal1 27324 14926 27324 14926 0 net115
rlabel via1 27273 13906 27273 13906 0 net116
rlabel metal1 26404 13906 26404 13906 0 net117
rlabel metal1 25300 14858 25300 14858 0 net118
rlabel metal1 25162 7378 25162 7378 0 net119
rlabel metal2 39422 68255 39422 68255 0 net12
rlabel metal1 11638 17170 11638 17170 0 net120
rlabel metal1 18354 7718 18354 7718 0 net121
rlabel metal1 30452 16150 30452 16150 0 net122
rlabel metal2 32890 20604 32890 20604 0 net123
rlabel metal2 32154 20706 32154 20706 0 net124
rlabel metal1 28336 22746 28336 22746 0 net125
rlabel metal1 36478 12274 36478 12274 0 net126
rlabel metal1 35696 24174 35696 24174 0 net127
rlabel metal2 28566 8636 28566 8636 0 net128
rlabel metal1 33810 26350 33810 26350 0 net129
rlabel metal3 751 64668 751 64668 0 net13
rlabel metal1 24104 27506 24104 27506 0 net130
rlabel metal1 22540 24922 22540 24922 0 net131
rlabel metal2 29164 12206 29164 12206 0 net132
rlabel metal1 31602 23086 31602 23086 0 net133
rlabel metal1 17204 14382 17204 14382 0 net134
rlabel metal1 17618 15130 17618 15130 0 net135
rlabel metal1 16514 23732 16514 23732 0 net136
rlabel metal1 14490 24208 14490 24208 0 net137
rlabel metal1 23230 15504 23230 15504 0 net138
rlabel via1 23133 16558 23133 16558 0 net139
rlabel metal1 33718 17544 33718 17544 0 net14
rlabel metal1 34316 9486 34316 9486 0 net140
rlabel metal1 20148 15538 20148 15538 0 net141
rlabel metal1 25024 10098 25024 10098 0 net142
rlabel metal1 27186 23630 27186 23630 0 net143
rlabel metal1 23046 25296 23046 25296 0 net144
rlabel metal1 27692 6290 27692 6290 0 net145
rlabel metal1 18354 10574 18354 10574 0 net146
rlabel metal2 12098 14518 12098 14518 0 net147
rlabel metal1 10672 23834 10672 23834 0 net148
rlabel metal1 13156 12750 13156 12750 0 net149
rlabel metal1 20608 12818 20608 12818 0 net15
rlabel metal1 23660 14994 23660 14994 0 net150
rlabel metal1 24472 23834 24472 23834 0 net151
rlabel metal1 25438 7922 25438 7922 0 net152
rlabel metal1 11040 20570 11040 20570 0 net153
rlabel metal1 9430 14246 9430 14246 0 net154
rlabel metal1 17388 9554 17388 9554 0 net155
rlabel metal2 10166 16762 10166 16762 0 net156
rlabel metal1 10994 24140 10994 24140 0 net157
rlabel metal1 20516 14858 20516 14858 0 net158
rlabel metal1 10442 22644 10442 22644 0 net159
rlabel metal1 16146 17170 16146 17170 0 net16
rlabel metal1 23092 28050 23092 28050 0 net160
rlabel metal1 37720 24174 37720 24174 0 net161
rlabel metal1 18354 9962 18354 9962 0 net162
rlabel metal1 10074 13294 10074 13294 0 net163
rlabel metal1 16560 20434 16560 20434 0 net164
rlabel metal2 24702 20740 24702 20740 0 net165
rlabel metal1 17480 16558 17480 16558 0 net166
rlabel metal2 20470 15470 20470 15470 0 net167
rlabel metal1 24288 19890 24288 19890 0 net168
rlabel metal1 36202 23154 36202 23154 0 net169
rlabel metal1 15410 17102 15410 17102 0 net17
rlabel metal1 30682 13367 30682 13367 0 net18
rlabel metal1 26542 18258 26542 18258 0 net19
rlabel metal2 68310 21658 68310 21658 0 net2
rlabel metal1 26036 18734 26036 18734 0 net20
rlabel metal1 20010 16150 20010 16150 0 net21
rlabel metal1 19228 16558 19228 16558 0 net22
rlabel metal2 20746 23596 20746 23596 0 net23
rlabel metal1 11960 18258 11960 18258 0 net24
rlabel metal1 25622 21454 25622 21454 0 net25
rlabel metal1 25760 21522 25760 21522 0 net26
rlabel metal1 17250 24174 17250 24174 0 net27
rlabel metal1 16514 24208 16514 24208 0 net28
rlabel metal1 27830 11730 27830 11730 0 net29
rlabel metal1 45540 14892 45540 14892 0 net3
rlabel metal1 21850 17646 21850 17646 0 net30
rlabel metal2 21850 16354 21850 16354 0 net31
rlabel metal1 18400 18258 18400 18258 0 net32
rlabel metal1 17357 18666 17357 18666 0 net33
rlabel metal1 14398 21522 14398 21522 0 net34
rlabel metal1 37352 21998 37352 21998 0 net35
rlabel metal1 20010 18394 20010 18394 0 net36
rlabel metal1 20792 20298 20792 20298 0 net37
rlabel metal1 19959 20842 19959 20842 0 net38
rlabel metal1 36708 17170 36708 17170 0 net39
rlabel metal2 1794 33116 1794 33116 0 net4
rlabel metal1 35558 15028 35558 15028 0 net40
rlabel metal2 19090 21641 19090 21641 0 net41
rlabel metal1 18542 20842 18542 20842 0 net42
rlabel metal1 30222 22610 30222 22610 0 net43
rlabel metal1 22356 20230 22356 20230 0 net44
rlabel metal1 28474 21114 28474 21114 0 net45
rlabel metal2 27738 21080 27738 21080 0 net46
rlabel metal1 31464 18734 31464 18734 0 net47
rlabel metal1 20194 18802 20194 18802 0 net48
rlabel metal1 26174 16524 26174 16524 0 net49
rlabel metal1 43654 2414 43654 2414 0 net5
rlabel metal1 28208 16082 28208 16082 0 net50
rlabel metal1 14720 23698 14720 23698 0 net51
rlabel metal2 17618 12517 17618 12517 0 net52
rlabel metal2 25714 24004 25714 24004 0 net53
rlabel metal1 22586 15606 22586 15606 0 net54
rlabel metal1 22555 14314 22555 14314 0 net55
rlabel metal1 32660 16014 32660 16014 0 net56
rlabel metal1 17894 13974 17894 13974 0 net57
rlabel metal1 17250 13940 17250 13940 0 net58
rlabel metal1 37812 18734 37812 18734 0 net59
rlabel metal1 12558 16150 12558 16150 0 net6
rlabel metal1 29440 26962 29440 26962 0 net60
rlabel metal1 23368 21930 23368 21930 0 net61
rlabel metal1 26450 22032 26450 22032 0 net62
rlabel metal1 16698 15062 16698 15062 0 net63
rlabel metal2 15226 14348 15226 14348 0 net64
rlabel metal1 16882 22950 16882 22950 0 net65
rlabel metal1 15226 22644 15226 22644 0 net66
rlabel metal1 33074 23766 33074 23766 0 net67
rlabel metal1 36018 20026 36018 20026 0 net68
rlabel via1 35558 19363 35558 19363 0 net69
rlabel metal2 13018 68255 13018 68255 0 net7
rlabel metal1 12282 24922 12282 24922 0 net70
rlabel metal2 23138 21828 23138 21828 0 net71
rlabel via1 23056 22678 23056 22678 0 net72
rlabel metal1 21344 8398 21344 8398 0 net73
rlabel metal1 33672 19346 33672 19346 0 net74
rlabel metal1 32890 18700 32890 18700 0 net75
rlabel via1 35190 22073 35190 22073 0 net76
rlabel metal1 29670 18598 29670 18598 0 net77
rlabel metal1 27370 26996 27370 26996 0 net78
rlabel metal1 20194 26384 20194 26384 0 net79
rlabel metal2 68494 9809 68494 9809 0 net8
rlabel metal1 27738 21930 27738 21930 0 net80
rlabel metal1 29900 17238 29900 17238 0 net81
rlabel metal1 30881 18326 30881 18326 0 net82
rlabel metal1 28014 11866 28014 11866 0 net83
rlabel metal1 30958 15062 30958 15062 0 net84
rlabel via1 33262 15062 33262 15062 0 net85
rlabel metal2 16974 22882 16974 22882 0 net86
rlabel via1 16610 21998 16610 21998 0 net87
rlabel metal1 36708 22746 36708 22746 0 net88
rlabel metal1 25346 13906 25346 13906 0 net89
rlabel metal2 26450 1027 26450 1027 0 net9
rlabel metal1 24988 13906 24988 13906 0 net90
rlabel metal1 29348 19754 29348 19754 0 net91
rlabel metal2 19642 12410 19642 12410 0 net92
rlabel metal1 21620 9622 21620 9622 0 net93
rlabel via1 27554 15011 27554 15011 0 net94
rlabel metal1 28336 14382 28336 14382 0 net95
rlabel metal1 15962 15470 15962 15470 0 net96
rlabel via1 15230 15470 15230 15470 0 net97
rlabel metal1 36248 13362 36248 13362 0 net98
rlabel metal1 34776 13498 34776 13498 0 net99
rlabel metal3 820 46308 820 46308 0 psram_ce_n
rlabel metal2 8418 2132 8418 2132 0 psram_d[0]
rlabel metal2 43838 1520 43838 1520 0 psram_sck
rlabel metal3 820 36788 820 36788 0 rst
rlabel metal1 33166 15368 33166 15368 0 softmax.addr\[11\]
rlabel metal1 32384 14790 32384 14790 0 softmax.addr\[8\]
rlabel metal1 30958 16048 30958 16048 0 softmax.data_valid
rlabel metal1 26151 12954 26151 12954 0 softmax.psram_ce_n
rlabel metal1 33534 8874 33534 8874 0 softmax.psram_ctrl.counter\[0\]
rlabel metal2 33718 9486 33718 9486 0 softmax.psram_ctrl.counter\[1\]
rlabel metal1 32522 12240 32522 12240 0 softmax.psram_ctrl.counter\[2\]
rlabel metal1 33488 9078 33488 9078 0 softmax.psram_ctrl.counter\[3\]
rlabel metal1 32982 10506 32982 10506 0 softmax.psram_ctrl.counter\[4\]
rlabel metal1 35282 12886 35282 12886 0 softmax.psram_ctrl.counter\[5\]
rlabel metal2 34178 13464 34178 13464 0 softmax.psram_ctrl.counter\[6\]
rlabel metal1 35006 12750 35006 12750 0 softmax.psram_ctrl.counter\[7\]
rlabel metal1 29486 14008 29486 14008 0 softmax.psram_ctrl.nstate
rlabel metal1 28290 12750 28290 12750 0 softmax.psram_ctrl.sck
rlabel metal1 29854 15436 29854 15436 0 softmax.psram_ctrl.start
rlabel metal1 31280 13838 31280 13838 0 softmax.psram_ctrl.state
rlabel metal2 30038 15300 30038 15300 0 softmax.start
rlabel metal1 68632 28050 68632 28050 0 start
rlabel metal1 35880 15674 35880 15674 0 state\[0\]
rlabel metal1 21942 19312 21942 19312 0 state\[1\]
rlabel metal1 34776 15470 34776 15470 0 state\[4\]
rlabel metal1 22402 13804 22402 13804 0 state\[5\]
<< properties >>
string FIXED_BBOX 0 0 70000 70000
<< end >>
