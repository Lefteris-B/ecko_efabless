VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cnn_kws_accel
  CLASS BLOCK ;
  FOREIGN cnn_kws_accel ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN audio_sample[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 346.000 0.370 350.000 ;
    END
  END audio_sample[0]
  PIN audio_sample[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 343.440 350.000 344.040 ;
    END
  END audio_sample[10]
  PIN audio_sample[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END audio_sample[11]
  PIN audio_sample[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END audio_sample[12]
  PIN audio_sample[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END audio_sample[13]
  PIN audio_sample[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 346.000 216.110 350.000 ;
    END
  END audio_sample[14]
  PIN audio_sample[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 346.000 332.030 350.000 ;
    END
  END audio_sample[15]
  PIN audio_sample[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 346.000 254.750 350.000 ;
    END
  END audio_sample[1]
  PIN audio_sample[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END audio_sample[2]
  PIN audio_sample[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 346.000 177.470 350.000 ;
    END
  END audio_sample[3]
  PIN audio_sample[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END audio_sample[4]
  PIN audio_sample[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 193.840 350.000 194.440 ;
    END
  END audio_sample[5]
  PIN audio_sample[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END audio_sample[6]
  PIN audio_sample[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END audio_sample[7]
  PIN audio_sample[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 346.000 241.870 350.000 ;
    END
  END audio_sample[8]
  PIN audio_sample[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END audio_sample[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 302.640 350.000 303.240 ;
    END
  END done
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 112.240 350.000 112.840 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 289.040 350.000 289.640 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 346.000 293.390 350.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 71.440 350.000 72.040 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 329.840 350.000 330.440 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 57.840 350.000 58.440 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 346.000 100.190 350.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 346.000 190.350 350.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 346.000 319.150 350.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 261.840 350.000 262.440 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 17.040 350.000 17.640 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 153.040 350.000 153.640 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 125.840 350.000 126.440 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 346.000 113.070 350.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 346.000 125.950 350.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 275.440 350.000 276.040 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 44.240 350.000 44.840 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 3.440 350.000 4.040 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 180.240 350.000 180.840 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 346.000 138.830 350.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 316.240 350.000 316.840 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 346.000 164.590 350.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 85.040 350.000 85.640 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 221.040 350.000 221.640 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 346.000 203.230 350.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 346.000 87.310 350.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 98.640 350.000 99.240 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 139.440 350.000 140.040 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 234.640 350.000 235.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 248.240 350.000 248.840 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 346.000 35.790 350.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 346.000 48.670 350.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 346.000 61.550 350.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 346.000 151.710 350.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 346.000 306.270 350.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 346.000 228.990 350.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 346.000 344.910 350.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 30.640 350.000 31.240 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 346.000 10.030 350.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END io_out[9]
  PIN psram_ce_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END psram_ce_n
  PIN psram_d[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END psram_d[0]
  PIN psram_d[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END psram_d[1]
  PIN psram_d[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 207.440 350.000 208.040 ;
    END
  END psram_d[2]
  PIN psram_d[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END psram_d[3]
  PIN psram_douten[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 346.000 280.510 350.000 ;
    END
  END psram_douten[0]
  PIN psram_douten[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 346.000 267.630 350.000 ;
    END
  END psram_douten[1]
  PIN psram_douten[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 346.000 22.910 350.000 ;
    END
  END psram_douten[2]
  PIN psram_douten[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 346.000 74.430 350.000 ;
    END
  END psram_douten[3]
  PIN psram_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END psram_sck
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END rst
  PIN sample_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END sample_valid
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 346.000 166.640 350.000 167.240 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 0.070 10.640 344.930 337.520 ;
      LAYER met2 ;
        RECT 0.650 345.720 9.470 346.530 ;
        RECT 10.310 345.720 22.350 346.530 ;
        RECT 23.190 345.720 35.230 346.530 ;
        RECT 36.070 345.720 48.110 346.530 ;
        RECT 48.950 345.720 60.990 346.530 ;
        RECT 61.830 345.720 73.870 346.530 ;
        RECT 74.710 345.720 86.750 346.530 ;
        RECT 87.590 345.720 99.630 346.530 ;
        RECT 100.470 345.720 112.510 346.530 ;
        RECT 113.350 345.720 125.390 346.530 ;
        RECT 126.230 345.720 138.270 346.530 ;
        RECT 139.110 345.720 151.150 346.530 ;
        RECT 151.990 345.720 164.030 346.530 ;
        RECT 164.870 345.720 176.910 346.530 ;
        RECT 177.750 345.720 189.790 346.530 ;
        RECT 190.630 345.720 202.670 346.530 ;
        RECT 203.510 345.720 215.550 346.530 ;
        RECT 216.390 345.720 228.430 346.530 ;
        RECT 229.270 345.720 241.310 346.530 ;
        RECT 242.150 345.720 254.190 346.530 ;
        RECT 255.030 345.720 267.070 346.530 ;
        RECT 267.910 345.720 279.950 346.530 ;
        RECT 280.790 345.720 292.830 346.530 ;
        RECT 293.670 345.720 305.710 346.530 ;
        RECT 306.550 345.720 318.590 346.530 ;
        RECT 319.430 345.720 331.470 346.530 ;
        RECT 332.310 345.720 344.350 346.530 ;
        RECT 0.100 4.280 344.900 345.720 ;
        RECT 0.650 3.555 9.470 4.280 ;
        RECT 10.310 3.555 22.350 4.280 ;
        RECT 23.190 3.555 35.230 4.280 ;
        RECT 36.070 3.555 48.110 4.280 ;
        RECT 48.950 3.555 60.990 4.280 ;
        RECT 61.830 3.555 73.870 4.280 ;
        RECT 74.710 3.555 86.750 4.280 ;
        RECT 87.590 3.555 99.630 4.280 ;
        RECT 100.470 3.555 112.510 4.280 ;
        RECT 113.350 3.555 125.390 4.280 ;
        RECT 126.230 3.555 138.270 4.280 ;
        RECT 139.110 3.555 151.150 4.280 ;
        RECT 151.990 3.555 164.030 4.280 ;
        RECT 164.870 3.555 176.910 4.280 ;
        RECT 177.750 3.555 189.790 4.280 ;
        RECT 190.630 3.555 202.670 4.280 ;
        RECT 203.510 3.555 215.550 4.280 ;
        RECT 216.390 3.555 228.430 4.280 ;
        RECT 229.270 3.555 241.310 4.280 ;
        RECT 242.150 3.555 254.190 4.280 ;
        RECT 255.030 3.555 267.070 4.280 ;
        RECT 267.910 3.555 279.950 4.280 ;
        RECT 280.790 3.555 292.830 4.280 ;
        RECT 293.670 3.555 305.710 4.280 ;
        RECT 306.550 3.555 318.590 4.280 ;
        RECT 319.430 3.555 331.470 4.280 ;
        RECT 332.310 3.555 341.130 4.280 ;
        RECT 341.970 3.555 344.900 4.280 ;
      LAYER met3 ;
        RECT 4.400 336.240 346.000 337.445 ;
        RECT 3.990 330.840 346.000 336.240 ;
        RECT 3.990 329.440 345.600 330.840 ;
        RECT 3.990 324.040 346.000 329.440 ;
        RECT 4.400 322.640 346.000 324.040 ;
        RECT 3.990 317.240 346.000 322.640 ;
        RECT 3.990 315.840 345.600 317.240 ;
        RECT 3.990 310.440 346.000 315.840 ;
        RECT 4.400 309.040 346.000 310.440 ;
        RECT 3.990 303.640 346.000 309.040 ;
        RECT 3.990 302.240 345.600 303.640 ;
        RECT 3.990 296.840 346.000 302.240 ;
        RECT 4.400 295.440 346.000 296.840 ;
        RECT 3.990 290.040 346.000 295.440 ;
        RECT 3.990 288.640 345.600 290.040 ;
        RECT 3.990 283.240 346.000 288.640 ;
        RECT 4.400 281.840 346.000 283.240 ;
        RECT 3.990 276.440 346.000 281.840 ;
        RECT 3.990 275.040 345.600 276.440 ;
        RECT 3.990 269.640 346.000 275.040 ;
        RECT 4.400 268.240 346.000 269.640 ;
        RECT 3.990 262.840 346.000 268.240 ;
        RECT 3.990 261.440 345.600 262.840 ;
        RECT 3.990 256.040 346.000 261.440 ;
        RECT 4.400 254.640 346.000 256.040 ;
        RECT 3.990 249.240 346.000 254.640 ;
        RECT 3.990 247.840 345.600 249.240 ;
        RECT 3.990 242.440 346.000 247.840 ;
        RECT 4.400 241.040 346.000 242.440 ;
        RECT 3.990 235.640 346.000 241.040 ;
        RECT 3.990 234.240 345.600 235.640 ;
        RECT 3.990 228.840 346.000 234.240 ;
        RECT 4.400 227.440 346.000 228.840 ;
        RECT 3.990 222.040 346.000 227.440 ;
        RECT 3.990 220.640 345.600 222.040 ;
        RECT 3.990 215.240 346.000 220.640 ;
        RECT 4.400 213.840 346.000 215.240 ;
        RECT 3.990 208.440 346.000 213.840 ;
        RECT 3.990 207.040 345.600 208.440 ;
        RECT 3.990 201.640 346.000 207.040 ;
        RECT 4.400 200.240 346.000 201.640 ;
        RECT 3.990 194.840 346.000 200.240 ;
        RECT 3.990 193.440 345.600 194.840 ;
        RECT 3.990 188.040 346.000 193.440 ;
        RECT 4.400 186.640 346.000 188.040 ;
        RECT 3.990 181.240 346.000 186.640 ;
        RECT 3.990 179.840 345.600 181.240 ;
        RECT 3.990 174.440 346.000 179.840 ;
        RECT 4.400 173.040 346.000 174.440 ;
        RECT 3.990 167.640 346.000 173.040 ;
        RECT 3.990 166.240 345.600 167.640 ;
        RECT 3.990 160.840 346.000 166.240 ;
        RECT 4.400 159.440 346.000 160.840 ;
        RECT 3.990 154.040 346.000 159.440 ;
        RECT 3.990 152.640 345.600 154.040 ;
        RECT 3.990 147.240 346.000 152.640 ;
        RECT 4.400 145.840 346.000 147.240 ;
        RECT 3.990 140.440 346.000 145.840 ;
        RECT 3.990 139.040 345.600 140.440 ;
        RECT 3.990 133.640 346.000 139.040 ;
        RECT 4.400 132.240 346.000 133.640 ;
        RECT 3.990 126.840 346.000 132.240 ;
        RECT 3.990 125.440 345.600 126.840 ;
        RECT 3.990 120.040 346.000 125.440 ;
        RECT 4.400 118.640 346.000 120.040 ;
        RECT 3.990 113.240 346.000 118.640 ;
        RECT 3.990 111.840 345.600 113.240 ;
        RECT 3.990 106.440 346.000 111.840 ;
        RECT 4.400 105.040 346.000 106.440 ;
        RECT 3.990 99.640 346.000 105.040 ;
        RECT 3.990 98.240 345.600 99.640 ;
        RECT 3.990 92.840 346.000 98.240 ;
        RECT 4.400 91.440 346.000 92.840 ;
        RECT 3.990 86.040 346.000 91.440 ;
        RECT 3.990 84.640 345.600 86.040 ;
        RECT 3.990 79.240 346.000 84.640 ;
        RECT 4.400 77.840 346.000 79.240 ;
        RECT 3.990 72.440 346.000 77.840 ;
        RECT 3.990 71.040 345.600 72.440 ;
        RECT 3.990 65.640 346.000 71.040 ;
        RECT 4.400 64.240 346.000 65.640 ;
        RECT 3.990 58.840 346.000 64.240 ;
        RECT 3.990 57.440 345.600 58.840 ;
        RECT 3.990 52.040 346.000 57.440 ;
        RECT 4.400 50.640 346.000 52.040 ;
        RECT 3.990 45.240 346.000 50.640 ;
        RECT 3.990 43.840 345.600 45.240 ;
        RECT 3.990 38.440 346.000 43.840 ;
        RECT 4.400 37.040 346.000 38.440 ;
        RECT 3.990 31.640 346.000 37.040 ;
        RECT 3.990 30.240 345.600 31.640 ;
        RECT 3.990 24.840 346.000 30.240 ;
        RECT 4.400 23.440 346.000 24.840 ;
        RECT 3.990 18.040 346.000 23.440 ;
        RECT 3.990 16.640 345.600 18.040 ;
        RECT 3.990 11.240 346.000 16.640 ;
        RECT 4.400 9.840 346.000 11.240 ;
        RECT 3.990 4.440 346.000 9.840 ;
        RECT 3.990 3.575 345.600 4.440 ;
      LAYER met4 ;
        RECT 187.975 16.495 188.305 69.185 ;
  END
END cnn_kws_accel
END LIBRARY

