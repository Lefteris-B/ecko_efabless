// This is the unpowered netlist.
module cnn_kws_accel (clk,
    done,
    psram_ce_n,
    psram_sck,
    rst_n,
    sample_valid,
    start,
    audio_sample,
    psram_d,
    psram_douten);
 input clk;
 output done;
 output psram_ce_n;
 output psram_sck;
 input rst_n;
 input sample_valid;
 input start;
 input [15:0] audio_sample;
 inout [3:0] psram_d;
 output [3:0] psram_douten;

 wire net23;
 wire net24;
 wire net25;
 wire net29;
 wire net26;
 wire net27;
 wire net28;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire \conv1.addr[8] ;
 wire \conv1.done ;
 wire \conv1.psram_ce_n ;
 wire \conv1.psram_ctrl.counter[0] ;
 wire \conv1.psram_ctrl.counter[1] ;
 wire \conv1.psram_ctrl.counter[2] ;
 wire \conv1.psram_ctrl.counter[3] ;
 wire \conv1.psram_ctrl.counter[4] ;
 wire \conv1.psram_ctrl.counter[5] ;
 wire \conv1.psram_ctrl.counter[6] ;
 wire \conv1.psram_ctrl.counter[7] ;
 wire \conv1.psram_ctrl.has_wait_states ;
 wire \conv1.psram_ctrl.nstate ;
 wire \conv1.psram_ctrl.sck ;
 wire \conv1.psram_ctrl.start ;
 wire \conv1.psram_ctrl.state ;
 wire \conv1.state[0] ;
 wire \conv1.state[1] ;
 wire \conv1.state[2] ;
 wire \conv1.state[3] ;
 wire \conv1.state[5] ;
 wire \conv2.addr[8] ;
 wire \conv2.addr[9] ;
 wire \conv2.data_out_valid ;
 wire \conv2.psram_ce_n ;
 wire \conv2.psram_ctrl.counter[0] ;
 wire \conv2.psram_ctrl.counter[1] ;
 wire \conv2.psram_ctrl.counter[2] ;
 wire \conv2.psram_ctrl.counter[3] ;
 wire \conv2.psram_ctrl.counter[4] ;
 wire \conv2.psram_ctrl.counter[5] ;
 wire \conv2.psram_ctrl.counter[6] ;
 wire \conv2.psram_ctrl.counter[7] ;
 wire \conv2.psram_ctrl.has_wait_states ;
 wire \conv2.psram_ctrl.nstate ;
 wire \conv2.psram_ctrl.sck ;
 wire \conv2.psram_ctrl.start ;
 wire \conv2.psram_ctrl.state ;
 wire \conv2.state[0] ;
 wire \conv2.state[1] ;
 wire \conv2.state[2] ;
 wire \conv2.state[3] ;
 wire \conv2.state[5] ;
 wire \fc1.addr[10] ;
 wire \fc1.addr[8] ;
 wire \fc1.data_out_valid ;
 wire \fc1.psram_ce_n ;
 wire \fc1.psram_ctrl.counter[0] ;
 wire \fc1.psram_ctrl.counter[1] ;
 wire \fc1.psram_ctrl.counter[2] ;
 wire \fc1.psram_ctrl.counter[3] ;
 wire \fc1.psram_ctrl.counter[4] ;
 wire \fc1.psram_ctrl.counter[5] ;
 wire \fc1.psram_ctrl.counter[6] ;
 wire \fc1.psram_ctrl.counter[7] ;
 wire \fc1.psram_ctrl.has_wait_states ;
 wire \fc1.psram_ctrl.nstate ;
 wire \fc1.psram_ctrl.sck ;
 wire \fc1.psram_ctrl.start ;
 wire \fc1.psram_ctrl.state ;
 wire \fc1.state[0] ;
 wire \fc1.state[1] ;
 wire \fc1.state[2] ;
 wire \fc1.state[3] ;
 wire \fc1.state[5] ;
 wire \fc2.addr[10] ;
 wire \fc2.addr[8] ;
 wire \fc2.done ;
 wire \fc2.psram_ce_n ;
 wire \fc2.psram_ctrl.counter[0] ;
 wire \fc2.psram_ctrl.counter[1] ;
 wire \fc2.psram_ctrl.counter[2] ;
 wire \fc2.psram_ctrl.counter[3] ;
 wire \fc2.psram_ctrl.counter[4] ;
 wire \fc2.psram_ctrl.counter[5] ;
 wire \fc2.psram_ctrl.counter[6] ;
 wire \fc2.psram_ctrl.counter[7] ;
 wire \fc2.psram_ctrl.has_wait_states ;
 wire \fc2.psram_ctrl.nstate ;
 wire \fc2.psram_ctrl.sck ;
 wire \fc2.psram_ctrl.start ;
 wire \fc2.psram_ctrl.state ;
 wire \fc2.state[0] ;
 wire \fc2.state[1] ;
 wire \fc2.state[2] ;
 wire \fc2.state[3] ;
 wire \fc2.state[5] ;
 wire \maxpool.addr[11] ;
 wire \maxpool.addr[8] ;
 wire \maxpool.psram_ce_n ;
 wire \maxpool.psram_ctrl.counter[0] ;
 wire \maxpool.psram_ctrl.counter[1] ;
 wire \maxpool.psram_ctrl.counter[2] ;
 wire \maxpool.psram_ctrl.counter[3] ;
 wire \maxpool.psram_ctrl.counter[4] ;
 wire \maxpool.psram_ctrl.counter[5] ;
 wire \maxpool.psram_ctrl.counter[6] ;
 wire \maxpool.psram_ctrl.counter[7] ;
 wire \maxpool.psram_ctrl.nstate ;
 wire \maxpool.psram_ctrl.sck ;
 wire \maxpool.psram_ctrl.start ;
 wire \maxpool.psram_ctrl.state ;
 wire \maxpool.state[0] ;
 wire \maxpool.state[1] ;
 wire \maxpool.state[2] ;
 wire \mfcc.dct.data_valid ;
 wire \mfcc.dct.dct_valid ;
 wire \mfcc.dct.input_counter[0] ;
 wire \mfcc.dct.input_counter[1] ;
 wire \mfcc.dct.input_counter[2] ;
 wire \mfcc.dct.input_counter[3] ;
 wire \mfcc.dct.input_counter[4] ;
 wire \mfcc.dct.output_counter[0] ;
 wire \mfcc.dct.output_counter[1] ;
 wire \mfcc.dct.output_counter[2] ;
 wire \mfcc.dct.output_counter[3] ;
 wire \mfcc.dct.output_counter[4] ;
 wire \mfcc.dct.output_counter[5] ;
 wire \mfcc.dct.state[0] ;
 wire \mfcc.dct.state[1] ;
 wire \mfcc.log.data_valid ;
 wire \mfcc.log.shift_count[0] ;
 wire \mfcc.log.shift_count[1] ;
 wire \mfcc.log.shift_count[2] ;
 wire \mfcc.log.shift_count[3] ;
 wire \mfcc.log.state[0] ;
 wire \mfcc.log.state[1] ;
 wire \mfcc.log.state[2] ;
 wire \mfcc.mel.coeff_counter[0] ;
 wire \mfcc.mel.coeff_counter[1] ;
 wire \mfcc.mel.coeff_counter[2] ;
 wire \mfcc.mel.coeff_counter[3] ;
 wire \mfcc.mel.coeff_counter[4] ;
 wire \mfcc.mel.filter_counter[0] ;
 wire \mfcc.mel.filter_counter[1] ;
 wire \mfcc.mel.filter_counter[2] ;
 wire \mfcc.mel.filter_counter[3] ;
 wire \mfcc.mel.filter_counter[4] ;
 wire \mfcc.mel.filter_counter[5] ;
 wire \mfcc.mel.state[0] ;
 wire \mfcc.mel.state[1] ;
 wire \mfcc.mfcc_valid ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \softmax.addr[11] ;
 wire \softmax.addr[8] ;
 wire \softmax.data_valid ;
 wire \softmax.psram_ce_n ;
 wire \softmax.psram_ctrl.counter[0] ;
 wire \softmax.psram_ctrl.counter[1] ;
 wire \softmax.psram_ctrl.counter[2] ;
 wire \softmax.psram_ctrl.counter[3] ;
 wire \softmax.psram_ctrl.counter[4] ;
 wire \softmax.psram_ctrl.counter[5] ;
 wire \softmax.psram_ctrl.counter[6] ;
 wire \softmax.psram_ctrl.counter[7] ;
 wire \softmax.psram_ctrl.nstate ;
 wire \softmax.psram_ctrl.sck ;
 wire \softmax.psram_ctrl.start ;
 wire \softmax.psram_ctrl.state ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;

 sky130_fd_sc_hd__decap_8 FILLER_0_0_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_80 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__or3_1 _0521_ (.A(\fc2.state[2] ),
    .B(\fc2.state[1] ),
    .C(\fc2.state[3] ),
    .X(_0149_));
 sky130_fd_sc_hd__buf_1 _0522_ (.A(_0149_),
    .X(_0028_));
 sky130_fd_sc_hd__or3b_1 _0523_ (.A(\state[2] ),
    .B(\state[0] ),
    .C_N(\state[1] ),
    .X(_0150_));
 sky130_fd_sc_hd__buf_2 _0524_ (.A(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__a21o_1 _0525_ (.A1(\conv1.state[0] ),
    .A2(_0151_),
    .B1(net55),
    .X(_0010_));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(\fc2.psram_ctrl.has_wait_states ),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _0527_ (.A(\fc2.psram_ctrl.counter[4] ),
    .Y(_0153_));
 sky130_fd_sc_hd__or3b_1 _0528_ (.A(_0153_),
    .B(\fc2.psram_ctrl.counter[2] ),
    .C_N(\fc2.psram_ctrl.counter[5] ),
    .X(_0154_));
 sky130_fd_sc_hd__or2_1 _0529_ (.A(\fc2.psram_ctrl.counter[1] ),
    .B(\fc2.psram_ctrl.counter[0] ),
    .X(_0155_));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(\fc2.psram_ctrl.counter[3] ),
    .Y(_0156_));
 sky130_fd_sc_hd__a211o_1 _0531_ (.A1(\fc2.psram_ctrl.has_wait_states ),
    .A2(_0156_),
    .B1(\fc2.psram_ctrl.counter[7] ),
    .C1(\fc2.psram_ctrl.counter[6] ),
    .X(_0157_));
 sky130_fd_sc_hd__a2111o_4 _0532_ (.A1(_0152_),
    .A2(\fc2.psram_ctrl.counter[3] ),
    .B1(_0154_),
    .C1(_0155_),
    .D1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__a21o_1 _0533_ (.A1(\fc2.state[1] ),
    .A2(_0158_),
    .B1(net38),
    .X(_0020_));
 sky130_fd_sc_hd__inv_2 _0534_ (.A(\fc1.data_out_valid ),
    .Y(_0159_));
 sky130_fd_sc_hd__a21o_1 _0535_ (.A1(\fc2.state[0] ),
    .A2(_0159_),
    .B1(net45),
    .X(_0019_));
 sky130_fd_sc_hd__or3_1 _0536_ (.A(\fc1.state[2] ),
    .B(\fc1.state[3] ),
    .C(\fc1.state[1] ),
    .X(_0160_));
 sky130_fd_sc_hd__buf_1 _0537_ (.A(_0160_),
    .X(_0029_));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(\conv2.psram_ctrl.counter[4] ),
    .Y(_0161_));
 sky130_fd_sc_hd__or3b_1 _0539_ (.A(_0161_),
    .B(\conv2.psram_ctrl.counter[2] ),
    .C_N(\conv2.psram_ctrl.counter[5] ),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _0540_ (.A(\conv2.psram_ctrl.counter[1] ),
    .B(\conv2.psram_ctrl.counter[0] ),
    .X(_0163_));
 sky130_fd_sc_hd__or2_1 _0541_ (.A(\conv2.psram_ctrl.counter[7] ),
    .B(\conv2.psram_ctrl.counter[6] ),
    .X(_0164_));
 sky130_fd_sc_hd__xor2_1 _0542_ (.A(\conv2.psram_ctrl.has_wait_states ),
    .B(\conv2.psram_ctrl.counter[3] ),
    .X(_0165_));
 sky130_fd_sc_hd__or4_1 _0543_ (.A(_0162_),
    .B(_0163_),
    .C(_0164_),
    .D(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__buf_2 _0544_ (.A(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__nand2_1 _0545_ (.A(\state[0] ),
    .B(\state[1] ),
    .Y(_0168_));
 sky130_fd_sc_hd__nor2_1 _0546_ (.A(\state[2] ),
    .B(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hd__a22o_1 _0547_ (.A1(net74),
    .A2(_0167_),
    .B1(_0169_),
    .B2(net129),
    .X(_0015_));
 sky130_fd_sc_hd__inv_2 _0548_ (.A(_0151_),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _0549_ (.A(\conv1.psram_ctrl.counter[4] ),
    .Y(_0171_));
 sky130_fd_sc_hd__or3b_1 _0550_ (.A(\conv1.psram_ctrl.counter[2] ),
    .B(_0171_),
    .C_N(\conv1.psram_ctrl.counter[5] ),
    .X(_0172_));
 sky130_fd_sc_hd__or2_1 _0551_ (.A(\conv1.psram_ctrl.counter[1] ),
    .B(\conv1.psram_ctrl.counter[0] ),
    .X(_0173_));
 sky130_fd_sc_hd__or2_1 _0552_ (.A(\conv1.psram_ctrl.counter[7] ),
    .B(\conv1.psram_ctrl.counter[6] ),
    .X(_0174_));
 sky130_fd_sc_hd__xor2_1 _0553_ (.A(\conv1.psram_ctrl.has_wait_states ),
    .B(\conv1.psram_ctrl.counter[3] ),
    .X(_0175_));
 sky130_fd_sc_hd__or4_1 _0554_ (.A(_0172_),
    .B(_0173_),
    .C(_0174_),
    .D(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__buf_2 _0555_ (.A(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_1 _0556_ (.A1(\conv1.state[0] ),
    .A2(_0170_),
    .B1(_0177_),
    .B2(net147),
    .X(_0012_));
 sky130_fd_sc_hd__a22o_1 _0557_ (.A1(\fc2.state[0] ),
    .A2(\fc1.data_out_valid ),
    .B1(_0158_),
    .B2(net70),
    .X(_0021_));
 sky130_fd_sc_hd__a21o_1 _0558_ (.A1(\conv1.state[1] ),
    .A2(_0177_),
    .B1(net40),
    .X(_0011_));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(\fc1.psram_ctrl.counter[2] ),
    .Y(_0178_));
 sky130_fd_sc_hd__nand3_1 _0560_ (.A(_0178_),
    .B(\fc1.psram_ctrl.counter[5] ),
    .C(\fc1.psram_ctrl.counter[4] ),
    .Y(_0179_));
 sky130_fd_sc_hd__xor2_1 _0561_ (.A(\fc1.psram_ctrl.has_wait_states ),
    .B(\fc1.psram_ctrl.counter[3] ),
    .X(_0180_));
 sky130_fd_sc_hd__or2_1 _0562_ (.A(\fc1.psram_ctrl.counter[7] ),
    .B(\fc1.psram_ctrl.counter[6] ),
    .X(_0181_));
 sky130_fd_sc_hd__or2_1 _0563_ (.A(\fc1.psram_ctrl.counter[1] ),
    .B(\fc1.psram_ctrl.counter[0] ),
    .X(_0182_));
 sky130_fd_sc_hd__or4_1 _0564_ (.A(_0179_),
    .B(_0180_),
    .C(_0181_),
    .D(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__buf_2 _0565_ (.A(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__a22o_1 _0566_ (.A1(net79),
    .A2(net108),
    .B1(_0184_),
    .B2(net106),
    .X(_0018_));
 sky130_fd_sc_hd__nor3b_2 _0567_ (.A(\mfcc.dct.output_counter[4] ),
    .B(\mfcc.dct.output_counter[3] ),
    .C_N(\mfcc.dct.output_counter[5] ),
    .Y(_0185_));
 sky130_fd_sc_hd__and3_1 _0568_ (.A(\mfcc.dct.input_counter[4] ),
    .B(\mfcc.dct.input_counter[3] ),
    .C(\mfcc.dct.input_counter[0] ),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _0569_ (.A(\mfcc.dct.input_counter[2] ),
    .B(\mfcc.dct.input_counter[1] ),
    .C(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_2 _0570_ (.A(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__and4_1 _0571_ (.A(\mfcc.dct.output_counter[1] ),
    .B(\mfcc.dct.output_counter[0] ),
    .C(\mfcc.dct.state[1] ),
    .D(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _0572_ (.A(\mfcc.dct.output_counter[2] ),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__buf_2 _0573_ (.A(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__nand2_1 _0574_ (.A(\mfcc.dct.data_valid ),
    .B(_0188_),
    .Y(_0192_));
 sky130_fd_sc_hd__clkbuf_4 _0575_ (.A(net21),
    .X(_0193_));
 sky130_fd_sc_hd__a221o_1 _0576_ (.A1(_0185_),
    .A2(_0191_),
    .B1(_0192_),
    .B2(net98),
    .C1(_0193_),
    .X(_0022_));
 sky130_fd_sc_hd__inv_2 _0577_ (.A(\mfcc.log.data_valid ),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _0578_ (.A(\mfcc.log.state[1] ),
    .Y(_0195_));
 sky130_fd_sc_hd__nand4_1 _0579_ (.A(\mfcc.log.shift_count[3] ),
    .B(\mfcc.log.shift_count[2] ),
    .C(\mfcc.log.shift_count[1] ),
    .D(\mfcc.log.shift_count[0] ),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _0580_ (.A(_0195_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__a2111o_1 _0581_ (.A1(_0194_),
    .A2(net53),
    .B1(\mfcc.log.state[2] ),
    .C1(_0197_),
    .D1(_0193_),
    .X(_0024_));
 sky130_fd_sc_hd__inv_2 _0582_ (.A(net20),
    .Y(_0198_));
 sky130_fd_sc_hd__clkbuf_4 _0583_ (.A(_0198_),
    .X(_0038_));
 sky130_fd_sc_hd__and4_1 _0584_ (.A(\mfcc.dct.output_counter[2] ),
    .B(\mfcc.dct.output_counter[1] ),
    .C(\mfcc.dct.output_counter[0] ),
    .D(_0185_),
    .X(_0199_));
 sky130_fd_sc_hd__nand2_1 _0585_ (.A(_0188_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__a32o_1 _0586_ (.A1(\mfcc.dct.data_valid ),
    .A2(\mfcc.dct.state[0] ),
    .A3(_0188_),
    .B1(_0200_),
    .B2(\mfcc.dct.state[1] ),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _0587_ (.A(_0038_),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_1 _0588_ (.A(_0202_),
    .X(_0023_));
 sky130_fd_sc_hd__or3_1 _0589_ (.A(\conv2.state[3] ),
    .B(\conv2.state[2] ),
    .C(\conv2.state[1] ),
    .X(_0203_));
 sky130_fd_sc_hd__buf_1 _0590_ (.A(_0203_),
    .X(_0030_));
 sky130_fd_sc_hd__and3b_1 _0591_ (.A_N(\mfcc.mel.coeff_counter[0] ),
    .B(\mfcc.mel.coeff_counter[1] ),
    .C(\mfcc.mel.coeff_counter[2] ),
    .X(_0204_));
 sky130_fd_sc_hd__and3b_1 _0592_ (.A_N(\mfcc.mel.coeff_counter[3] ),
    .B(_0204_),
    .C(\mfcc.mel.coeff_counter[4] ),
    .X(_0205_));
 sky130_fd_sc_hd__or4b_1 _0593_ (.A(\mfcc.mel.filter_counter[2] ),
    .B(\mfcc.mel.filter_counter[1] ),
    .C(\mfcc.mel.filter_counter[0] ),
    .D_N(\mfcc.mel.filter_counter[3] ),
    .X(_0206_));
 sky130_fd_sc_hd__nor3b_1 _0594_ (.A(\mfcc.mel.filter_counter[4] ),
    .B(_0206_),
    .C_N(\mfcc.mel.filter_counter[5] ),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _0595_ (.A(_0205_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__and3_1 _0596_ (.A(\mfcc.mel.state[1] ),
    .B(_0198_),
    .C(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0209_),
    .X(_0026_));
 sky130_fd_sc_hd__and2_2 _0598_ (.A(\mfcc.mel.state[1] ),
    .B(_0205_),
    .X(_0210_));
 sky130_fd_sc_hd__a211o_1 _0599_ (.A1(_0207_),
    .A2(_0210_),
    .B1(_0193_),
    .C1(net48),
    .X(_0025_));
 sky130_fd_sc_hd__or2_2 _0600_ (.A(\state[2] ),
    .B(_0168_),
    .X(_0211_));
 sky130_fd_sc_hd__a21o_1 _0601_ (.A1(\conv2.state[0] ),
    .A2(_0211_),
    .B1(net79),
    .X(_0013_));
 sky130_fd_sc_hd__a21o_1 _0602_ (.A1(\fc1.state[1] ),
    .A2(_0184_),
    .B1(net36),
    .X(_0017_));
 sky130_fd_sc_hd__inv_2 _0603_ (.A(\conv2.data_out_valid ),
    .Y(_0212_));
 sky130_fd_sc_hd__a21o_1 _0604_ (.A1(_0212_),
    .A2(net108),
    .B1(net111),
    .X(_0016_));
 sky130_fd_sc_hd__a21o_1 _0605_ (.A1(\conv2.state[1] ),
    .A2(_0167_),
    .B1(net34),
    .X(_0014_));
 sky130_fd_sc_hd__inv_2 _0606_ (.A(net58),
    .Y(_0213_));
 sky130_fd_sc_hd__and2_1 _0607_ (.A(_0213_),
    .B(\maxpool.state[0] ),
    .X(_0214_));
 sky130_fd_sc_hd__buf_1 _0608_ (.A(_0214_),
    .X(_0027_));
 sky130_fd_sc_hd__or3_1 _0609_ (.A(\conv1.state[3] ),
    .B(\conv1.state[1] ),
    .C(\conv1.state[2] ),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_1 _0610_ (.A(_0215_),
    .X(_0031_));
 sky130_fd_sc_hd__nand3_2 _0611_ (.A(\state[2] ),
    .B(\state[0] ),
    .C(\state[1] ),
    .Y(_0216_));
 sky130_fd_sc_hd__or3b_1 _0612_ (.A(\softmax.psram_ctrl.counter[7] ),
    .B(\softmax.psram_ctrl.counter[3] ),
    .C_N(\softmax.psram_ctrl.counter[4] ),
    .X(_0217_));
 sky130_fd_sc_hd__or2_1 _0613_ (.A(\softmax.psram_ctrl.counter[1] ),
    .B(\softmax.psram_ctrl.counter[0] ),
    .X(_0218_));
 sky130_fd_sc_hd__or3b_1 _0614_ (.A(\softmax.psram_ctrl.counter[6] ),
    .B(\softmax.psram_ctrl.counter[2] ),
    .C_N(\softmax.psram_ctrl.counter[5] ),
    .X(_0219_));
 sky130_fd_sc_hd__or3_1 _0615_ (.A(_0217_),
    .B(_0218_),
    .C(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__buf_2 _0616_ (.A(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__nor3_1 _0617_ (.A(\softmax.data_valid ),
    .B(\softmax.psram_ctrl.start ),
    .C(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__mux2_1 _0618_ (.A0(net2),
    .A1(\mfcc.mfcc_valid ),
    .S(\state[0] ),
    .X(_0223_));
 sky130_fd_sc_hd__or2b_1 _0619_ (.A(\state[1] ),
    .B_N(\state[2] ),
    .X(_0224_));
 sky130_fd_sc_hd__or2_2 _0620_ (.A(\state[0] ),
    .B(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__o32a_1 _0621_ (.A1(\state[2] ),
    .A2(\state[1] ),
    .A3(_0223_),
    .B1(_0225_),
    .B2(\fc1.data_out_valid ),
    .X(_0226_));
 sky130_fd_sc_hd__inv_2 _0622_ (.A(\state[0] ),
    .Y(_0227_));
 sky130_fd_sc_hd__or2_1 _0623_ (.A(_0227_),
    .B(_0224_),
    .X(_0228_));
 sky130_fd_sc_hd__and3b_2 _0624_ (.A_N(\state[0] ),
    .B(\state[1] ),
    .C(\state[2] ),
    .X(_0229_));
 sky130_fd_sc_hd__or3b_1 _0625_ (.A(\maxpool.state[0] ),
    .B(\maxpool.state[1] ),
    .C_N(\maxpool.state[2] ),
    .X(_0230_));
 sky130_fd_sc_hd__o2bb2a_1 _0626_ (.A1_N(_0229_),
    .A2_N(_0230_),
    .B1(\conv1.done ),
    .B2(_0151_),
    .X(_0231_));
 sky130_fd_sc_hd__o221a_1 _0627_ (.A1(\conv2.data_out_valid ),
    .A2(_0211_),
    .B1(_0228_),
    .B2(\fc2.done ),
    .C1(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__o211ai_2 _0628_ (.A1(_0216_),
    .A2(_0222_),
    .B1(_0226_),
    .C1(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__nor2_1 _0629_ (.A(_0216_),
    .B(_0233_),
    .Y(net3));
 sky130_fd_sc_hd__nor2_1 _0630_ (.A(_0227_),
    .B(_0224_),
    .Y(_0234_));
 sky130_fd_sc_hd__mux2_1 _0631_ (.A0(\softmax.psram_ctrl.sck ),
    .A1(\maxpool.psram_ctrl.sck ),
    .S(_0229_),
    .X(_0235_));
 sky130_fd_sc_hd__inv_2 _0632_ (.A(\fc1.psram_ctrl.sck ),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _0633_ (.A(_0236_),
    .B(_0225_),
    .Y(_0237_));
 sky130_fd_sc_hd__a221o_1 _0634_ (.A1(\fc2.psram_ctrl.sck ),
    .A2(_0234_),
    .B1(_0235_),
    .B2(_0224_),
    .C1(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _0635_ (.A0(\conv2.psram_ctrl.sck ),
    .A1(_0238_),
    .S(_0211_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(\conv1.psram_ctrl.sck ),
    .A1(_0239_),
    .S(_0151_),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_1 _0637_ (.A(_0240_),
    .X(net5));
 sky130_fd_sc_hd__mux2_1 _0638_ (.A0(\softmax.psram_ce_n ),
    .A1(\maxpool.psram_ce_n ),
    .S(_0229_),
    .X(_0241_));
 sky130_fd_sc_hd__inv_2 _0639_ (.A(\fc1.psram_ce_n ),
    .Y(_0242_));
 sky130_fd_sc_hd__nor2_1 _0640_ (.A(_0242_),
    .B(_0225_),
    .Y(_0243_));
 sky130_fd_sc_hd__a221o_1 _0641_ (.A1(\fc2.psram_ce_n ),
    .A2(_0234_),
    .B1(_0241_),
    .B2(_0224_),
    .C1(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(\conv2.psram_ce_n ),
    .A1(_0244_),
    .S(_0211_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _0643_ (.A0(\conv1.psram_ce_n ),
    .A1(_0245_),
    .S(_0151_),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_1 _0644_ (.A(_0246_),
    .X(net4));
 sky130_fd_sc_hd__a21o_1 _0645_ (.A1(\conv1.psram_ctrl.counter[0] ),
    .A2(\conv1.addr[8] ),
    .B1(_0171_),
    .X(_0247_));
 sky130_fd_sc_hd__o21ai_1 _0646_ (.A1(\conv1.psram_ctrl.counter[1] ),
    .A2(\conv1.psram_ctrl.counter[2] ),
    .B1(\conv1.psram_ctrl.counter[0] ),
    .Y(_0248_));
 sky130_fd_sc_hd__a32o_1 _0647_ (.A1(\conv1.psram_ctrl.counter[1] ),
    .A2(\conv1.psram_ctrl.counter[2] ),
    .A3(_0247_),
    .B1(_0248_),
    .B2(_0171_),
    .X(_0249_));
 sky130_fd_sc_hd__or4b_2 _0648_ (.A(\conv1.psram_ctrl.counter[3] ),
    .B(\conv1.psram_ctrl.counter[5] ),
    .C(_0174_),
    .D_N(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__or3b_1 _0649_ (.A(\maxpool.psram_ctrl.counter[1] ),
    .B(\maxpool.psram_ctrl.counter[0] ),
    .C_N(\maxpool.addr[11] ),
    .X(_0251_));
 sky130_fd_sc_hd__nand3_1 _0650_ (.A(\maxpool.psram_ctrl.counter[1] ),
    .B(\maxpool.psram_ctrl.counter[0] ),
    .C(\maxpool.addr[8] ),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _0651_ (.A(\maxpool.psram_ctrl.counter[2] ),
    .Y(_0253_));
 sky130_fd_sc_hd__a21o_1 _0652_ (.A1(_0251_),
    .A2(_0252_),
    .B1(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__and2b_1 _0653_ (.A_N(\maxpool.psram_ctrl.counter[1] ),
    .B(\maxpool.psram_ctrl.counter[0] ),
    .X(_0255_));
 sky130_fd_sc_hd__a21o_1 _0654_ (.A1(\maxpool.psram_ctrl.counter[1] ),
    .A2(\maxpool.psram_ctrl.counter[0] ),
    .B1(\maxpool.psram_ctrl.counter[2] ),
    .X(_0256_));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(\maxpool.psram_ctrl.counter[4] ),
    .Y(_0257_));
 sky130_fd_sc_hd__o211a_1 _0656_ (.A1(_0253_),
    .A2(_0255_),
    .B1(_0256_),
    .C1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__or4_1 _0657_ (.A(\maxpool.psram_ctrl.counter[6] ),
    .B(\maxpool.psram_ctrl.counter[7] ),
    .C(\maxpool.psram_ctrl.counter[5] ),
    .D(\maxpool.psram_ctrl.counter[3] ),
    .X(_0259_));
 sky130_fd_sc_hd__a211o_1 _0658_ (.A1(\maxpool.psram_ctrl.counter[4] ),
    .A2(_0254_),
    .B1(_0258_),
    .C1(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__xor2_1 _0659_ (.A(\softmax.psram_ctrl.counter[2] ),
    .B(\softmax.psram_ctrl.counter[1] ),
    .X(_0261_));
 sky130_fd_sc_hd__or3_1 _0660_ (.A(\softmax.psram_ctrl.counter[4] ),
    .B(\softmax.psram_ctrl.counter[7] ),
    .C(\softmax.psram_ctrl.counter[3] ),
    .X(_0262_));
 sky130_fd_sc_hd__a2111o_1 _0661_ (.A1(\softmax.psram_ctrl.counter[0] ),
    .A2(_0261_),
    .B1(_0262_),
    .C1(\softmax.psram_ctrl.counter[6] ),
    .D1(\softmax.psram_ctrl.counter[5] ),
    .X(_0263_));
 sky130_fd_sc_hd__or2b_1 _0662_ (.A(\softmax.psram_ctrl.counter[0] ),
    .B_N(\softmax.addr[11] ),
    .X(_0264_));
 sky130_fd_sc_hd__nand3_1 _0663_ (.A(\softmax.psram_ctrl.counter[1] ),
    .B(\softmax.psram_ctrl.counter[0] ),
    .C(\softmax.addr[8] ),
    .Y(_0265_));
 sky130_fd_sc_hd__or3b_1 _0664_ (.A(\softmax.psram_ctrl.counter[5] ),
    .B(\softmax.psram_ctrl.counter[6] ),
    .C_N(\softmax.psram_ctrl.counter[2] ),
    .X(_0266_));
 sky130_fd_sc_hd__a211o_1 _0665_ (.A1(_0264_),
    .A2(_0265_),
    .B1(_0266_),
    .C1(_0217_),
    .X(_0267_));
 sky130_fd_sc_hd__and3b_1 _0666_ (.A_N(_0229_),
    .B(_0263_),
    .C(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__a211o_1 _0667_ (.A1(_0229_),
    .A2(_0260_),
    .B1(_0268_),
    .C1(_0234_),
    .X(_0269_));
 sky130_fd_sc_hd__xor2_1 _0668_ (.A(\fc2.psram_ctrl.counter[1] ),
    .B(\fc2.psram_ctrl.counter[2] ),
    .X(_0270_));
 sky130_fd_sc_hd__or4_1 _0669_ (.A(\fc2.psram_ctrl.counter[3] ),
    .B(\fc2.psram_ctrl.counter[5] ),
    .C(\fc2.psram_ctrl.counter[7] ),
    .D(\fc2.psram_ctrl.counter[6] ),
    .X(_0271_));
 sky130_fd_sc_hd__a31o_1 _0670_ (.A1(\fc2.psram_ctrl.counter[0] ),
    .A2(_0153_),
    .A3(_0270_),
    .B1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _0671_ (.A(\fc2.psram_ctrl.counter[1] ),
    .B(\fc2.psram_ctrl.counter[0] ),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _0672_ (.A0(\fc2.addr[10] ),
    .A1(\fc2.addr[8] ),
    .S(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__a31o_1 _0673_ (.A1(\fc2.psram_ctrl.counter[2] ),
    .A2(_0155_),
    .A3(_0274_),
    .B1(_0153_),
    .X(_0275_));
 sky130_fd_sc_hd__or3b_1 _0674_ (.A(_0228_),
    .B(_0272_),
    .C_N(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__or2b_1 _0675_ (.A(\fc1.addr[8] ),
    .B_N(\fc1.psram_ctrl.counter[1] ),
    .X(_0277_));
 sky130_fd_sc_hd__a21boi_1 _0676_ (.A1(\fc1.psram_ctrl.counter[0] ),
    .A2(_0277_),
    .B1_N(\fc1.psram_ctrl.counter[4] ),
    .Y(_0278_));
 sky130_fd_sc_hd__a21oi_1 _0677_ (.A1(\fc1.psram_ctrl.counter[4] ),
    .A2(\fc1.addr[10] ),
    .B1(\fc1.psram_ctrl.counter[1] ),
    .Y(_0279_));
 sky130_fd_sc_hd__o21a_1 _0678_ (.A1(\fc1.psram_ctrl.counter[1] ),
    .A2(\fc1.psram_ctrl.counter[2] ),
    .B1(\fc1.psram_ctrl.counter[0] ),
    .X(_0280_));
 sky130_fd_sc_hd__o32a_1 _0679_ (.A1(_0178_),
    .A2(_0278_),
    .A3(_0279_),
    .B1(\fc1.psram_ctrl.counter[4] ),
    .B2(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__or3_1 _0680_ (.A(\fc1.psram_ctrl.counter[3] ),
    .B(\fc1.psram_ctrl.counter[5] ),
    .C(_0181_),
    .X(_0282_));
 sky130_fd_sc_hd__o21ba_1 _0681_ (.A1(_0281_),
    .A2(_0282_),
    .B1_N(_0225_),
    .X(_0283_));
 sky130_fd_sc_hd__a311o_1 _0682_ (.A1(_0225_),
    .A2(_0269_),
    .A3(_0276_),
    .B1(_0283_),
    .C1(_0169_),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _0683_ (.A(\conv2.psram_ctrl.counter[3] ),
    .B(\conv2.psram_ctrl.counter[5] ),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _0684_ (.A0(\conv2.addr[9] ),
    .A1(\conv2.addr[8] ),
    .S(\conv2.psram_ctrl.counter[0] ),
    .X(_0286_));
 sky130_fd_sc_hd__o21ai_1 _0685_ (.A1(\conv2.psram_ctrl.counter[1] ),
    .A2(\conv2.psram_ctrl.counter[2] ),
    .B1(\conv2.psram_ctrl.counter[0] ),
    .Y(_0287_));
 sky130_fd_sc_hd__a21o_1 _0686_ (.A1(\conv2.psram_ctrl.counter[1] ),
    .A2(\conv2.psram_ctrl.counter[2] ),
    .B1(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__a32o_1 _0687_ (.A1(\conv2.psram_ctrl.counter[1] ),
    .A2(\conv2.psram_ctrl.counter[2] ),
    .A3(_0286_),
    .B1(_0288_),
    .B2(_0161_),
    .X(_0289_));
 sky130_fd_sc_hd__or4b_1 _0688_ (.A(_0164_),
    .B(_0211_),
    .C(_0285_),
    .D_N(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__a21o_1 _0689_ (.A1(_0284_),
    .A2(_0290_),
    .B1(_0170_),
    .X(_0291_));
 sky130_fd_sc_hd__o21ai_4 _0690_ (.A1(_0151_),
    .A2(_0250_),
    .B1(_0291_),
    .Y(psram_d[0]));
 sky130_fd_sc_hd__mux2_1 _0691_ (.A0(net89),
    .A1(_0177_),
    .S(\conv1.psram_ctrl.state ),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _0692_ (.A(_0292_),
    .X(\conv1.psram_ctrl.nstate ));
 sky130_fd_sc_hd__mux2_1 _0693_ (.A0(net124),
    .A1(_0167_),
    .S(\conv2.psram_ctrl.state ),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _0694_ (.A(_0293_),
    .X(\conv2.psram_ctrl.nstate ));
 sky130_fd_sc_hd__mux2_1 _0695_ (.A0(net92),
    .A1(_0184_),
    .S(\fc1.psram_ctrl.state ),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _0696_ (.A(_0294_),
    .X(\fc1.psram_ctrl.nstate ));
 sky130_fd_sc_hd__mux2_1 _0697_ (.A0(net116),
    .A1(_0158_),
    .S(\fc2.psram_ctrl.state ),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _0698_ (.A(_0295_),
    .X(\fc2.psram_ctrl.nstate ));
 sky130_fd_sc_hd__nand2_1 _0699_ (.A(\maxpool.psram_ctrl.counter[5] ),
    .B(\maxpool.psram_ctrl.counter[4] ),
    .Y(_0296_));
 sky130_fd_sc_hd__or2_1 _0700_ (.A(\maxpool.psram_ctrl.counter[1] ),
    .B(\maxpool.psram_ctrl.counter[0] ),
    .X(_0297_));
 sky130_fd_sc_hd__or3_1 _0701_ (.A(\maxpool.psram_ctrl.counter[6] ),
    .B(\maxpool.psram_ctrl.counter[7] ),
    .C(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__or4_2 _0702_ (.A(\maxpool.psram_ctrl.counter[3] ),
    .B(\maxpool.psram_ctrl.counter[2] ),
    .C(_0296_),
    .D(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _0703_ (.A0(net131),
    .A1(_0299_),
    .S(\maxpool.psram_ctrl.state ),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_1 _0704_ (.A(_0300_),
    .X(\maxpool.psram_ctrl.nstate ));
 sky130_fd_sc_hd__mux2_1 _0705_ (.A0(net81),
    .A1(_0221_),
    .S(\softmax.psram_ctrl.state ),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0706_ (.A(_0301_),
    .X(\softmax.psram_ctrl.nstate ));
 sky130_fd_sc_hd__inv_2 _0707_ (.A(net87),
    .Y(_0302_));
 sky130_fd_sc_hd__nor2_1 _0708_ (.A(_0302_),
    .B(_0158_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0709_ (.A(net130),
    .Y(_0303_));
 sky130_fd_sc_hd__nor2_1 _0710_ (.A(_0303_),
    .B(_0158_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(net150),
    .Y(_0304_));
 sky130_fd_sc_hd__nor2_1 _0712_ (.A(_0304_),
    .B(_0177_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(net94),
    .Y(_0305_));
 sky130_fd_sc_hd__nor2_1 _0714_ (.A(_0305_),
    .B(_0177_),
    .Y(_0001_));
 sky130_fd_sc_hd__nand2_1 _0715_ (.A(net47),
    .B(_0177_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _0716_ (.A(net77),
    .Y(_0306_));
 sky130_fd_sc_hd__nor2_1 _0717_ (.A(_0306_),
    .B(_0184_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(net125),
    .Y(_0307_));
 sky130_fd_sc_hd__nor2_1 _0719_ (.A(_0307_),
    .B(_0184_),
    .Y(_0004_));
 sky130_fd_sc_hd__and3_1 _0720_ (.A(\mfcc.log.data_valid ),
    .B(_0198_),
    .C(net53),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _0721_ (.A(_0308_),
    .X(_0009_));
 sky130_fd_sc_hd__and3_1 _0722_ (.A(_0198_),
    .B(\mfcc.log.state[1] ),
    .C(_0196_),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _0723_ (.A(_0309_),
    .X(_0008_));
 sky130_fd_sc_hd__nand2_1 _0724_ (.A(net31),
    .B(_0167_),
    .Y(_0033_));
 sky130_fd_sc_hd__nand2_1 _0725_ (.A(net42),
    .B(_0184_),
    .Y(_0034_));
 sky130_fd_sc_hd__nand2_1 _0726_ (.A(net43),
    .B(_0158_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(net113),
    .Y(_0310_));
 sky130_fd_sc_hd__nor2_1 _0728_ (.A(_0310_),
    .B(_0167_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(net69),
    .Y(_0311_));
 sky130_fd_sc_hd__nor2_1 _0730_ (.A(_0311_),
    .B(_0167_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand2_1 _0731_ (.A(net44),
    .B(_0299_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand2_1 _0732_ (.A(net52),
    .B(_0221_),
    .Y(_0037_));
 sky130_fd_sc_hd__nor2_1 _0733_ (.A(\softmax.psram_ctrl.sck ),
    .B(\softmax.psram_ce_n ),
    .Y(_0312_));
 sky130_fd_sc_hd__and2_1 _0734_ (.A(\softmax.psram_ctrl.sck ),
    .B(\softmax.psram_ce_n ),
    .X(_0313_));
 sky130_fd_sc_hd__o21a_1 _0735_ (.A1(_0312_),
    .A2(_0313_),
    .B1(_0221_),
    .X(_0039_));
 sky130_fd_sc_hd__a21oi_1 _0736_ (.A1(\mfcc.dct.state[1] ),
    .A2(_0188_),
    .B1(net104),
    .Y(_0314_));
 sky130_fd_sc_hd__clkbuf_4 _0737_ (.A(net22),
    .X(_0315_));
 sky130_fd_sc_hd__a31o_1 _0738_ (.A1(\mfcc.dct.output_counter[0] ),
    .A2(\mfcc.dct.state[1] ),
    .A3(_0188_),
    .B1(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__nor2_1 _0739_ (.A(_0314_),
    .B(_0316_),
    .Y(_0040_));
 sky130_fd_sc_hd__a31o_1 _0740_ (.A1(\mfcc.dct.output_counter[0] ),
    .A2(\mfcc.dct.state[1] ),
    .A3(_0188_),
    .B1(\mfcc.dct.output_counter[1] ),
    .X(_0317_));
 sky130_fd_sc_hd__nor3b_1 _0741_ (.A(_0193_),
    .B(_0189_),
    .C_N(_0317_),
    .Y(_0041_));
 sky130_fd_sc_hd__nor2_1 _0742_ (.A(_0315_),
    .B(_0191_),
    .Y(_0318_));
 sky130_fd_sc_hd__o21a_1 _0743_ (.A1(net57),
    .A2(_0189_),
    .B1(_0318_),
    .X(_0042_));
 sky130_fd_sc_hd__a211o_1 _0744_ (.A1(\mfcc.dct.output_counter[3] ),
    .A2(_0191_),
    .B1(_0185_),
    .C1(_0315_),
    .X(_0319_));
 sky130_fd_sc_hd__o21ba_1 _0745_ (.A1(net110),
    .A2(_0191_),
    .B1_N(_0319_),
    .X(_0043_));
 sky130_fd_sc_hd__a21oi_1 _0746_ (.A1(\mfcc.dct.output_counter[3] ),
    .A2(_0191_),
    .B1(net50),
    .Y(_0320_));
 sky130_fd_sc_hd__and3_1 _0747_ (.A(\mfcc.dct.output_counter[4] ),
    .B(\mfcc.dct.output_counter[3] ),
    .C(_0191_),
    .X(_0321_));
 sky130_fd_sc_hd__nor3_1 _0748_ (.A(_0193_),
    .B(_0320_),
    .C(_0321_),
    .Y(_0044_));
 sky130_fd_sc_hd__a221o_1 _0749_ (.A1(_0185_),
    .A2(_0191_),
    .B1(_0321_),
    .B2(\mfcc.dct.output_counter[5] ),
    .C1(_0315_),
    .X(_0322_));
 sky130_fd_sc_hd__o21ba_1 _0750_ (.A1(net63),
    .A2(_0321_),
    .B1_N(_0322_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0751_ (.A0(\mfcc.dct.state[1] ),
    .A1(\mfcc.dct.data_valid ),
    .S(\mfcc.dct.state[0] ),
    .X(_0323_));
 sky130_fd_sc_hd__and2_1 _0752_ (.A(\mfcc.dct.input_counter[0] ),
    .B(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__nor2_1 _0753_ (.A(_0315_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__o21a_1 _0754_ (.A1(net68),
    .A2(_0323_),
    .B1(_0325_),
    .X(_0046_));
 sky130_fd_sc_hd__and3_1 _0755_ (.A(\mfcc.dct.input_counter[1] ),
    .B(\mfcc.dct.input_counter[0] ),
    .C(_0323_),
    .X(_0326_));
 sky130_fd_sc_hd__o21ai_1 _0756_ (.A1(net158),
    .A2(_0324_),
    .B1(_0038_),
    .Y(_0327_));
 sky130_fd_sc_hd__nor2_1 _0757_ (.A(_0326_),
    .B(_0327_),
    .Y(_0047_));
 sky130_fd_sc_hd__a31o_1 _0758_ (.A1(\mfcc.dct.input_counter[2] ),
    .A2(\mfcc.dct.input_counter[1] ),
    .A3(_0324_),
    .B1(_0315_),
    .X(_0328_));
 sky130_fd_sc_hd__o21ba_1 _0759_ (.A1(net119),
    .A2(_0326_),
    .B1_N(_0328_),
    .X(_0048_));
 sky130_fd_sc_hd__a31oi_1 _0760_ (.A1(net168),
    .A2(\mfcc.dct.input_counter[1] ),
    .A3(_0324_),
    .B1(net72),
    .Y(_0329_));
 sky130_fd_sc_hd__and4_1 _0761_ (.A(\mfcc.dct.input_counter[3] ),
    .B(\mfcc.dct.input_counter[2] ),
    .C(\mfcc.dct.input_counter[1] ),
    .D(_0324_),
    .X(_0330_));
 sky130_fd_sc_hd__nor3_1 _0762_ (.A(_0193_),
    .B(_0329_),
    .C(_0330_),
    .Y(_0049_));
 sky130_fd_sc_hd__o21ai_1 _0763_ (.A1(net49),
    .A2(_0330_),
    .B1(_0038_),
    .Y(_0331_));
 sky130_fd_sc_hd__a21oi_1 _0764_ (.A1(net49),
    .A2(_0330_),
    .B1(_0331_),
    .Y(_0050_));
 sky130_fd_sc_hd__a21oi_1 _0765_ (.A1(_0185_),
    .A2(_0191_),
    .B1(net30),
    .Y(_0332_));
 sky130_fd_sc_hd__nor2_1 _0766_ (.A(_0193_),
    .B(_0332_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(\mfcc.log.state[2] ),
    .Y(_0333_));
 sky130_fd_sc_hd__a21oi_1 _0768_ (.A1(\mfcc.log.state[1] ),
    .A2(_0333_),
    .B1(net82),
    .Y(_0334_));
 sky130_fd_sc_hd__and4_1 _0769_ (.A(\mfcc.log.shift_count[0] ),
    .B(\mfcc.log.state[1] ),
    .C(_0333_),
    .D(_0196_),
    .X(_0335_));
 sky130_fd_sc_hd__nor3_1 _0770_ (.A(_0193_),
    .B(_0334_),
    .C(_0335_),
    .Y(_0052_));
 sky130_fd_sc_hd__o21ai_1 _0771_ (.A1(net67),
    .A2(_0335_),
    .B1(_0038_),
    .Y(_0336_));
 sky130_fd_sc_hd__a21oi_1 _0772_ (.A1(net67),
    .A2(_0335_),
    .B1(_0336_),
    .Y(_0053_));
 sky130_fd_sc_hd__a21oi_1 _0773_ (.A1(\mfcc.log.shift_count[1] ),
    .A2(_0335_),
    .B1(net96),
    .Y(_0337_));
 sky130_fd_sc_hd__and3_1 _0774_ (.A(\mfcc.log.shift_count[2] ),
    .B(\mfcc.log.shift_count[1] ),
    .C(_0335_),
    .X(_0338_));
 sky130_fd_sc_hd__nor3_1 _0775_ (.A(_0193_),
    .B(net97),
    .C(_0338_),
    .Y(_0054_));
 sky130_fd_sc_hd__o21a_1 _0776_ (.A1(net51),
    .A2(_0338_),
    .B1(_0038_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(net161),
    .A1(\maxpool.state[1] ),
    .S(_0027_),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _0778_ (.A(_0339_),
    .X(_0056_));
 sky130_fd_sc_hd__or2_1 _0779_ (.A(net128),
    .B(_0027_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _0780_ (.A(_0340_),
    .X(_0057_));
 sky130_fd_sc_hd__nor2_1 _0781_ (.A(\mfcc.log.state[1] ),
    .B(_0333_),
    .Y(_0341_));
 sky130_fd_sc_hd__o31a_1 _0782_ (.A1(net120),
    .A2(_0197_),
    .A3(_0341_),
    .B1(_0038_),
    .X(_0058_));
 sky130_fd_sc_hd__o21a_1 _0783_ (.A1(net73),
    .A2(_0210_),
    .B1(_0038_),
    .X(_0059_));
 sky130_fd_sc_hd__or2b_1 _0784_ (.A(\mfcc.mel.state[0] ),
    .B_N(_0210_),
    .X(_0342_));
 sky130_fd_sc_hd__nor2_1 _0785_ (.A(_0207_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__and2b_1 _0786_ (.A_N(\mfcc.mel.state[0] ),
    .B(_0210_),
    .X(_0344_));
 sky130_fd_sc_hd__and2_1 _0787_ (.A(\mfcc.mel.filter_counter[0] ),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__nor2_1 _0788_ (.A(_0315_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__o21a_1 _0789_ (.A1(net115),
    .A2(_0343_),
    .B1(_0346_),
    .X(_0060_));
 sky130_fd_sc_hd__and3_1 _0790_ (.A(\mfcc.mel.filter_counter[1] ),
    .B(\mfcc.mel.filter_counter[0] ),
    .C(_0344_),
    .X(_0347_));
 sky130_fd_sc_hd__nor2_1 _0791_ (.A(_0315_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__o21a_1 _0792_ (.A1(net105),
    .A2(_0345_),
    .B1(_0348_),
    .X(_0061_));
 sky130_fd_sc_hd__o21ai_1 _0793_ (.A1(net66),
    .A2(_0347_),
    .B1(_0038_),
    .Y(_0349_));
 sky130_fd_sc_hd__a21oi_1 _0794_ (.A1(net66),
    .A2(_0347_),
    .B1(_0349_),
    .Y(_0062_));
 sky130_fd_sc_hd__and4_2 _0795_ (.A(\mfcc.mel.filter_counter[3] ),
    .B(\mfcc.mel.filter_counter[2] ),
    .C(\mfcc.mel.filter_counter[1] ),
    .D(\mfcc.mel.filter_counter[0] ),
    .X(_0350_));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__a22o_1 _0797_ (.A1(\mfcc.mel.filter_counter[3] ),
    .A2(_0342_),
    .B1(_0343_),
    .B2(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__a31o_1 _0798_ (.A1(\mfcc.mel.filter_counter[2] ),
    .A2(\mfcc.mel.filter_counter[1] ),
    .A3(\mfcc.mel.filter_counter[0] ),
    .B1(\mfcc.mel.filter_counter[3] ),
    .X(_0353_));
 sky130_fd_sc_hd__and3_1 _0799_ (.A(_0198_),
    .B(_0352_),
    .C(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _0800_ (.A(_0354_),
    .X(_0063_));
 sky130_fd_sc_hd__a21oi_1 _0801_ (.A1(_0344_),
    .A2(_0350_),
    .B1(net127),
    .Y(_0355_));
 sky130_fd_sc_hd__a31o_1 _0802_ (.A1(\mfcc.mel.filter_counter[4] ),
    .A2(_0344_),
    .A3(_0350_),
    .B1(_0315_),
    .X(_0356_));
 sky130_fd_sc_hd__nor2_1 _0803_ (.A(_0355_),
    .B(_0356_),
    .Y(_0064_));
 sky130_fd_sc_hd__a21o_1 _0804_ (.A1(\mfcc.mel.filter_counter[4] ),
    .A2(_0350_),
    .B1(\mfcc.mel.filter_counter[5] ),
    .X(_0357_));
 sky130_fd_sc_hd__nand3_1 _0805_ (.A(\mfcc.mel.filter_counter[5] ),
    .B(\mfcc.mel.filter_counter[4] ),
    .C(_0350_),
    .Y(_0358_));
 sky130_fd_sc_hd__a32o_1 _0806_ (.A1(_0343_),
    .A2(_0357_),
    .A3(_0358_),
    .B1(_0342_),
    .B2(\mfcc.mel.filter_counter[5] ),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _0807_ (.A(_0198_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _0808_ (.A(_0360_),
    .X(_0065_));
 sky130_fd_sc_hd__o21a_1 _0809_ (.A1(\mfcc.mel.coeff_counter[0] ),
    .A2(_0205_),
    .B1(\mfcc.mel.state[1] ),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _0810_ (.A(\mfcc.mel.state[1] ),
    .B(\mfcc.mel.coeff_counter[0] ),
    .X(_0362_));
 sky130_fd_sc_hd__and3b_1 _0811_ (.A_N(_0361_),
    .B(_0362_),
    .C(_0198_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _0812_ (.A(_0363_),
    .X(_0066_));
 sky130_fd_sc_hd__xnor2_1 _0813_ (.A(net145),
    .B(_0361_),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _0814_ (.A(_0193_),
    .B(_0364_),
    .Y(_0067_));
 sky130_fd_sc_hd__and4_1 _0815_ (.A(\mfcc.mel.state[1] ),
    .B(\mfcc.mel.coeff_counter[2] ),
    .C(\mfcc.mel.coeff_counter[1] ),
    .D(\mfcc.mel.coeff_counter[0] ),
    .X(_0365_));
 sky130_fd_sc_hd__a31o_1 _0816_ (.A1(\mfcc.mel.state[1] ),
    .A2(\mfcc.mel.coeff_counter[1] ),
    .A3(\mfcc.mel.coeff_counter[0] ),
    .B1(\mfcc.mel.coeff_counter[2] ),
    .X(_0366_));
 sky130_fd_sc_hd__or4b_1 _0817_ (.A(net12),
    .B(_0210_),
    .C(_0365_),
    .D_N(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__inv_2 _0818_ (.A(_0367_),
    .Y(_0068_));
 sky130_fd_sc_hd__and2_1 _0819_ (.A(\mfcc.mel.coeff_counter[3] ),
    .B(_0365_),
    .X(_0368_));
 sky130_fd_sc_hd__o21ai_1 _0820_ (.A1(net76),
    .A2(_0365_),
    .B1(_0038_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _0821_ (.A(_0368_),
    .B(_0369_),
    .Y(_0069_));
 sky130_fd_sc_hd__a211o_1 _0822_ (.A1(\mfcc.mel.coeff_counter[4] ),
    .A2(_0368_),
    .B1(_0210_),
    .C1(_0315_),
    .X(_0370_));
 sky130_fd_sc_hd__o21ba_1 _0823_ (.A1(net59),
    .A2(_0368_),
    .B1_N(_0370_),
    .X(_0070_));
 sky130_fd_sc_hd__or2_1 _0824_ (.A(\maxpool.psram_ctrl.sck ),
    .B(\maxpool.psram_ce_n ),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_1 _0825_ (.A(\maxpool.psram_ctrl.sck ),
    .B(net136),
    .Y(_0372_));
 sky130_fd_sc_hd__nor4_1 _0826_ (.A(\maxpool.psram_ctrl.counter[3] ),
    .B(\maxpool.psram_ctrl.counter[2] ),
    .C(_0296_),
    .D(_0298_),
    .Y(_0373_));
 sky130_fd_sc_hd__a21oi_1 _0827_ (.A1(_0371_),
    .A2(_0372_),
    .B1(net6),
    .Y(_0071_));
 sky130_fd_sc_hd__o21a_1 _0828_ (.A1(net90),
    .A2(_0031_),
    .B1(_0304_),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _0829_ (.A(\conv1.psram_ctrl.sck ),
    .B(_0177_),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _0830_ (.A(\conv1.psram_ctrl.sck ),
    .B(_0176_),
    .Y(_0375_));
 sky130_fd_sc_hd__and2_1 _0831_ (.A(\conv1.psram_ctrl.state ),
    .B(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _0832_ (.A0(_0374_),
    .A1(_0376_),
    .S(\conv1.psram_ctrl.counter[0] ),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _0833_ (.A(_0377_),
    .X(_0073_));
 sky130_fd_sc_hd__nand2_1 _0834_ (.A(\conv1.psram_ctrl.counter[1] ),
    .B(\conv1.psram_ctrl.counter[0] ),
    .Y(_0378_));
 sky130_fd_sc_hd__a32o_1 _0835_ (.A1(\conv1.psram_ctrl.sck ),
    .A2(_0173_),
    .A3(_0378_),
    .B1(_0376_),
    .B2(net134),
    .X(_0074_));
 sky130_fd_sc_hd__a21o_1 _0836_ (.A1(\conv1.psram_ctrl.counter[1] ),
    .A2(\conv1.psram_ctrl.counter[0] ),
    .B1(\conv1.psram_ctrl.counter[2] ),
    .X(_0379_));
 sky130_fd_sc_hd__and3_1 _0837_ (.A(\conv1.psram_ctrl.counter[1] ),
    .B(\conv1.psram_ctrl.counter[0] ),
    .C(\conv1.psram_ctrl.counter[2] ),
    .X(_0380_));
 sky130_fd_sc_hd__inv_2 _0838_ (.A(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__a32o_1 _0839_ (.A1(_0374_),
    .A2(_0379_),
    .A3(_0381_),
    .B1(_0376_),
    .B2(net157),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _0840_ (.A(\conv1.psram_ctrl.counter[3] ),
    .B(_0380_),
    .X(_0382_));
 sky130_fd_sc_hd__o21ai_1 _0841_ (.A1(\conv1.psram_ctrl.counter[3] ),
    .A2(_0380_),
    .B1(_0374_),
    .Y(_0383_));
 sky130_fd_sc_hd__a2bb2o_1 _0842_ (.A1_N(_0382_),
    .A2_N(_0383_),
    .B1(\conv1.psram_ctrl.counter[3] ),
    .B2(_0376_),
    .X(_0076_));
 sky130_fd_sc_hd__and3_1 _0843_ (.A(\conv1.psram_ctrl.counter[3] ),
    .B(\conv1.psram_ctrl.counter[4] ),
    .C(_0380_),
    .X(_0384_));
 sky130_fd_sc_hd__o21bai_1 _0844_ (.A1(_0375_),
    .A2(_0384_),
    .B1_N(_0376_),
    .Y(_0385_));
 sky130_fd_sc_hd__and3_1 _0845_ (.A(_0171_),
    .B(\conv1.psram_ctrl.sck ),
    .C(_0382_),
    .X(_0386_));
 sky130_fd_sc_hd__a21o_1 _0846_ (.A1(net93),
    .A2(_0385_),
    .B1(_0386_),
    .X(_0077_));
 sky130_fd_sc_hd__and3_1 _0847_ (.A(\conv1.psram_ctrl.sck ),
    .B(_0177_),
    .C(_0384_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(_0387_),
    .A1(_0385_),
    .S(\conv1.psram_ctrl.counter[5] ),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _0849_ (.A(_0388_),
    .X(_0078_));
 sky130_fd_sc_hd__and3_1 _0850_ (.A(\conv1.psram_ctrl.counter[5] ),
    .B(\conv1.psram_ctrl.counter[6] ),
    .C(_0384_),
    .X(_0389_));
 sky130_fd_sc_hd__nor2_1 _0851_ (.A(_0375_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__or2_1 _0852_ (.A(_0376_),
    .B(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__a32o_1 _0853_ (.A1(\conv1.psram_ctrl.counter[5] ),
    .A2(_0384_),
    .A3(_0390_),
    .B1(_0391_),
    .B2(net60),
    .X(_0079_));
 sky130_fd_sc_hd__nor2_1 _0854_ (.A(net95),
    .B(_0375_),
    .Y(_0392_));
 sky130_fd_sc_hd__a22o_1 _0855_ (.A1(net95),
    .A2(_0391_),
    .B1(_0392_),
    .B2(_0389_),
    .X(_0080_));
 sky130_fd_sc_hd__o31a_1 _0856_ (.A1(\conv2.psram_ctrl.has_wait_states ),
    .A2(net74),
    .A3(\conv2.state[2] ),
    .B1(_0311_),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _0857_ (.A(\conv2.psram_ctrl.sck ),
    .B(_0167_),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_1 _0858_ (.A(\conv2.psram_ctrl.sck ),
    .B(_0166_),
    .Y(_0394_));
 sky130_fd_sc_hd__and2_2 _0859_ (.A(\conv2.psram_ctrl.state ),
    .B(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _0860_ (.A0(_0393_),
    .A1(_0395_),
    .S(\conv2.psram_ctrl.counter[0] ),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _0861_ (.A(_0396_),
    .X(_0082_));
 sky130_fd_sc_hd__nand2_1 _0862_ (.A(\conv2.psram_ctrl.counter[1] ),
    .B(\conv2.psram_ctrl.counter[0] ),
    .Y(_0397_));
 sky130_fd_sc_hd__a32o_1 _0863_ (.A1(net154),
    .A2(_0163_),
    .A3(_0397_),
    .B1(_0395_),
    .B2(\conv2.psram_ctrl.counter[1] ),
    .X(_0083_));
 sky130_fd_sc_hd__a21o_1 _0864_ (.A1(\conv2.psram_ctrl.counter[1] ),
    .A2(\conv2.psram_ctrl.counter[0] ),
    .B1(\conv2.psram_ctrl.counter[2] ),
    .X(_0398_));
 sky130_fd_sc_hd__nand3_1 _0865_ (.A(\conv2.psram_ctrl.counter[1] ),
    .B(\conv2.psram_ctrl.counter[0] ),
    .C(\conv2.psram_ctrl.counter[2] ),
    .Y(_0399_));
 sky130_fd_sc_hd__a32o_1 _0866_ (.A1(_0393_),
    .A2(_0398_),
    .A3(_0399_),
    .B1(_0395_),
    .B2(\conv2.psram_ctrl.counter[2] ),
    .X(_0084_));
 sky130_fd_sc_hd__a31o_1 _0867_ (.A1(\conv2.psram_ctrl.counter[1] ),
    .A2(\conv2.psram_ctrl.counter[0] ),
    .A3(\conv2.psram_ctrl.counter[2] ),
    .B1(\conv2.psram_ctrl.counter[3] ),
    .X(_0400_));
 sky130_fd_sc_hd__and4_1 _0868_ (.A(\conv2.psram_ctrl.counter[1] ),
    .B(\conv2.psram_ctrl.counter[0] ),
    .C(\conv2.psram_ctrl.counter[3] ),
    .D(\conv2.psram_ctrl.counter[2] ),
    .X(_0401_));
 sky130_fd_sc_hd__inv_2 _0869_ (.A(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__a32o_1 _0870_ (.A1(_0393_),
    .A2(_0400_),
    .A3(_0402_),
    .B1(_0395_),
    .B2(net151),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _0871_ (.A(\conv2.psram_ctrl.counter[4] ),
    .B(_0401_),
    .X(_0403_));
 sky130_fd_sc_hd__nor2_1 _0872_ (.A(_0394_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__or2_1 _0873_ (.A(_0395_),
    .B(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _0874_ (.A1(_0401_),
    .A2(_0404_),
    .B1(_0405_),
    .B2(net103),
    .X(_0086_));
 sky130_fd_sc_hd__and3_1 _0875_ (.A(\conv2.psram_ctrl.sck ),
    .B(_0167_),
    .C(_0403_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _0876_ (.A0(_0406_),
    .A1(_0405_),
    .S(\conv2.psram_ctrl.counter[5] ),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _0877_ (.A(_0407_),
    .X(_0087_));
 sky130_fd_sc_hd__and3_1 _0878_ (.A(\conv2.psram_ctrl.counter[5] ),
    .B(\conv2.psram_ctrl.counter[6] ),
    .C(_0403_),
    .X(_0408_));
 sky130_fd_sc_hd__nor2_1 _0879_ (.A(_0394_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__or2_1 _0880_ (.A(_0395_),
    .B(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__a32o_1 _0881_ (.A1(\conv2.psram_ctrl.counter[5] ),
    .A2(_0403_),
    .A3(_0409_),
    .B1(_0410_),
    .B2(net64),
    .X(_0088_));
 sky130_fd_sc_hd__nor2_1 _0882_ (.A(net83),
    .B(_0394_),
    .Y(_0411_));
 sky130_fd_sc_hd__a22o_1 _0883_ (.A1(net83),
    .A2(_0410_),
    .B1(_0411_),
    .B2(_0408_),
    .X(_0089_));
 sky130_fd_sc_hd__inv_2 _0884_ (.A(\conv1.state[3] ),
    .Y(_0412_));
 sky130_fd_sc_hd__a31o_1 _0885_ (.A1(_0412_),
    .A2(_0304_),
    .A3(net84),
    .B1(\conv1.state[2] ),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_1 _0886_ (.A(\conv1.psram_ce_n ),
    .B(\conv1.psram_ctrl.sck ),
    .Y(_0413_));
 sky130_fd_sc_hd__and2_1 _0887_ (.A(\conv1.psram_ce_n ),
    .B(\conv1.psram_ctrl.sck ),
    .X(_0414_));
 sky130_fd_sc_hd__o21a_1 _0888_ (.A1(_0413_),
    .A2(_0414_),
    .B1(_0177_),
    .X(_0091_));
 sky130_fd_sc_hd__o31a_1 _0889_ (.A1(\fc1.psram_ctrl.has_wait_states ),
    .A2(net77),
    .A3(net106),
    .B1(_0307_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _0890_ (.A(\fc1.psram_ctrl.sck ),
    .B(_0184_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_1 _0891_ (.A(\fc1.psram_ctrl.sck ),
    .B(_0184_),
    .Y(_0416_));
 sky130_fd_sc_hd__and2_2 _0892_ (.A(\fc1.psram_ctrl.state ),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _0893_ (.A0(_0415_),
    .A1(_0417_),
    .S(\fc1.psram_ctrl.counter[0] ),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _0894_ (.A(_0418_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _0895_ (.A(\fc1.psram_ctrl.counter[1] ),
    .B(\fc1.psram_ctrl.counter[0] ),
    .Y(_0419_));
 sky130_fd_sc_hd__a32o_1 _0896_ (.A1(net117),
    .A2(_0182_),
    .A3(_0419_),
    .B1(_0417_),
    .B2(\fc1.psram_ctrl.counter[1] ),
    .X(_0094_));
 sky130_fd_sc_hd__nand2_1 _0897_ (.A(_0178_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__or2_1 _0898_ (.A(_0178_),
    .B(_0419_),
    .X(_0421_));
 sky130_fd_sc_hd__a32o_1 _0899_ (.A1(_0415_),
    .A2(_0420_),
    .A3(_0421_),
    .B1(_0417_),
    .B2(net156),
    .X(_0095_));
 sky130_fd_sc_hd__a31o_1 _0900_ (.A1(\fc1.psram_ctrl.counter[1] ),
    .A2(\fc1.psram_ctrl.counter[0] ),
    .A3(\fc1.psram_ctrl.counter[2] ),
    .B1(\fc1.psram_ctrl.counter[3] ),
    .X(_0422_));
 sky130_fd_sc_hd__and4_1 _0901_ (.A(\fc1.psram_ctrl.counter[1] ),
    .B(\fc1.psram_ctrl.counter[0] ),
    .C(\fc1.psram_ctrl.counter[3] ),
    .D(\fc1.psram_ctrl.counter[2] ),
    .X(_0423_));
 sky130_fd_sc_hd__inv_2 _0902_ (.A(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__a32o_1 _0903_ (.A1(_0415_),
    .A2(_0422_),
    .A3(_0424_),
    .B1(_0417_),
    .B2(net159),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _0904_ (.A(\fc1.psram_ctrl.counter[4] ),
    .B(_0423_),
    .X(_0425_));
 sky130_fd_sc_hd__inv_2 _0905_ (.A(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21o_1 _0906_ (.A1(_0415_),
    .A2(_0426_),
    .B1(_0417_),
    .X(_0427_));
 sky130_fd_sc_hd__and3_1 _0907_ (.A(_0415_),
    .B(_0423_),
    .C(_0426_),
    .X(_0428_));
 sky130_fd_sc_hd__a21o_1 _0908_ (.A1(net163),
    .A2(_0427_),
    .B1(_0428_),
    .X(_0097_));
 sky130_fd_sc_hd__nor2_1 _0909_ (.A(_0416_),
    .B(_0426_),
    .Y(_0429_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(_0429_),
    .A1(_0427_),
    .S(\fc1.psram_ctrl.counter[5] ),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _0911_ (.A(_0430_),
    .X(_0098_));
 sky130_fd_sc_hd__and3_1 _0912_ (.A(\fc1.psram_ctrl.counter[5] ),
    .B(\fc1.psram_ctrl.counter[6] ),
    .C(_0425_),
    .X(_0431_));
 sky130_fd_sc_hd__nor2_1 _0913_ (.A(_0416_),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__or2_1 _0914_ (.A(_0417_),
    .B(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__a32o_1 _0915_ (.A1(\fc1.psram_ctrl.counter[5] ),
    .A2(_0425_),
    .A3(_0432_),
    .B1(_0433_),
    .B2(net62),
    .X(_0099_));
 sky130_fd_sc_hd__nor2_1 _0916_ (.A(net86),
    .B(_0416_),
    .Y(_0434_));
 sky130_fd_sc_hd__a22o_1 _0917_ (.A1(net86),
    .A2(_0433_),
    .B1(_0434_),
    .B2(_0431_),
    .X(_0100_));
 sky130_fd_sc_hd__inv_2 _0918_ (.A(\conv2.addr[8] ),
    .Y(_0435_));
 sky130_fd_sc_hd__o21ai_1 _0919_ (.A1(_0435_),
    .A2(_0030_),
    .B1(_0310_),
    .Y(_0101_));
 sky130_fd_sc_hd__or2_1 _0920_ (.A(net122),
    .B(_0030_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _0921_ (.A(_0436_),
    .X(_0102_));
 sky130_fd_sc_hd__nor2_1 _0922_ (.A(\conv2.psram_ce_n ),
    .B(\conv2.psram_ctrl.sck ),
    .Y(_0437_));
 sky130_fd_sc_hd__and2_1 _0923_ (.A(\conv2.psram_ce_n ),
    .B(\conv2.psram_ctrl.sck ),
    .X(_0438_));
 sky130_fd_sc_hd__o21a_1 _0924_ (.A1(_0437_),
    .A2(_0438_),
    .B1(_0167_),
    .X(_0103_));
 sky130_fd_sc_hd__nor2_1 _0925_ (.A(_0227_),
    .B(_0233_),
    .Y(_0439_));
 sky130_fd_sc_hd__and2_1 _0926_ (.A(_0227_),
    .B(_0233_),
    .X(_0440_));
 sky130_fd_sc_hd__nor2_1 _0927_ (.A(_0439_),
    .B(_0440_),
    .Y(_0104_));
 sky130_fd_sc_hd__xor2_1 _0928_ (.A(net142),
    .B(_0439_),
    .X(_0105_));
 sky130_fd_sc_hd__a21oi_1 _0929_ (.A1(\state[1] ),
    .A2(_0439_),
    .B1(net155),
    .Y(_0441_));
 sky130_fd_sc_hd__nor2_1 _0930_ (.A(net3),
    .B(_0441_),
    .Y(_0106_));
 sky130_fd_sc_hd__o21a_1 _0931_ (.A1(net132),
    .A2(_0028_),
    .B1(_0303_),
    .X(_0107_));
 sky130_fd_sc_hd__and2_1 _0932_ (.A(\fc2.psram_ctrl.sck ),
    .B(_0158_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_2 _0933_ (.A(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _0934_ (.A(\fc2.psram_ctrl.sck ),
    .B(_0158_),
    .Y(_0444_));
 sky130_fd_sc_hd__and2_2 _0935_ (.A(\fc2.psram_ctrl.state ),
    .B(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(_0443_),
    .A1(_0445_),
    .S(\fc2.psram_ctrl.counter[0] ),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0937_ (.A(_0446_),
    .X(_0108_));
 sky130_fd_sc_hd__nor2_1 _0938_ (.A(_0273_),
    .B(_0444_),
    .Y(_0447_));
 sky130_fd_sc_hd__a22o_1 _0939_ (.A1(net144),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0155_),
    .X(_0109_));
 sky130_fd_sc_hd__or2_1 _0940_ (.A(\fc2.psram_ctrl.counter[2] ),
    .B(_0273_),
    .X(_0448_));
 sky130_fd_sc_hd__nand2_1 _0941_ (.A(\fc2.psram_ctrl.counter[2] ),
    .B(_0273_),
    .Y(_0449_));
 sky130_fd_sc_hd__a32o_1 _0942_ (.A1(_0443_),
    .A2(_0448_),
    .A3(_0449_),
    .B1(_0445_),
    .B2(net133),
    .X(_0110_));
 sky130_fd_sc_hd__nand2_1 _0943_ (.A(_0156_),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__nor2_1 _0944_ (.A(_0156_),
    .B(_0449_),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _0945_ (.A(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__a32o_1 _0946_ (.A1(_0443_),
    .A2(_0450_),
    .A3(_0452_),
    .B1(_0445_),
    .B2(net149),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_1 _0947_ (.A(\fc2.psram_ctrl.counter[4] ),
    .B(_0451_),
    .Y(_0453_));
 sky130_fd_sc_hd__a21o_1 _0948_ (.A1(_0443_),
    .A2(_0453_),
    .B1(_0445_),
    .X(_0454_));
 sky130_fd_sc_hd__nor2_1 _0949_ (.A(\fc2.psram_ctrl.counter[4] ),
    .B(_0452_),
    .Y(_0455_));
 sky130_fd_sc_hd__a22o_1 _0950_ (.A1(net165),
    .A2(_0454_),
    .B1(_0455_),
    .B2(_0443_),
    .X(_0112_));
 sky130_fd_sc_hd__nor2_1 _0951_ (.A(\fc2.psram_ctrl.counter[5] ),
    .B(_0453_),
    .Y(_0456_));
 sky130_fd_sc_hd__a22o_1 _0952_ (.A1(net162),
    .A2(_0454_),
    .B1(_0456_),
    .B2(_0443_),
    .X(_0113_));
 sky130_fd_sc_hd__and4_1 _0953_ (.A(\fc2.psram_ctrl.counter[5] ),
    .B(\fc2.psram_ctrl.counter[4] ),
    .C(\fc2.psram_ctrl.counter[6] ),
    .D(_0451_),
    .X(_0457_));
 sky130_fd_sc_hd__o21bai_1 _0954_ (.A1(_0444_),
    .A2(_0457_),
    .B1_N(_0445_),
    .Y(_0458_));
 sky130_fd_sc_hd__or4b_1 _0955_ (.A(\fc2.psram_ctrl.counter[6] ),
    .B(_0444_),
    .C(_0453_),
    .D_N(\fc2.psram_ctrl.counter[5] ),
    .X(_0459_));
 sky130_fd_sc_hd__a21bo_1 _0956_ (.A1(net109),
    .A2(_0458_),
    .B1_N(_0459_),
    .X(_0114_));
 sky130_fd_sc_hd__and2_1 _0957_ (.A(_0443_),
    .B(_0457_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(_0460_),
    .A1(_0458_),
    .S(\fc2.psram_ctrl.counter[7] ),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0959_ (.A(_0461_),
    .X(_0115_));
 sky130_fd_sc_hd__inv_2 _0960_ (.A(\fc1.addr[8] ),
    .Y(_0462_));
 sky130_fd_sc_hd__o21ai_1 _0961_ (.A1(_0462_),
    .A2(_0029_),
    .B1(_0306_),
    .Y(_0116_));
 sky130_fd_sc_hd__or2_1 _0962_ (.A(net143),
    .B(_0029_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _0963_ (.A(_0463_),
    .X(_0117_));
 sky130_fd_sc_hd__nor2_1 _0964_ (.A(\fc1.psram_ctrl.sck ),
    .B(\fc1.psram_ce_n ),
    .Y(_0464_));
 sky130_fd_sc_hd__nor2_1 _0965_ (.A(_0236_),
    .B(_0242_),
    .Y(_0465_));
 sky130_fd_sc_hd__o21a_1 _0966_ (.A1(_0464_),
    .A2(_0465_),
    .B1(_0184_),
    .X(_0118_));
 sky130_fd_sc_hd__nand2_1 _0967_ (.A(\maxpool.state[0] ),
    .B(net6),
    .Y(_0466_));
 sky130_fd_sc_hd__o311a_1 _0968_ (.A1(\maxpool.state[0] ),
    .A2(net138),
    .A3(_0229_),
    .B1(_0466_),
    .C1(_0213_),
    .X(_0119_));
 sky130_fd_sc_hd__and3_1 _0969_ (.A(\maxpool.state[0] ),
    .B(\maxpool.state[1] ),
    .C(net6),
    .X(_0467_));
 sky130_fd_sc_hd__a21oi_1 _0970_ (.A1(\maxpool.state[0] ),
    .A2(net6),
    .B1(\maxpool.state[1] ),
    .Y(_0468_));
 sky130_fd_sc_hd__nor3_1 _0971_ (.A(net58),
    .B(_0467_),
    .C(_0468_),
    .Y(_0120_));
 sky130_fd_sc_hd__and2_1 _0972_ (.A(_0213_),
    .B(_0467_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _0973_ (.A(_0469_),
    .X(_0121_));
 sky130_fd_sc_hd__and2_2 _0974_ (.A(\maxpool.psram_ctrl.sck ),
    .B(_0299_),
    .X(_0470_));
 sky130_fd_sc_hd__nor2b_2 _0975_ (.A(_0470_),
    .B_N(\maxpool.psram_ctrl.state ),
    .Y(_0471_));
 sky130_fd_sc_hd__mux2_1 _0976_ (.A0(_0470_),
    .A1(_0471_),
    .S(\maxpool.psram_ctrl.counter[0] ),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0472_),
    .X(_0122_));
 sky130_fd_sc_hd__nand2_1 _0978_ (.A(\maxpool.psram_ctrl.counter[1] ),
    .B(\maxpool.psram_ctrl.counter[0] ),
    .Y(_0473_));
 sky130_fd_sc_hd__a32o_1 _0979_ (.A1(net101),
    .A2(_0297_),
    .A3(_0473_),
    .B1(_0471_),
    .B2(\maxpool.psram_ctrl.counter[1] ),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _0980_ (.A(_0253_),
    .B(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__a32o_1 _0981_ (.A1(_0256_),
    .A2(_0470_),
    .A3(_0474_),
    .B1(_0471_),
    .B2(net153),
    .X(_0124_));
 sky130_fd_sc_hd__a31o_1 _0982_ (.A1(\maxpool.psram_ctrl.counter[2] ),
    .A2(\maxpool.psram_ctrl.counter[1] ),
    .A3(\maxpool.psram_ctrl.counter[0] ),
    .B1(\maxpool.psram_ctrl.counter[3] ),
    .X(_0475_));
 sky130_fd_sc_hd__and4_1 _0983_ (.A(\maxpool.psram_ctrl.counter[3] ),
    .B(\maxpool.psram_ctrl.counter[2] ),
    .C(\maxpool.psram_ctrl.counter[1] ),
    .D(\maxpool.psram_ctrl.counter[0] ),
    .X(_0476_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__a32o_1 _0985_ (.A1(_0470_),
    .A2(_0475_),
    .A3(_0477_),
    .B1(_0471_),
    .B2(net152),
    .X(_0125_));
 sky130_fd_sc_hd__nor2_1 _0986_ (.A(_0257_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_2 _0987_ (.A(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__a21o_1 _0988_ (.A1(_0470_),
    .A2(_0479_),
    .B1(_0471_),
    .X(_0480_));
 sky130_fd_sc_hd__and3_1 _0989_ (.A(_0257_),
    .B(\maxpool.psram_ctrl.sck ),
    .C(_0476_),
    .X(_0481_));
 sky130_fd_sc_hd__a21o_1 _0990_ (.A1(net123),
    .A2(_0480_),
    .B1(_0481_),
    .X(_0126_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(\maxpool.psram_ctrl.counter[5] ),
    .Y(_0482_));
 sky130_fd_sc_hd__a31o_1 _0992_ (.A1(\maxpool.psram_ctrl.sck ),
    .A2(_0299_),
    .A3(_0478_),
    .B1(\maxpool.psram_ctrl.counter[5] ),
    .X(_0483_));
 sky130_fd_sc_hd__o21a_1 _0993_ (.A1(_0482_),
    .A2(_0480_),
    .B1(_0483_),
    .X(_0127_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(\maxpool.psram_ctrl.counter[6] ),
    .Y(_0484_));
 sky130_fd_sc_hd__o31a_1 _0995_ (.A1(_0484_),
    .A2(_0482_),
    .A3(_0479_),
    .B1(_0470_),
    .X(_0485_));
 sky130_fd_sc_hd__or2_1 _0996_ (.A(_0471_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__a32o_1 _0997_ (.A1(\maxpool.psram_ctrl.counter[5] ),
    .A2(_0478_),
    .A3(_0485_),
    .B1(_0486_),
    .B2(net139),
    .X(_0128_));
 sky130_fd_sc_hd__and4_1 _0998_ (.A(\maxpool.psram_ctrl.counter[6] ),
    .B(\maxpool.psram_ctrl.counter[5] ),
    .C(_0470_),
    .D(_0478_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(_0487_),
    .A1(_0486_),
    .S(\maxpool.psram_ctrl.counter[7] ),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(_0488_),
    .X(_0129_));
 sky130_fd_sc_hd__inv_2 _1001_ (.A(\fc2.addr[8] ),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_1 _1002_ (.A1(_0489_),
    .A2(_0028_),
    .B1(_0302_),
    .Y(_0130_));
 sky130_fd_sc_hd__or2_1 _1003_ (.A(net126),
    .B(_0028_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _1004_ (.A(_0490_),
    .X(_0131_));
 sky130_fd_sc_hd__nor2_1 _1005_ (.A(\fc2.psram_ce_n ),
    .B(\fc2.psram_ctrl.sck ),
    .Y(_0491_));
 sky130_fd_sc_hd__and2_1 _1006_ (.A(\fc2.psram_ce_n ),
    .B(\fc2.psram_ctrl.sck ),
    .X(_0492_));
 sky130_fd_sc_hd__o21a_1 _1007_ (.A1(_0491_),
    .A2(_0492_),
    .B1(_0158_),
    .X(_0132_));
 sky130_fd_sc_hd__or2_1 _1008_ (.A(\softmax.psram_ctrl.start ),
    .B(_0216_),
    .X(_0493_));
 sky130_fd_sc_hd__a21o_1 _1009_ (.A1(\softmax.addr[8] ),
    .A2(_0493_),
    .B1(net32),
    .X(_0133_));
 sky130_fd_sc_hd__or2b_1 _1010_ (.A(net167),
    .B_N(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__or2_1 _1011_ (.A(net135),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _1012_ (.A(_0495_),
    .X(_0134_));
 sky130_fd_sc_hd__and2_1 _1013_ (.A(\softmax.psram_ctrl.sck ),
    .B(_0221_),
    .X(_0496_));
 sky130_fd_sc_hd__nand2_1 _1014_ (.A(\softmax.psram_ctrl.sck ),
    .B(_0221_),
    .Y(_0497_));
 sky130_fd_sc_hd__and2_1 _1015_ (.A(\softmax.psram_ctrl.state ),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(_0496_),
    .A1(_0498_),
    .S(\softmax.psram_ctrl.counter[0] ),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _1017_ (.A(_0499_),
    .X(_0135_));
 sky130_fd_sc_hd__nand2_1 _1018_ (.A(\softmax.psram_ctrl.counter[1] ),
    .B(\softmax.psram_ctrl.counter[0] ),
    .Y(_0500_));
 sky130_fd_sc_hd__a32o_1 _1019_ (.A1(net146),
    .A2(_0218_),
    .A3(_0500_),
    .B1(_0498_),
    .B2(\softmax.psram_ctrl.counter[1] ),
    .X(_0136_));
 sky130_fd_sc_hd__a21o_1 _1020_ (.A1(\softmax.psram_ctrl.counter[1] ),
    .A2(\softmax.psram_ctrl.counter[0] ),
    .B1(\softmax.psram_ctrl.counter[2] ),
    .X(_0501_));
 sky130_fd_sc_hd__nand3_1 _1021_ (.A(\softmax.psram_ctrl.counter[2] ),
    .B(\softmax.psram_ctrl.counter[1] ),
    .C(\softmax.psram_ctrl.counter[0] ),
    .Y(_0502_));
 sky130_fd_sc_hd__a32o_1 _1022_ (.A1(_0501_),
    .A2(_0496_),
    .A3(_0502_),
    .B1(_0498_),
    .B2(net160),
    .X(_0137_));
 sky130_fd_sc_hd__a31o_1 _1023_ (.A1(\softmax.psram_ctrl.counter[2] ),
    .A2(\softmax.psram_ctrl.counter[1] ),
    .A3(\softmax.psram_ctrl.counter[0] ),
    .B1(\softmax.psram_ctrl.counter[3] ),
    .X(_0503_));
 sky130_fd_sc_hd__and4_1 _1024_ (.A(\softmax.psram_ctrl.counter[3] ),
    .B(\softmax.psram_ctrl.counter[2] ),
    .C(\softmax.psram_ctrl.counter[1] ),
    .D(\softmax.psram_ctrl.counter[0] ),
    .X(_0504_));
 sky130_fd_sc_hd__inv_2 _1025_ (.A(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__a32o_1 _1026_ (.A1(_0496_),
    .A2(_0503_),
    .A3(_0505_),
    .B1(_0498_),
    .B2(net137),
    .X(_0138_));
 sky130_fd_sc_hd__and2_1 _1027_ (.A(\softmax.psram_ctrl.counter[4] ),
    .B(_0504_),
    .X(_0506_));
 sky130_fd_sc_hd__nor2_1 _1028_ (.A(_0497_),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__or2_1 _1029_ (.A(_0498_),
    .B(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__a22o_1 _1030_ (.A1(_0504_),
    .A2(_0507_),
    .B1(_0508_),
    .B2(net100),
    .X(_0139_));
 sky130_fd_sc_hd__and3_1 _1031_ (.A(\softmax.psram_ctrl.sck ),
    .B(_0221_),
    .C(_0506_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _1032_ (.A0(_0509_),
    .A1(_0508_),
    .S(\softmax.psram_ctrl.counter[5] ),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_1 _1033_ (.A(_0510_),
    .X(_0140_));
 sky130_fd_sc_hd__nand2_1 _1034_ (.A(\softmax.psram_ctrl.state ),
    .B(_0497_),
    .Y(_0511_));
 sky130_fd_sc_hd__a31o_1 _1035_ (.A1(\softmax.psram_ctrl.counter[5] ),
    .A2(\softmax.psram_ctrl.counter[6] ),
    .A3(_0506_),
    .B1(_0497_),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_1 _1036_ (.A(_0511_),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__and3b_1 _1037_ (.A_N(\softmax.psram_ctrl.counter[6] ),
    .B(_0509_),
    .C(\softmax.psram_ctrl.counter[5] ),
    .X(_0514_));
 sky130_fd_sc_hd__a21o_1 _1038_ (.A1(net141),
    .A2(_0513_),
    .B1(_0514_),
    .X(_0141_));
 sky130_fd_sc_hd__and4_1 _1039_ (.A(\softmax.psram_ctrl.counter[5] ),
    .B(\softmax.psram_ctrl.counter[6] ),
    .C(\softmax.psram_ctrl.sck ),
    .D(_0506_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _1040_ (.A0(_0515_),
    .A1(_0513_),
    .S(\softmax.psram_ctrl.counter[7] ),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _1041_ (.A(_0516_),
    .X(_0142_));
 sky130_fd_sc_hd__a21o_1 _1042_ (.A1(net81),
    .A2(_0221_),
    .B1(_0494_),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_1 _1043_ (.A(_0221_),
    .B(_0494_),
    .Y(_0144_));
 sky130_fd_sc_hd__mux2_1 _1044_ (.A0(net106),
    .A1(net164),
    .S(_0184_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _1045_ (.A(_0517_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _1046_ (.A0(net70),
    .A1(\fc2.state[2] ),
    .S(_0158_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _1047_ (.A(_0518_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _1048_ (.A0(net166),
    .A1(\conv2.state[2] ),
    .S(_0167_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_1 _1049_ (.A(_0519_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\conv1.state[3] ),
    .A1(\conv1.state[2] ),
    .S(_0177_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(_0520_),
    .X(_0148_));
 sky130_fd_sc_hd__dfrtp_4 _1052_ (.CLK(clknet_4_11_0_clk),
    .D(_0039_),
    .RESET_B(net16),
    .Q(\softmax.psram_ctrl.sck ));
 sky130_fd_sc_hd__dfstp_1 _1053_ (.CLK(clknet_4_3_0_clk),
    .D(net56),
    .SET_B(net10),
    .Q(\conv1.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1054_ (.CLK(clknet_4_2_0_clk),
    .D(net41),
    .RESET_B(net9),
    .Q(\conv1.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1055_ (.CLK(clknet_4_3_0_clk),
    .D(net148),
    .RESET_B(net10),
    .Q(\conv1.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1056_ (.CLK(clknet_4_2_0_clk),
    .D(_0000_),
    .RESET_B(net9),
    .Q(\conv1.done ));
 sky130_fd_sc_hd__dfrtp_1 _1057_ (.CLK(clknet_4_2_0_clk),
    .D(_0001_),
    .RESET_B(net9),
    .Q(\conv1.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(clknet_4_15_0_clk),
    .D(_0040_),
    .Q(\mfcc.dct.output_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(clknet_4_15_0_clk),
    .D(_0041_),
    .Q(\mfcc.dct.output_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_4_15_0_clk),
    .D(_0042_),
    .Q(\mfcc.dct.output_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_4_14_0_clk),
    .D(_0043_),
    .Q(\mfcc.dct.output_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_4_14_0_clk),
    .D(_0044_),
    .Q(\mfcc.dct.output_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_4_14_0_clk),
    .D(_0045_),
    .Q(\mfcc.dct.output_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_4_15_0_clk),
    .D(_0046_),
    .Q(\mfcc.dct.input_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_4_15_0_clk),
    .D(_0047_),
    .Q(\mfcc.dct.input_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(clknet_4_15_0_clk),
    .D(_0048_),
    .Q(\mfcc.dct.input_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_4_15_0_clk),
    .D(_0049_),
    .Q(\mfcc.dct.input_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_4_15_0_clk),
    .D(_0050_),
    .Q(\mfcc.dct.input_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_4_14_0_clk),
    .D(_0051_),
    .Q(\mfcc.dct.dct_valid ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_4_13_0_clk),
    .D(_0052_),
    .Q(\mfcc.log.shift_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_4_12_0_clk),
    .D(_0053_),
    .Q(\mfcc.log.shift_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_4_12_0_clk),
    .D(_0054_),
    .Q(\mfcc.log.shift_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_4_12_0_clk),
    .D(_0055_),
    .Q(\mfcc.log.shift_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1074_ (.CLK(clknet_4_2_0_clk),
    .D(_0056_),
    .RESET_B(net9),
    .Q(\maxpool.addr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1075_ (.CLK(clknet_4_2_0_clk),
    .D(_0057_),
    .RESET_B(net9),
    .Q(\maxpool.addr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_4_15_0_clk),
    .D(net121),
    .Q(\mfcc.dct.data_valid ));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_4_13_0_clk),
    .D(_0059_),
    .Q(\mfcc.log.data_valid ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_4_13_0_clk),
    .D(_0060_),
    .Q(\mfcc.mel.filter_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_4_15_0_clk),
    .D(_0061_),
    .Q(\mfcc.mel.filter_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_4_13_0_clk),
    .D(_0062_),
    .Q(\mfcc.mel.filter_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_4_13_0_clk),
    .D(_0063_),
    .Q(\mfcc.mel.filter_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_4_7_0_clk),
    .D(_0064_),
    .Q(\mfcc.mel.filter_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_4_7_0_clk),
    .D(_0065_),
    .Q(\mfcc.mel.filter_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_4_7_0_clk),
    .D(_0066_),
    .Q(\mfcc.mel.coeff_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_4_7_0_clk),
    .D(_0067_),
    .Q(\mfcc.mel.coeff_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_4_7_0_clk),
    .D(_0068_),
    .Q(\mfcc.mel.coeff_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_4_13_0_clk),
    .D(_0069_),
    .Q(\mfcc.mel.coeff_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_4_7_0_clk),
    .D(_0070_),
    .Q(\mfcc.mel.coeff_counter[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1089_ (.CLK(clknet_4_8_0_clk),
    .D(_0071_),
    .RESET_B(net15),
    .Q(\maxpool.psram_ctrl.sck ));
 sky130_fd_sc_hd__dfrtp_1 _1090_ (.CLK(clknet_4_14_0_clk),
    .D(net30),
    .RESET_B(_0038_),
    .Q(\mfcc.mfcc_valid ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_4_15_0_clk),
    .D(net99),
    .Q(\mfcc.dct.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_4_15_0_clk),
    .D(_0023_),
    .Q(\mfcc.dct.state[1] ));
 sky130_fd_sc_hd__dfstp_1 _1093_ (.CLK(clknet_4_3_0_clk),
    .D(net80),
    .SET_B(net10),
    .Q(\conv2.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1094_ (.CLK(clknet_4_5_0_clk),
    .D(net35),
    .RESET_B(net12),
    .Q(\conv2.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1095_ (.CLK(clknet_4_3_0_clk),
    .D(_0015_),
    .RESET_B(net10),
    .Q(\conv2.state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1096_ (.CLK(clknet_4_4_0_clk),
    .D(_0002_),
    .RESET_B(net12),
    .Q(\conv2.data_out_valid ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_4_4_0_clk),
    .D(_0003_),
    .RESET_B(net11),
    .Q(\conv2.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1098_ (.CLK(clknet_4_0_0_clk),
    .D(net91),
    .RESET_B(net7),
    .Q(\conv1.psram_ctrl.has_wait_states ));
 sky130_fd_sc_hd__dfstp_1 _1099_ (.CLK(clknet_4_1_0_clk),
    .D(_0032_),
    .SET_B(net7),
    .Q(\conv1.psram_ce_n ));
 sky130_fd_sc_hd__dfrtp_2 _1100_ (.CLK(clknet_4_0_0_clk),
    .D(_0073_),
    .RESET_B(net7),
    .Q(\conv1.psram_ctrl.counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1101_ (.CLK(clknet_4_0_0_clk),
    .D(_0074_),
    .RESET_B(net7),
    .Q(\conv1.psram_ctrl.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_4_0_0_clk),
    .D(_0075_),
    .RESET_B(net7),
    .Q(\conv1.psram_ctrl.counter[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1103_ (.CLK(clknet_4_0_0_clk),
    .D(_0076_),
    .RESET_B(net7),
    .Q(\conv1.psram_ctrl.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1104_ (.CLK(clknet_4_0_0_clk),
    .D(_0077_),
    .RESET_B(net7),
    .Q(\conv1.psram_ctrl.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1105_ (.CLK(clknet_4_1_0_clk),
    .D(_0078_),
    .RESET_B(net8),
    .Q(\conv1.psram_ctrl.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1106_ (.CLK(clknet_4_1_0_clk),
    .D(net61),
    .RESET_B(net7),
    .Q(\conv1.psram_ctrl.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1107_ (.CLK(clknet_4_0_0_clk),
    .D(_0080_),
    .RESET_B(net7),
    .Q(\conv1.psram_ctrl.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1108_ (.CLK(clknet_4_2_0_clk),
    .D(\conv1.psram_ctrl.nstate ),
    .RESET_B(net9),
    .Q(\conv1.psram_ctrl.state ));
 sky130_fd_sc_hd__dfrtp_1 _1109_ (.CLK(clknet_4_0_0_clk),
    .D(_0031_),
    .RESET_B(net9),
    .Q(\conv1.psram_ctrl.start ));
 sky130_fd_sc_hd__dfstp_1 _1110_ (.CLK(clknet_4_3_0_clk),
    .D(net46),
    .SET_B(net19),
    .Q(\fc2.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1111_ (.CLK(clknet_4_12_0_clk),
    .D(net39),
    .RESET_B(net19),
    .Q(\fc2.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_4_6_0_clk),
    .D(net71),
    .RESET_B(net19),
    .Q(\fc2.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1113_ (.CLK(clknet_4_6_0_clk),
    .D(_0006_),
    .RESET_B(net12),
    .Q(\fc2.done ));
 sky130_fd_sc_hd__dfrtp_1 _1114_ (.CLK(clknet_4_12_0_clk),
    .D(_0007_),
    .RESET_B(net19),
    .Q(\fc2.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_4_13_0_clk),
    .D(net54),
    .Q(\mfcc.log.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_4_13_0_clk),
    .D(_0008_),
    .Q(\mfcc.log.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_4_13_0_clk),
    .D(_0009_),
    .Q(\mfcc.log.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_4_7_0_clk),
    .D(_0025_),
    .Q(\mfcc.mel.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_4_7_0_clk),
    .D(_0026_),
    .Q(\mfcc.mel.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_4_4_0_clk),
    .D(net75),
    .RESET_B(net12),
    .Q(\conv2.psram_ctrl.has_wait_states ));
 sky130_fd_sc_hd__dfstp_1 _1121_ (.CLK(clknet_4_1_0_clk),
    .D(_0033_),
    .SET_B(net8),
    .Q(\conv2.psram_ce_n ));
 sky130_fd_sc_hd__dfrtp_4 _1122_ (.CLK(clknet_4_4_0_clk),
    .D(_0082_),
    .RESET_B(net11),
    .Q(\conv2.psram_ctrl.counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1123_ (.CLK(clknet_4_4_0_clk),
    .D(_0083_),
    .RESET_B(net11),
    .Q(\conv2.psram_ctrl.counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1124_ (.CLK(clknet_4_4_0_clk),
    .D(_0084_),
    .RESET_B(net11),
    .Q(\conv2.psram_ctrl.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_4_4_0_clk),
    .D(_0085_),
    .RESET_B(net11),
    .Q(\conv2.psram_ctrl.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_4_1_0_clk),
    .D(_0086_),
    .RESET_B(net8),
    .Q(\conv2.psram_ctrl.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_4_1_0_clk),
    .D(_0087_),
    .RESET_B(net8),
    .Q(\conv2.psram_ctrl.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_4_1_0_clk),
    .D(net65),
    .RESET_B(net8),
    .Q(\conv2.psram_ctrl.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(clknet_4_1_0_clk),
    .D(_0089_),
    .RESET_B(net8),
    .Q(\conv2.psram_ctrl.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(clknet_4_5_0_clk),
    .D(\conv2.psram_ctrl.nstate ),
    .RESET_B(net11),
    .Q(\conv2.psram_ctrl.state ));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(clknet_4_4_0_clk),
    .D(_0030_),
    .RESET_B(net11),
    .Q(\conv2.psram_ctrl.start ));
 sky130_fd_sc_hd__dfrtp_1 _1132_ (.CLK(clknet_4_0_0_clk),
    .D(net85),
    .RESET_B(net7),
    .Q(\conv1.addr[8] ));
 sky130_fd_sc_hd__dfrtp_4 _1133_ (.CLK(clknet_4_0_0_clk),
    .D(_0091_),
    .RESET_B(net8),
    .Q(\conv1.psram_ctrl.sck ));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(clknet_4_9_0_clk),
    .D(net107),
    .RESET_B(net19),
    .Q(\fc1.psram_ctrl.has_wait_states ));
 sky130_fd_sc_hd__dfstp_1 _1135_ (.CLK(clknet_4_11_0_clk),
    .D(_0034_),
    .SET_B(net21),
    .Q(\fc1.psram_ce_n ));
 sky130_fd_sc_hd__dfrtp_4 _1136_ (.CLK(clknet_4_14_0_clk),
    .D(_0093_),
    .RESET_B(net22),
    .Q(\fc1.psram_ctrl.counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1137_ (.CLK(clknet_4_14_0_clk),
    .D(net118),
    .RESET_B(net21),
    .Q(\fc1.psram_ctrl.counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1138_ (.CLK(clknet_4_14_0_clk),
    .D(_0095_),
    .RESET_B(net21),
    .Q(\fc1.psram_ctrl.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(clknet_4_14_0_clk),
    .D(_0096_),
    .RESET_B(net21),
    .Q(\fc1.psram_ctrl.counter[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1140_ (.CLK(clknet_4_11_0_clk),
    .D(_0097_),
    .RESET_B(net21),
    .Q(\fc1.psram_ctrl.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1141_ (.CLK(clknet_4_11_0_clk),
    .D(_0098_),
    .RESET_B(net16),
    .Q(\fc1.psram_ctrl.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1142_ (.CLK(clknet_4_11_0_clk),
    .D(_0099_),
    .RESET_B(net17),
    .Q(\fc1.psram_ctrl.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1143_ (.CLK(clknet_4_11_0_clk),
    .D(_0100_),
    .RESET_B(net17),
    .Q(\fc1.psram_ctrl.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1144_ (.CLK(clknet_4_11_0_clk),
    .D(\fc1.psram_ctrl.nstate ),
    .RESET_B(net21),
    .Q(\fc1.psram_ctrl.state ));
 sky130_fd_sc_hd__dfrtp_1 _1145_ (.CLK(clknet_4_9_0_clk),
    .D(_0029_),
    .RESET_B(net21),
    .Q(\fc1.psram_ctrl.start ));
 sky130_fd_sc_hd__dfrtp_1 _1146_ (.CLK(clknet_4_5_0_clk),
    .D(net114),
    .RESET_B(net11),
    .Q(\conv2.addr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1147_ (.CLK(clknet_4_5_0_clk),
    .D(_0102_),
    .RESET_B(net11),
    .Q(\conv2.addr[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1148_ (.CLK(clknet_4_1_0_clk),
    .D(_0103_),
    .RESET_B(net10),
    .Q(\conv2.psram_ctrl.sck ));
 sky130_fd_sc_hd__dfrtp_4 _1149_ (.CLK(clknet_4_9_0_clk),
    .D(_0104_),
    .RESET_B(net18),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1150_ (.CLK(clknet_4_9_0_clk),
    .D(_0105_),
    .RESET_B(net18),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1151_ (.CLK(clknet_4_8_0_clk),
    .D(_0106_),
    .RESET_B(net18),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1152_ (.CLK(clknet_4_6_0_clk),
    .D(_0107_),
    .RESET_B(net12),
    .Q(\fc2.psram_ctrl.has_wait_states ));
 sky130_fd_sc_hd__dfstp_1 _1153_ (.CLK(clknet_4_6_0_clk),
    .D(_0035_),
    .SET_B(net12),
    .Q(\fc2.psram_ce_n ));
 sky130_fd_sc_hd__dfrtp_1 _1154_ (.CLK(clknet_4_7_0_clk),
    .D(_0108_),
    .RESET_B(net13),
    .Q(\fc2.psram_ctrl.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1155_ (.CLK(clknet_4_12_0_clk),
    .D(_0109_),
    .RESET_B(net13),
    .Q(\fc2.psram_ctrl.counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1156_ (.CLK(clknet_4_6_0_clk),
    .D(_0110_),
    .RESET_B(net13),
    .Q(\fc2.psram_ctrl.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1157_ (.CLK(clknet_4_6_0_clk),
    .D(_0111_),
    .RESET_B(net13),
    .Q(\fc2.psram_ctrl.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1158_ (.CLK(clknet_4_7_0_clk),
    .D(_0112_),
    .RESET_B(net13),
    .Q(\fc2.psram_ctrl.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1159_ (.CLK(clknet_4_7_0_clk),
    .D(_0113_),
    .RESET_B(net13),
    .Q(\fc2.psram_ctrl.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1160_ (.CLK(clknet_4_5_0_clk),
    .D(_0114_),
    .RESET_B(net11),
    .Q(\fc2.psram_ctrl.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1161_ (.CLK(clknet_4_5_0_clk),
    .D(_0115_),
    .RESET_B(net14),
    .Q(\fc2.psram_ctrl.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1162_ (.CLK(clknet_4_6_0_clk),
    .D(\fc2.psram_ctrl.nstate ),
    .RESET_B(net12),
    .Q(\fc2.psram_ctrl.state ));
 sky130_fd_sc_hd__dfrtp_1 _1163_ (.CLK(clknet_4_6_0_clk),
    .D(_0028_),
    .RESET_B(net12),
    .Q(\fc2.psram_ctrl.start ));
 sky130_fd_sc_hd__dfrtp_1 _1164_ (.CLK(clknet_4_14_0_clk),
    .D(net78),
    .RESET_B(net21),
    .Q(\fc1.addr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1165_ (.CLK(clknet_4_14_0_clk),
    .D(_0117_),
    .RESET_B(net21),
    .Q(\fc1.addr[10] ));
 sky130_fd_sc_hd__dfrtp_2 _1166_ (.CLK(clknet_4_11_0_clk),
    .D(_0118_),
    .RESET_B(net17),
    .Q(\fc1.psram_ctrl.sck ));
 sky130_fd_sc_hd__dfstp_1 _1167_ (.CLK(clknet_4_9_0_clk),
    .D(net112),
    .SET_B(net19),
    .Q(\fc1.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1168_ (.CLK(clknet_4_12_0_clk),
    .D(net37),
    .RESET_B(net19),
    .Q(\fc1.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1169_ (.CLK(clknet_4_9_0_clk),
    .D(_0018_),
    .RESET_B(net19),
    .Q(\fc1.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1170_ (.CLK(clknet_4_9_0_clk),
    .D(_0004_),
    .RESET_B(net19),
    .Q(\fc1.data_out_valid ));
 sky130_fd_sc_hd__dfrtp_1 _1171_ (.CLK(clknet_4_12_0_clk),
    .D(_0005_),
    .RESET_B(net20),
    .Q(\fc1.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1172_ (.CLK(clknet_4_3_0_clk),
    .D(_0119_),
    .RESET_B(net10),
    .Q(\maxpool.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1173_ (.CLK(clknet_4_3_0_clk),
    .D(_0120_),
    .RESET_B(net10),
    .Q(\maxpool.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1174_ (.CLK(clknet_4_3_0_clk),
    .D(_0121_),
    .RESET_B(net14),
    .Q(\maxpool.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _1175_ (.CLK(clknet_4_2_0_clk),
    .D(_0036_),
    .SET_B(net15),
    .Q(\maxpool.psram_ce_n ));
 sky130_fd_sc_hd__dfrtp_4 _1176_ (.CLK(clknet_4_2_0_clk),
    .D(_0122_),
    .RESET_B(net9),
    .Q(\maxpool.psram_ctrl.counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1177_ (.CLK(clknet_4_2_0_clk),
    .D(net102),
    .RESET_B(net9),
    .Q(\maxpool.psram_ctrl.counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1178_ (.CLK(clknet_4_2_0_clk),
    .D(_0124_),
    .RESET_B(net10),
    .Q(\maxpool.psram_ctrl.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1179_ (.CLK(clknet_4_2_0_clk),
    .D(_0125_),
    .RESET_B(net15),
    .Q(\maxpool.psram_ctrl.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1180_ (.CLK(clknet_4_8_0_clk),
    .D(_0126_),
    .RESET_B(net15),
    .Q(\maxpool.psram_ctrl.counter[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1181_ (.CLK(clknet_4_8_0_clk),
    .D(_0127_),
    .RESET_B(net15),
    .Q(\maxpool.psram_ctrl.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1182_ (.CLK(clknet_4_8_0_clk),
    .D(net140),
    .RESET_B(net15),
    .Q(\maxpool.psram_ctrl.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1183_ (.CLK(clknet_4_10_0_clk),
    .D(_0129_),
    .RESET_B(net15),
    .Q(\maxpool.psram_ctrl.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1184_ (.CLK(clknet_4_2_0_clk),
    .D(\maxpool.psram_ctrl.nstate ),
    .RESET_B(net15),
    .Q(\maxpool.psram_ctrl.state ));
 sky130_fd_sc_hd__dfrtp_1 _1185_ (.CLK(clknet_4_12_0_clk),
    .D(net88),
    .RESET_B(net20),
    .Q(\fc2.addr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1186_ (.CLK(clknet_4_12_0_clk),
    .D(_0131_),
    .RESET_B(net20),
    .Q(\fc2.addr[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1187_ (.CLK(clknet_4_2_0_clk),
    .D(_0027_),
    .RESET_B(net10),
    .Q(\maxpool.psram_ctrl.start ));
 sky130_fd_sc_hd__dfrtp_1 _1188_ (.CLK(clknet_4_3_0_clk),
    .D(_0132_),
    .RESET_B(net14),
    .Q(\fc2.psram_ctrl.sck ));
 sky130_fd_sc_hd__dfrtp_1 _1189_ (.CLK(clknet_4_10_0_clk),
    .D(net33),
    .RESET_B(net16),
    .Q(\softmax.addr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1190_ (.CLK(clknet_4_10_0_clk),
    .D(_0134_),
    .RESET_B(net16),
    .Q(\softmax.addr[11] ));
 sky130_fd_sc_hd__dfstp_1 _1191_ (.CLK(clknet_4_10_0_clk),
    .D(_0037_),
    .SET_B(net17),
    .Q(\softmax.psram_ce_n ));
 sky130_fd_sc_hd__dfrtp_4 _1192_ (.CLK(clknet_4_10_0_clk),
    .D(_0135_),
    .RESET_B(net16),
    .Q(\softmax.psram_ctrl.counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1193_ (.CLK(clknet_4_10_0_clk),
    .D(_0136_),
    .RESET_B(net16),
    .Q(\softmax.psram_ctrl.counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1194_ (.CLK(clknet_4_10_0_clk),
    .D(_0137_),
    .RESET_B(net16),
    .Q(\softmax.psram_ctrl.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1195_ (.CLK(clknet_4_10_0_clk),
    .D(_0138_),
    .RESET_B(net16),
    .Q(\softmax.psram_ctrl.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1196_ (.CLK(clknet_4_10_0_clk),
    .D(_0139_),
    .RESET_B(net16),
    .Q(\softmax.psram_ctrl.counter[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1197_ (.CLK(clknet_4_10_0_clk),
    .D(_0140_),
    .RESET_B(net17),
    .Q(\softmax.psram_ctrl.counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _1198_ (.CLK(clknet_4_10_0_clk),
    .D(_0141_),
    .RESET_B(net17),
    .Q(\softmax.psram_ctrl.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1199_ (.CLK(clknet_4_10_0_clk),
    .D(_0142_),
    .RESET_B(net17),
    .Q(\softmax.psram_ctrl.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1200_ (.CLK(clknet_4_10_0_clk),
    .D(\softmax.psram_ctrl.nstate ),
    .RESET_B(net16),
    .Q(\softmax.psram_ctrl.state ));
 sky130_fd_sc_hd__dfrtp_1 _1201_ (.CLK(clknet_4_8_0_clk),
    .D(_0143_),
    .RESET_B(net15),
    .Q(\softmax.psram_ctrl.start ));
 sky130_fd_sc_hd__dfrtp_1 _1202_ (.CLK(clknet_4_8_0_clk),
    .D(_0144_),
    .RESET_B(net15),
    .Q(\softmax.data_valid ));
 sky130_fd_sc_hd__dfrtp_1 _1203_ (.CLK(clknet_4_12_0_clk),
    .D(_0145_),
    .RESET_B(net20),
    .Q(\fc1.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1204_ (.CLK(clknet_4_12_0_clk),
    .D(_0146_),
    .RESET_B(net19),
    .Q(\fc2.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1205_ (.CLK(clknet_4_4_0_clk),
    .D(_0147_),
    .RESET_B(net12),
    .Q(\conv2.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1206_ (.CLK(clknet_4_0_0_clk),
    .D(_0148_),
    .RESET_B(net9),
    .Q(\conv1.state[2] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__conb_1 cnn_kws_accel_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 cnn_kws_accel_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 cnn_kws_accel_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 cnn_kws_accel_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 cnn_kws_accel_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 cnn_kws_accel_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 cnn_kws_accel_29 (.HI(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net14),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 fanout11 (.A(net14),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net14),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net1),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net18),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net18),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net18),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 fanout18 (.A(net22),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net22),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(net1),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(net8),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net14),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\mfcc.dct.dct_valid ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0020_),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\conv2.state[0] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\fc2.state[1] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\maxpool.psram_ctrl.start ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\fc2.psram_ctrl.has_wait_states ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\fc2.psram_ctrl.counter[2] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\conv1.psram_ctrl.counter[1] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\softmax.addr[11] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\maxpool.psram_ce_n ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\softmax.psram_ctrl.counter[3] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\maxpool.state[1] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\conv1.state[5] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\maxpool.psram_ctrl.counter[6] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0128_),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\softmax.psram_ctrl.counter[6] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\state[1] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\fc1.addr[10] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\fc2.psram_ctrl.counter[1] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\mfcc.mel.coeff_counter[1] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\softmax.psram_ctrl.sck ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\conv1.state[3] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0012_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0011_),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\fc2.psram_ctrl.counter[3] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\conv1.state[1] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\conv2.psram_ctrl.counter[3] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\maxpool.psram_ctrl.counter[3] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\maxpool.psram_ctrl.counter[2] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\conv2.psram_ctrl.sck ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\state[2] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\fc1.psram_ctrl.counter[2] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\conv1.psram_ctrl.counter[2] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\mfcc.dct.input_counter[1] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\fc1.psram_ctrl.state ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\fc1.psram_ctrl.counter[3] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\softmax.psram_ctrl.counter[2] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\maxpool.addr[8] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\fc2.psram_ctrl.counter[5] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\fc1.psram_ctrl.counter[4] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\fc1.state[2] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\fc2.psram_ctrl.counter[4] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\conv2.state[3] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\softmax.data_valid ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\mfcc.dct.input_counter[2] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\fc2.psram_ctrl.state ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\maxpool.psram_ctrl.state ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\fc2.done ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0019_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\conv1.psram_ctrl.state ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\mfcc.mel.state[0] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\conv2.psram_ctrl.state ),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\mfcc.dct.input_counter[4] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\mfcc.dct.output_counter[4] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\mfcc.log.shift_count[3] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\softmax.psram_ctrl.state ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\mfcc.log.state[0] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0024_),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\conv1.done ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0010_),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\mfcc.dct.output_counter[2] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\maxpool.state[2] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\softmax.data_valid ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\mfcc.mel.coeff_counter[4] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\conv1.psram_ctrl.counter[6] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0079_),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\fc1.psram_ctrl.counter[6] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\mfcc.dct.output_counter[5] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\conv2.psram_ctrl.counter[6] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0088_),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\mfcc.mel.filter_counter[2] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\mfcc.log.shift_count[1] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\mfcc.dct.input_counter[0] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0133_),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\conv2.state[1] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\fc2.state[3] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0021_),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\mfcc.dct.input_counter[3] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\mfcc.log.data_valid ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\conv2.state[3] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0081_),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\mfcc.mel.coeff_counter[3] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\fc1.state[2] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0116_),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\conv2.state[5] ),
    .X(net34));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold50 (.A(\conv2.data_out_valid ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0013_),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\softmax.psram_ctrl.start ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\mfcc.log.shift_count[0] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\conv2.psram_ctrl.counter[7] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\conv1.addr[8] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0090_),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\fc1.psram_ctrl.counter[7] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\fc2.state[2] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0130_),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0014_),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\conv1.psram_ctrl.start ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\conv1.psram_ctrl.has_wait_states ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0072_),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\fc1.psram_ctrl.start ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\conv1.psram_ctrl.counter[4] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\conv1.state[2] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\conv1.psram_ctrl.counter[7] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\mfcc.log.shift_count[2] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0337_),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\mfcc.dct.state[0] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\fc1.state[5] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0022_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\softmax.psram_ctrl.counter[4] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\maxpool.psram_ctrl.sck ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0123_),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\conv2.psram_ctrl.counter[4] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\mfcc.dct.output_counter[0] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\mfcc.mel.filter_counter[1] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\fc1.state[3] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0092_),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\fc1.state[0] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0017_),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\fc2.psram_ctrl.counter[6] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\mfcc.dct.output_counter[3] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\fc1.data_out_valid ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0016_),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\conv2.state[2] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0101_),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\mfcc.mel.filter_counter[0] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\fc2.psram_ctrl.start ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\fc1.psram_ctrl.sck ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0094_),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\fc2.state[5] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\mfcc.dct.input_counter[2] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\mfcc.dct.data_valid ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0058_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\conv2.addr[9] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\maxpool.psram_ctrl.counter[4] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\conv2.psram_ctrl.start ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\fc1.state[1] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\fc2.addr[10] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\mfcc.mel.filter_counter[4] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\maxpool.addr[11] ),
    .X(net128));
 sky130_fd_sc_hd__buf_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(start),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 output3 (.A(net3),
    .X(done));
 sky130_fd_sc_hd__clkbuf_4 output4 (.A(net4),
    .X(psram_ce_n));
 sky130_fd_sc_hd__clkbuf_4 output5 (.A(net5),
    .X(psram_sck));
 sky130_fd_sc_hd__buf_1 wire6 (.A(_0373_),
    .X(net6));
 assign psram_d[1] = net23;
 assign psram_d[2] = net24;
 assign psram_d[3] = net25;
 assign psram_douten[0] = net29;
 assign psram_douten[1] = net26;
 assign psram_douten[2] = net27;
 assign psram_douten[3] = net28;
endmodule

