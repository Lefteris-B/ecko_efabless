VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -38.270 12.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -38.270 192.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -38.270 372.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -38.270 552.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -38.270 732.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -38.270 912.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -38.270 1092.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -38.270 1272.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -38.270 1452.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -38.270 1632.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -38.270 1812.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -38.270 1992.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -38.270 2172.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -38.270 2352.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -38.270 2532.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -38.270 2712.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -38.270 2892.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 14.330 2963.250 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 194.330 2963.250 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 374.330 2963.250 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 554.330 2963.250 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 734.330 2963.250 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 914.330 2963.250 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1094.330 2963.250 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1274.330 2963.250 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1454.330 2963.250 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1634.330 2963.250 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1814.330 2963.250 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1994.330 2963.250 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2174.330 2963.250 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2354.330 2963.250 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2534.330 2963.250 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2714.330 2963.250 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2894.330 2963.250 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3074.330 2963.250 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3254.330 2963.250 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3434.330 2963.250 3437.430 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -38.270 49.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 -38.270 229.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 -38.270 409.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 -38.270 589.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 -38.270 769.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 -38.270 949.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 -38.270 1129.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 -38.270 1309.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 -38.270 1489.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 -38.270 1669.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 -38.270 1849.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 -38.270 2029.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 -38.270 2209.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 -38.270 2389.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 -38.270 2569.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 -38.270 2749.270 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 51.530 2963.250 54.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 231.530 2963.250 234.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 411.530 2963.250 414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 591.530 2963.250 594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 771.530 2963.250 774.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 951.530 2963.250 954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1131.530 2963.250 1134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1311.530 2963.250 1314.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1491.530 2963.250 1494.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1671.530 2963.250 1674.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1851.530 2963.250 1854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2031.530 2963.250 2034.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2211.530 2963.250 2214.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2391.530 2963.250 2394.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2571.530 2963.250 2574.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2751.530 2963.250 2754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2931.530 2963.250 2934.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3111.530 2963.250 3114.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3291.530 2963.250 3294.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3471.530 2963.250 3474.630 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.370 -38.270 86.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.370 -38.270 266.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.370 -38.270 446.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.370 -38.270 626.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.370 -38.270 806.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 983.370 -38.270 986.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1163.370 -38.270 1166.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1343.370 -38.270 1346.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.370 -38.270 1526.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1703.370 -38.270 1706.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1883.370 -38.270 1886.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2063.370 -38.270 2066.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2243.370 -38.270 2246.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.370 -38.270 2426.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2603.370 -38.270 2606.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2783.370 -38.270 2786.470 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 88.730 2963.250 91.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 268.730 2963.250 271.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 448.730 2963.250 451.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 628.730 2963.250 631.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 808.730 2963.250 811.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 988.730 2963.250 991.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1168.730 2963.250 1171.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1348.730 2963.250 1351.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1528.730 2963.250 1531.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1708.730 2963.250 1711.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1888.730 2963.250 1891.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2068.730 2963.250 2071.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2248.730 2963.250 2251.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2428.730 2963.250 2431.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2608.730 2963.250 2611.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2788.730 2963.250 2791.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2968.730 2963.250 2971.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3148.730 2963.250 3151.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3328.730 2963.250 3331.830 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.570 -38.270 123.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 300.570 -38.270 303.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 480.570 -38.270 483.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 660.570 -38.270 663.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 840.570 -38.270 843.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1020.570 -38.270 1023.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1200.570 -38.270 1203.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1380.570 -38.270 1383.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1560.570 -38.270 1563.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1740.570 -38.270 1743.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1920.570 -38.270 1923.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2100.570 -38.270 2103.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2280.570 -38.270 2283.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2460.570 -38.270 2463.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2640.570 -38.270 2643.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2820.570 -38.270 2823.670 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 125.930 2963.250 129.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 305.930 2963.250 309.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 485.930 2963.250 489.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 665.930 2963.250 669.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 845.930 2963.250 849.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1025.930 2963.250 1029.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1205.930 2963.250 1209.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1385.930 2963.250 1389.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1565.930 2963.250 1569.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1745.930 2963.250 1749.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1925.930 2963.250 1929.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2105.930 2963.250 2109.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2285.930 2963.250 2289.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2465.930 2963.250 2469.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2645.930 2963.250 2649.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2825.930 2963.250 2829.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3005.930 2963.250 3009.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3185.930 2963.250 3189.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3365.930 2963.250 3369.030 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.970 -38.270 105.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 281.970 -38.270 285.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.970 -38.270 465.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 641.970 -38.270 645.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.970 -38.270 825.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.970 -38.270 1005.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1181.970 -38.270 1185.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1361.970 -38.270 1365.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1541.970 -38.270 1545.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.970 -38.270 1725.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1901.970 -38.270 1905.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2081.970 -38.270 2085.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2261.970 -38.270 2265.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2441.970 -38.270 2445.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2621.970 -38.270 2625.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2801.970 -38.270 2805.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 107.330 2963.250 110.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 287.330 2963.250 290.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 467.330 2963.250 470.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 647.330 2963.250 650.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 827.330 2963.250 830.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1007.330 2963.250 1010.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1187.330 2963.250 1190.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1367.330 2963.250 1370.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1547.330 2963.250 1550.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1727.330 2963.250 1730.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1907.330 2963.250 1910.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2087.330 2963.250 2090.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2267.330 2963.250 2270.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2447.330 2963.250 2450.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2627.330 2963.250 2630.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2807.330 2963.250 2810.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2987.330 2963.250 2990.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3167.330 2963.250 3170.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3347.330 2963.250 3350.430 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.170 -38.270 142.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.170 -38.270 322.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 499.170 -38.270 502.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.170 -38.270 682.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 859.170 -38.270 862.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1039.170 -38.270 1042.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1219.170 -38.270 1222.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1399.170 -38.270 1402.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1579.170 -38.270 1582.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1759.170 -38.270 1762.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1939.170 -38.270 1942.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2119.170 -38.270 2122.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2299.170 -38.270 2302.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2479.170 -38.270 2482.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2659.170 -38.270 2662.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2839.170 -38.270 2842.270 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 144.530 2963.250 147.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 324.530 2963.250 327.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 504.530 2963.250 507.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 684.530 2963.250 687.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 864.530 2963.250 867.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1044.530 2963.250 1047.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1224.530 2963.250 1227.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1404.530 2963.250 1407.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1584.530 2963.250 1587.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1764.530 2963.250 1767.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1944.530 2963.250 1947.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2124.530 2963.250 2127.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2304.530 2963.250 2307.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2484.530 2963.250 2487.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2664.530 2963.250 2667.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2844.530 2963.250 2847.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3024.530 2963.250 3027.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3204.530 2963.250 3207.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3384.530 2963.250 3387.630 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -38.270 30.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 -38.270 210.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 363.220 390.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 -38.270 570.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 -38.270 750.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 -38.270 930.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 -38.270 1110.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 -38.270 1290.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 -38.270 1470.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 -38.270 1650.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 -38.270 1830.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 -38.270 2010.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 -38.270 2190.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 -38.270 2370.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 -38.270 2550.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 -38.270 2730.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.570 -38.270 2910.670 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 32.930 2963.250 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 212.930 2963.250 216.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 392.930 2963.250 396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 572.930 2963.250 576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 752.930 2963.250 756.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 932.930 2963.250 936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1112.930 2963.250 1116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1292.930 2963.250 1296.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1472.930 2963.250 1476.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1652.930 2963.250 1656.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1832.930 2963.250 1836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2012.930 2963.250 2016.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2192.930 2963.250 2196.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2372.930 2963.250 2376.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2552.930 2963.250 2556.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2732.930 2963.250 2736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2912.930 2963.250 2916.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3092.930 2963.250 3096.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3272.930 2963.250 3276.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3452.930 2963.250 3456.030 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 -38.270 247.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 -38.270 427.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 -38.270 607.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 -38.270 787.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 -38.270 967.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 -38.270 1147.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 -38.270 1327.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 -38.270 1507.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 -38.270 1687.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 -38.270 1867.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 -38.270 2047.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 -38.270 2227.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 -38.270 2407.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 -38.270 2587.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 -38.270 2767.870 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 250.130 2963.250 253.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 430.130 2963.250 433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 610.130 2963.250 613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 790.130 2963.250 793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.130 2963.250 973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 65.520 25.795 404.080 352.365 ;
      LAYER met1 ;
        RECT 64.670 25.640 404.470 352.520 ;
      LAYER met2 ;
        RECT 2.850 3517.320 40.150 3517.600 ;
        RECT 41.270 3517.320 121.110 3517.600 ;
        RECT 122.230 3517.320 202.070 3517.600 ;
        RECT 203.190 3517.320 283.490 3517.600 ;
        RECT 284.610 3517.320 364.450 3517.600 ;
        RECT 365.570 3517.320 445.410 3517.600 ;
        RECT 446.530 3517.320 526.830 3517.600 ;
        RECT 527.950 3517.320 607.790 3517.600 ;
        RECT 608.910 3517.320 688.750 3517.600 ;
        RECT 689.870 3517.320 770.170 3517.600 ;
        RECT 771.290 3517.320 851.130 3517.600 ;
        RECT 852.250 3517.320 932.090 3517.600 ;
        RECT 933.210 3517.320 1013.510 3517.600 ;
        RECT 1014.630 3517.320 1094.470 3517.600 ;
        RECT 1095.590 3517.320 1175.430 3517.600 ;
        RECT 1176.550 3517.320 1256.850 3517.600 ;
        RECT 1257.970 3517.320 1337.810 3517.600 ;
        RECT 1338.930 3517.320 1418.770 3517.600 ;
        RECT 1419.890 3517.320 1500.190 3517.600 ;
        RECT 1501.310 3517.320 1581.150 3517.600 ;
        RECT 1582.270 3517.320 1662.110 3517.600 ;
        RECT 1663.230 3517.320 1743.530 3517.600 ;
        RECT 1744.650 3517.320 1824.490 3517.600 ;
        RECT 1825.610 3517.320 1905.450 3517.600 ;
        RECT 1906.570 3517.320 1986.870 3517.600 ;
        RECT 1987.990 3517.320 2067.830 3517.600 ;
        RECT 2068.950 3517.320 2148.790 3517.600 ;
        RECT 2149.910 3517.320 2230.210 3517.600 ;
        RECT 2231.330 3517.320 2311.170 3517.600 ;
        RECT 2312.290 3517.320 2392.130 3517.600 ;
        RECT 2393.250 3517.320 2473.550 3517.600 ;
        RECT 2474.670 3517.320 2554.510 3517.600 ;
        RECT 2555.630 3517.320 2635.470 3517.600 ;
        RECT 2636.590 3517.320 2716.890 3517.600 ;
        RECT 2718.010 3517.320 2797.850 3517.600 ;
        RECT 2798.970 3517.320 2878.810 3517.600 ;
        RECT 2879.930 3517.320 2903.890 3517.600 ;
        RECT 2.850 2.680 2903.890 3517.320 ;
        RECT 3.550 2.400 7.950 2.680 ;
        RECT 9.070 2.400 13.930 2.680 ;
        RECT 15.050 2.400 19.910 2.680 ;
        RECT 21.030 2.400 25.890 2.680 ;
        RECT 27.010 2.400 31.870 2.680 ;
        RECT 32.990 2.400 37.850 2.680 ;
        RECT 38.970 2.400 43.370 2.680 ;
        RECT 44.490 2.400 49.350 2.680 ;
        RECT 50.470 2.400 55.330 2.680 ;
        RECT 56.450 2.400 61.310 2.680 ;
        RECT 62.430 2.400 67.290 2.680 ;
        RECT 68.410 2.400 73.270 2.680 ;
        RECT 74.390 2.400 79.250 2.680 ;
        RECT 80.370 2.400 84.770 2.680 ;
        RECT 85.890 2.400 90.750 2.680 ;
        RECT 91.870 2.400 96.730 2.680 ;
        RECT 97.850 2.400 102.710 2.680 ;
        RECT 103.830 2.400 108.690 2.680 ;
        RECT 109.810 2.400 114.670 2.680 ;
        RECT 115.790 2.400 120.650 2.680 ;
        RECT 121.770 2.400 126.170 2.680 ;
        RECT 127.290 2.400 132.150 2.680 ;
        RECT 133.270 2.400 138.130 2.680 ;
        RECT 139.250 2.400 144.110 2.680 ;
        RECT 145.230 2.400 150.090 2.680 ;
        RECT 151.210 2.400 156.070 2.680 ;
        RECT 157.190 2.400 161.590 2.680 ;
        RECT 162.710 2.400 167.570 2.680 ;
        RECT 168.690 2.400 173.550 2.680 ;
        RECT 174.670 2.400 179.530 2.680 ;
        RECT 180.650 2.400 185.510 2.680 ;
        RECT 186.630 2.400 191.490 2.680 ;
        RECT 192.610 2.400 197.470 2.680 ;
        RECT 198.590 2.400 202.990 2.680 ;
        RECT 204.110 2.400 208.970 2.680 ;
        RECT 210.090 2.400 214.950 2.680 ;
        RECT 216.070 2.400 220.930 2.680 ;
        RECT 222.050 2.400 226.910 2.680 ;
        RECT 228.030 2.400 232.890 2.680 ;
        RECT 234.010 2.400 238.870 2.680 ;
        RECT 239.990 2.400 244.390 2.680 ;
        RECT 245.510 2.400 250.370 2.680 ;
        RECT 251.490 2.400 256.350 2.680 ;
        RECT 257.470 2.400 262.330 2.680 ;
        RECT 263.450 2.400 268.310 2.680 ;
        RECT 269.430 2.400 274.290 2.680 ;
        RECT 275.410 2.400 279.810 2.680 ;
        RECT 280.930 2.400 285.790 2.680 ;
        RECT 286.910 2.400 291.770 2.680 ;
        RECT 292.890 2.400 297.750 2.680 ;
        RECT 298.870 2.400 303.730 2.680 ;
        RECT 304.850 2.400 309.710 2.680 ;
        RECT 310.830 2.400 315.690 2.680 ;
        RECT 316.810 2.400 321.210 2.680 ;
        RECT 322.330 2.400 327.190 2.680 ;
        RECT 328.310 2.400 333.170 2.680 ;
        RECT 334.290 2.400 339.150 2.680 ;
        RECT 340.270 2.400 345.130 2.680 ;
        RECT 346.250 2.400 351.110 2.680 ;
        RECT 352.230 2.400 357.090 2.680 ;
        RECT 358.210 2.400 362.610 2.680 ;
        RECT 363.730 2.400 368.590 2.680 ;
        RECT 369.710 2.400 374.570 2.680 ;
        RECT 375.690 2.400 380.550 2.680 ;
        RECT 381.670 2.400 386.530 2.680 ;
        RECT 387.650 2.400 392.510 2.680 ;
        RECT 393.630 2.400 398.030 2.680 ;
        RECT 399.150 2.400 404.010 2.680 ;
        RECT 405.130 2.400 409.990 2.680 ;
        RECT 411.110 2.400 415.970 2.680 ;
        RECT 417.090 2.400 421.950 2.680 ;
        RECT 423.070 2.400 427.930 2.680 ;
        RECT 429.050 2.400 433.910 2.680 ;
        RECT 435.030 2.400 439.430 2.680 ;
        RECT 440.550 2.400 445.410 2.680 ;
        RECT 446.530 2.400 451.390 2.680 ;
        RECT 452.510 2.400 457.370 2.680 ;
        RECT 458.490 2.400 463.350 2.680 ;
        RECT 464.470 2.400 469.330 2.680 ;
        RECT 470.450 2.400 475.310 2.680 ;
        RECT 476.430 2.400 480.830 2.680 ;
        RECT 481.950 2.400 486.810 2.680 ;
        RECT 487.930 2.400 492.790 2.680 ;
        RECT 493.910 2.400 498.770 2.680 ;
        RECT 499.890 2.400 504.750 2.680 ;
        RECT 505.870 2.400 510.730 2.680 ;
        RECT 511.850 2.400 516.250 2.680 ;
        RECT 517.370 2.400 522.230 2.680 ;
        RECT 523.350 2.400 528.210 2.680 ;
        RECT 529.330 2.400 534.190 2.680 ;
        RECT 535.310 2.400 540.170 2.680 ;
        RECT 541.290 2.400 546.150 2.680 ;
        RECT 547.270 2.400 552.130 2.680 ;
        RECT 553.250 2.400 557.650 2.680 ;
        RECT 558.770 2.400 563.630 2.680 ;
        RECT 564.750 2.400 569.610 2.680 ;
        RECT 570.730 2.400 575.590 2.680 ;
        RECT 576.710 2.400 581.570 2.680 ;
        RECT 582.690 2.400 587.550 2.680 ;
        RECT 588.670 2.400 593.530 2.680 ;
        RECT 594.650 2.400 599.050 2.680 ;
        RECT 600.170 2.400 605.030 2.680 ;
        RECT 606.150 2.400 611.010 2.680 ;
        RECT 612.130 2.400 616.990 2.680 ;
        RECT 618.110 2.400 622.970 2.680 ;
        RECT 624.090 2.400 628.950 2.680 ;
        RECT 630.070 2.400 634.470 2.680 ;
        RECT 635.590 2.400 640.450 2.680 ;
        RECT 641.570 2.400 646.430 2.680 ;
        RECT 647.550 2.400 652.410 2.680 ;
        RECT 653.530 2.400 658.390 2.680 ;
        RECT 659.510 2.400 664.370 2.680 ;
        RECT 665.490 2.400 670.350 2.680 ;
        RECT 671.470 2.400 675.870 2.680 ;
        RECT 676.990 2.400 681.850 2.680 ;
        RECT 682.970 2.400 687.830 2.680 ;
        RECT 688.950 2.400 693.810 2.680 ;
        RECT 694.930 2.400 699.790 2.680 ;
        RECT 700.910 2.400 705.770 2.680 ;
        RECT 706.890 2.400 711.750 2.680 ;
        RECT 712.870 2.400 717.270 2.680 ;
        RECT 718.390 2.400 723.250 2.680 ;
        RECT 724.370 2.400 729.230 2.680 ;
        RECT 730.350 2.400 735.210 2.680 ;
        RECT 736.330 2.400 741.190 2.680 ;
        RECT 742.310 2.400 747.170 2.680 ;
        RECT 748.290 2.400 752.690 2.680 ;
        RECT 753.810 2.400 758.670 2.680 ;
        RECT 759.790 2.400 764.650 2.680 ;
        RECT 765.770 2.400 770.630 2.680 ;
        RECT 771.750 2.400 776.610 2.680 ;
        RECT 777.730 2.400 782.590 2.680 ;
        RECT 783.710 2.400 788.570 2.680 ;
        RECT 789.690 2.400 794.090 2.680 ;
        RECT 795.210 2.400 800.070 2.680 ;
        RECT 801.190 2.400 806.050 2.680 ;
        RECT 807.170 2.400 812.030 2.680 ;
        RECT 813.150 2.400 818.010 2.680 ;
        RECT 819.130 2.400 823.990 2.680 ;
        RECT 825.110 2.400 829.970 2.680 ;
        RECT 831.090 2.400 835.490 2.680 ;
        RECT 836.610 2.400 841.470 2.680 ;
        RECT 842.590 2.400 847.450 2.680 ;
        RECT 848.570 2.400 853.430 2.680 ;
        RECT 854.550 2.400 859.410 2.680 ;
        RECT 860.530 2.400 865.390 2.680 ;
        RECT 866.510 2.400 870.910 2.680 ;
        RECT 872.030 2.400 876.890 2.680 ;
        RECT 878.010 2.400 882.870 2.680 ;
        RECT 883.990 2.400 888.850 2.680 ;
        RECT 889.970 2.400 894.830 2.680 ;
        RECT 895.950 2.400 900.810 2.680 ;
        RECT 901.930 2.400 906.790 2.680 ;
        RECT 907.910 2.400 912.310 2.680 ;
        RECT 913.430 2.400 918.290 2.680 ;
        RECT 919.410 2.400 924.270 2.680 ;
        RECT 925.390 2.400 930.250 2.680 ;
        RECT 931.370 2.400 936.230 2.680 ;
        RECT 937.350 2.400 942.210 2.680 ;
        RECT 943.330 2.400 948.190 2.680 ;
        RECT 949.310 2.400 953.710 2.680 ;
        RECT 954.830 2.400 959.690 2.680 ;
        RECT 960.810 2.400 965.670 2.680 ;
        RECT 966.790 2.400 971.650 2.680 ;
        RECT 972.770 2.400 977.630 2.680 ;
        RECT 978.750 2.400 983.610 2.680 ;
        RECT 984.730 2.400 989.130 2.680 ;
        RECT 990.250 2.400 995.110 2.680 ;
        RECT 996.230 2.400 1001.090 2.680 ;
        RECT 1002.210 2.400 1007.070 2.680 ;
        RECT 1008.190 2.400 1013.050 2.680 ;
        RECT 1014.170 2.400 1019.030 2.680 ;
        RECT 1020.150 2.400 1025.010 2.680 ;
        RECT 1026.130 2.400 1030.530 2.680 ;
        RECT 1031.650 2.400 1036.510 2.680 ;
        RECT 1037.630 2.400 1042.490 2.680 ;
        RECT 1043.610 2.400 1048.470 2.680 ;
        RECT 1049.590 2.400 1054.450 2.680 ;
        RECT 1055.570 2.400 1060.430 2.680 ;
        RECT 1061.550 2.400 1066.410 2.680 ;
        RECT 1067.530 2.400 1071.930 2.680 ;
        RECT 1073.050 2.400 1077.910 2.680 ;
        RECT 1079.030 2.400 1083.890 2.680 ;
        RECT 1085.010 2.400 1089.870 2.680 ;
        RECT 1090.990 2.400 1095.850 2.680 ;
        RECT 1096.970 2.400 1101.830 2.680 ;
        RECT 1102.950 2.400 1107.350 2.680 ;
        RECT 1108.470 2.400 1113.330 2.680 ;
        RECT 1114.450 2.400 1119.310 2.680 ;
        RECT 1120.430 2.400 1125.290 2.680 ;
        RECT 1126.410 2.400 1131.270 2.680 ;
        RECT 1132.390 2.400 1137.250 2.680 ;
        RECT 1138.370 2.400 1143.230 2.680 ;
        RECT 1144.350 2.400 1148.750 2.680 ;
        RECT 1149.870 2.400 1154.730 2.680 ;
        RECT 1155.850 2.400 1160.710 2.680 ;
        RECT 1161.830 2.400 1166.690 2.680 ;
        RECT 1167.810 2.400 1172.670 2.680 ;
        RECT 1173.790 2.400 1178.650 2.680 ;
        RECT 1179.770 2.400 1184.630 2.680 ;
        RECT 1185.750 2.400 1190.150 2.680 ;
        RECT 1191.270 2.400 1196.130 2.680 ;
        RECT 1197.250 2.400 1202.110 2.680 ;
        RECT 1203.230 2.400 1208.090 2.680 ;
        RECT 1209.210 2.400 1214.070 2.680 ;
        RECT 1215.190 2.400 1220.050 2.680 ;
        RECT 1221.170 2.400 1225.570 2.680 ;
        RECT 1226.690 2.400 1231.550 2.680 ;
        RECT 1232.670 2.400 1237.530 2.680 ;
        RECT 1238.650 2.400 1243.510 2.680 ;
        RECT 1244.630 2.400 1249.490 2.680 ;
        RECT 1250.610 2.400 1255.470 2.680 ;
        RECT 1256.590 2.400 1261.450 2.680 ;
        RECT 1262.570 2.400 1266.970 2.680 ;
        RECT 1268.090 2.400 1272.950 2.680 ;
        RECT 1274.070 2.400 1278.930 2.680 ;
        RECT 1280.050 2.400 1284.910 2.680 ;
        RECT 1286.030 2.400 1290.890 2.680 ;
        RECT 1292.010 2.400 1296.870 2.680 ;
        RECT 1297.990 2.400 1302.850 2.680 ;
        RECT 1303.970 2.400 1308.370 2.680 ;
        RECT 1309.490 2.400 1314.350 2.680 ;
        RECT 1315.470 2.400 1320.330 2.680 ;
        RECT 1321.450 2.400 1326.310 2.680 ;
        RECT 1327.430 2.400 1332.290 2.680 ;
        RECT 1333.410 2.400 1338.270 2.680 ;
        RECT 1339.390 2.400 1343.790 2.680 ;
        RECT 1344.910 2.400 1349.770 2.680 ;
        RECT 1350.890 2.400 1355.750 2.680 ;
        RECT 1356.870 2.400 1361.730 2.680 ;
        RECT 1362.850 2.400 1367.710 2.680 ;
        RECT 1368.830 2.400 1373.690 2.680 ;
        RECT 1374.810 2.400 1379.670 2.680 ;
        RECT 1380.790 2.400 1385.190 2.680 ;
        RECT 1386.310 2.400 1391.170 2.680 ;
        RECT 1392.290 2.400 1397.150 2.680 ;
        RECT 1398.270 2.400 1403.130 2.680 ;
        RECT 1404.250 2.400 1409.110 2.680 ;
        RECT 1410.230 2.400 1415.090 2.680 ;
        RECT 1416.210 2.400 1421.070 2.680 ;
        RECT 1422.190 2.400 1426.590 2.680 ;
        RECT 1427.710 2.400 1432.570 2.680 ;
        RECT 1433.690 2.400 1438.550 2.680 ;
        RECT 1439.670 2.400 1444.530 2.680 ;
        RECT 1445.650 2.400 1450.510 2.680 ;
        RECT 1451.630 2.400 1456.490 2.680 ;
        RECT 1457.610 2.400 1462.470 2.680 ;
        RECT 1463.590 2.400 1467.990 2.680 ;
        RECT 1469.110 2.400 1473.970 2.680 ;
        RECT 1475.090 2.400 1479.950 2.680 ;
        RECT 1481.070 2.400 1485.930 2.680 ;
        RECT 1487.050 2.400 1491.910 2.680 ;
        RECT 1493.030 2.400 1497.890 2.680 ;
        RECT 1499.010 2.400 1503.410 2.680 ;
        RECT 1504.530 2.400 1509.390 2.680 ;
        RECT 1510.510 2.400 1515.370 2.680 ;
        RECT 1516.490 2.400 1521.350 2.680 ;
        RECT 1522.470 2.400 1527.330 2.680 ;
        RECT 1528.450 2.400 1533.310 2.680 ;
        RECT 1534.430 2.400 1539.290 2.680 ;
        RECT 1540.410 2.400 1544.810 2.680 ;
        RECT 1545.930 2.400 1550.790 2.680 ;
        RECT 1551.910 2.400 1556.770 2.680 ;
        RECT 1557.890 2.400 1562.750 2.680 ;
        RECT 1563.870 2.400 1568.730 2.680 ;
        RECT 1569.850 2.400 1574.710 2.680 ;
        RECT 1575.830 2.400 1580.690 2.680 ;
        RECT 1581.810 2.400 1586.210 2.680 ;
        RECT 1587.330 2.400 1592.190 2.680 ;
        RECT 1593.310 2.400 1598.170 2.680 ;
        RECT 1599.290 2.400 1604.150 2.680 ;
        RECT 1605.270 2.400 1610.130 2.680 ;
        RECT 1611.250 2.400 1616.110 2.680 ;
        RECT 1617.230 2.400 1621.630 2.680 ;
        RECT 1622.750 2.400 1627.610 2.680 ;
        RECT 1628.730 2.400 1633.590 2.680 ;
        RECT 1634.710 2.400 1639.570 2.680 ;
        RECT 1640.690 2.400 1645.550 2.680 ;
        RECT 1646.670 2.400 1651.530 2.680 ;
        RECT 1652.650 2.400 1657.510 2.680 ;
        RECT 1658.630 2.400 1663.030 2.680 ;
        RECT 1664.150 2.400 1669.010 2.680 ;
        RECT 1670.130 2.400 1674.990 2.680 ;
        RECT 1676.110 2.400 1680.970 2.680 ;
        RECT 1682.090 2.400 1686.950 2.680 ;
        RECT 1688.070 2.400 1692.930 2.680 ;
        RECT 1694.050 2.400 1698.910 2.680 ;
        RECT 1700.030 2.400 1704.430 2.680 ;
        RECT 1705.550 2.400 1710.410 2.680 ;
        RECT 1711.530 2.400 1716.390 2.680 ;
        RECT 1717.510 2.400 1722.370 2.680 ;
        RECT 1723.490 2.400 1728.350 2.680 ;
        RECT 1729.470 2.400 1734.330 2.680 ;
        RECT 1735.450 2.400 1739.850 2.680 ;
        RECT 1740.970 2.400 1745.830 2.680 ;
        RECT 1746.950 2.400 1751.810 2.680 ;
        RECT 1752.930 2.400 1757.790 2.680 ;
        RECT 1758.910 2.400 1763.770 2.680 ;
        RECT 1764.890 2.400 1769.750 2.680 ;
        RECT 1770.870 2.400 1775.730 2.680 ;
        RECT 1776.850 2.400 1781.250 2.680 ;
        RECT 1782.370 2.400 1787.230 2.680 ;
        RECT 1788.350 2.400 1793.210 2.680 ;
        RECT 1794.330 2.400 1799.190 2.680 ;
        RECT 1800.310 2.400 1805.170 2.680 ;
        RECT 1806.290 2.400 1811.150 2.680 ;
        RECT 1812.270 2.400 1817.130 2.680 ;
        RECT 1818.250 2.400 1822.650 2.680 ;
        RECT 1823.770 2.400 1828.630 2.680 ;
        RECT 1829.750 2.400 1834.610 2.680 ;
        RECT 1835.730 2.400 1840.590 2.680 ;
        RECT 1841.710 2.400 1846.570 2.680 ;
        RECT 1847.690 2.400 1852.550 2.680 ;
        RECT 1853.670 2.400 1858.070 2.680 ;
        RECT 1859.190 2.400 1864.050 2.680 ;
        RECT 1865.170 2.400 1870.030 2.680 ;
        RECT 1871.150 2.400 1876.010 2.680 ;
        RECT 1877.130 2.400 1881.990 2.680 ;
        RECT 1883.110 2.400 1887.970 2.680 ;
        RECT 1889.090 2.400 1893.950 2.680 ;
        RECT 1895.070 2.400 1899.470 2.680 ;
        RECT 1900.590 2.400 1905.450 2.680 ;
        RECT 1906.570 2.400 1911.430 2.680 ;
        RECT 1912.550 2.400 1917.410 2.680 ;
        RECT 1918.530 2.400 1923.390 2.680 ;
        RECT 1924.510 2.400 1929.370 2.680 ;
        RECT 1930.490 2.400 1935.350 2.680 ;
        RECT 1936.470 2.400 1940.870 2.680 ;
        RECT 1941.990 2.400 1946.850 2.680 ;
        RECT 1947.970 2.400 1952.830 2.680 ;
        RECT 1953.950 2.400 1958.810 2.680 ;
        RECT 1959.930 2.400 1964.790 2.680 ;
        RECT 1965.910 2.400 1970.770 2.680 ;
        RECT 1971.890 2.400 1976.290 2.680 ;
        RECT 1977.410 2.400 1982.270 2.680 ;
        RECT 1983.390 2.400 1988.250 2.680 ;
        RECT 1989.370 2.400 1994.230 2.680 ;
        RECT 1995.350 2.400 2000.210 2.680 ;
        RECT 2001.330 2.400 2006.190 2.680 ;
        RECT 2007.310 2.400 2012.170 2.680 ;
        RECT 2013.290 2.400 2017.690 2.680 ;
        RECT 2018.810 2.400 2023.670 2.680 ;
        RECT 2024.790 2.400 2029.650 2.680 ;
        RECT 2030.770 2.400 2035.630 2.680 ;
        RECT 2036.750 2.400 2041.610 2.680 ;
        RECT 2042.730 2.400 2047.590 2.680 ;
        RECT 2048.710 2.400 2053.570 2.680 ;
        RECT 2054.690 2.400 2059.090 2.680 ;
        RECT 2060.210 2.400 2065.070 2.680 ;
        RECT 2066.190 2.400 2071.050 2.680 ;
        RECT 2072.170 2.400 2077.030 2.680 ;
        RECT 2078.150 2.400 2083.010 2.680 ;
        RECT 2084.130 2.400 2088.990 2.680 ;
        RECT 2090.110 2.400 2094.510 2.680 ;
        RECT 2095.630 2.400 2100.490 2.680 ;
        RECT 2101.610 2.400 2106.470 2.680 ;
        RECT 2107.590 2.400 2112.450 2.680 ;
        RECT 2113.570 2.400 2118.430 2.680 ;
        RECT 2119.550 2.400 2124.410 2.680 ;
        RECT 2125.530 2.400 2130.390 2.680 ;
        RECT 2131.510 2.400 2135.910 2.680 ;
        RECT 2137.030 2.400 2141.890 2.680 ;
        RECT 2143.010 2.400 2147.870 2.680 ;
        RECT 2148.990 2.400 2153.850 2.680 ;
        RECT 2154.970 2.400 2159.830 2.680 ;
        RECT 2160.950 2.400 2165.810 2.680 ;
        RECT 2166.930 2.400 2171.790 2.680 ;
        RECT 2172.910 2.400 2177.310 2.680 ;
        RECT 2178.430 2.400 2183.290 2.680 ;
        RECT 2184.410 2.400 2189.270 2.680 ;
        RECT 2190.390 2.400 2195.250 2.680 ;
        RECT 2196.370 2.400 2201.230 2.680 ;
        RECT 2202.350 2.400 2207.210 2.680 ;
        RECT 2208.330 2.400 2212.730 2.680 ;
        RECT 2213.850 2.400 2218.710 2.680 ;
        RECT 2219.830 2.400 2224.690 2.680 ;
        RECT 2225.810 2.400 2230.670 2.680 ;
        RECT 2231.790 2.400 2236.650 2.680 ;
        RECT 2237.770 2.400 2242.630 2.680 ;
        RECT 2243.750 2.400 2248.610 2.680 ;
        RECT 2249.730 2.400 2254.130 2.680 ;
        RECT 2255.250 2.400 2260.110 2.680 ;
        RECT 2261.230 2.400 2266.090 2.680 ;
        RECT 2267.210 2.400 2272.070 2.680 ;
        RECT 2273.190 2.400 2278.050 2.680 ;
        RECT 2279.170 2.400 2284.030 2.680 ;
        RECT 2285.150 2.400 2290.010 2.680 ;
        RECT 2291.130 2.400 2295.530 2.680 ;
        RECT 2296.650 2.400 2301.510 2.680 ;
        RECT 2302.630 2.400 2307.490 2.680 ;
        RECT 2308.610 2.400 2313.470 2.680 ;
        RECT 2314.590 2.400 2319.450 2.680 ;
        RECT 2320.570 2.400 2325.430 2.680 ;
        RECT 2326.550 2.400 2330.950 2.680 ;
        RECT 2332.070 2.400 2336.930 2.680 ;
        RECT 2338.050 2.400 2342.910 2.680 ;
        RECT 2344.030 2.400 2348.890 2.680 ;
        RECT 2350.010 2.400 2354.870 2.680 ;
        RECT 2355.990 2.400 2360.850 2.680 ;
        RECT 2361.970 2.400 2366.830 2.680 ;
        RECT 2367.950 2.400 2372.350 2.680 ;
        RECT 2373.470 2.400 2378.330 2.680 ;
        RECT 2379.450 2.400 2384.310 2.680 ;
        RECT 2385.430 2.400 2390.290 2.680 ;
        RECT 2391.410 2.400 2396.270 2.680 ;
        RECT 2397.390 2.400 2402.250 2.680 ;
        RECT 2403.370 2.400 2408.230 2.680 ;
        RECT 2409.350 2.400 2413.750 2.680 ;
        RECT 2414.870 2.400 2419.730 2.680 ;
        RECT 2420.850 2.400 2425.710 2.680 ;
        RECT 2426.830 2.400 2431.690 2.680 ;
        RECT 2432.810 2.400 2437.670 2.680 ;
        RECT 2438.790 2.400 2443.650 2.680 ;
        RECT 2444.770 2.400 2449.170 2.680 ;
        RECT 2450.290 2.400 2455.150 2.680 ;
        RECT 2456.270 2.400 2461.130 2.680 ;
        RECT 2462.250 2.400 2467.110 2.680 ;
        RECT 2468.230 2.400 2473.090 2.680 ;
        RECT 2474.210 2.400 2479.070 2.680 ;
        RECT 2480.190 2.400 2485.050 2.680 ;
        RECT 2486.170 2.400 2490.570 2.680 ;
        RECT 2491.690 2.400 2496.550 2.680 ;
        RECT 2497.670 2.400 2502.530 2.680 ;
        RECT 2503.650 2.400 2508.510 2.680 ;
        RECT 2509.630 2.400 2514.490 2.680 ;
        RECT 2515.610 2.400 2520.470 2.680 ;
        RECT 2521.590 2.400 2526.450 2.680 ;
        RECT 2527.570 2.400 2531.970 2.680 ;
        RECT 2533.090 2.400 2537.950 2.680 ;
        RECT 2539.070 2.400 2543.930 2.680 ;
        RECT 2545.050 2.400 2549.910 2.680 ;
        RECT 2551.030 2.400 2555.890 2.680 ;
        RECT 2557.010 2.400 2561.870 2.680 ;
        RECT 2562.990 2.400 2567.390 2.680 ;
        RECT 2568.510 2.400 2573.370 2.680 ;
        RECT 2574.490 2.400 2579.350 2.680 ;
        RECT 2580.470 2.400 2585.330 2.680 ;
        RECT 2586.450 2.400 2591.310 2.680 ;
        RECT 2592.430 2.400 2597.290 2.680 ;
        RECT 2598.410 2.400 2603.270 2.680 ;
        RECT 2604.390 2.400 2608.790 2.680 ;
        RECT 2609.910 2.400 2614.770 2.680 ;
        RECT 2615.890 2.400 2620.750 2.680 ;
        RECT 2621.870 2.400 2626.730 2.680 ;
        RECT 2627.850 2.400 2632.710 2.680 ;
        RECT 2633.830 2.400 2638.690 2.680 ;
        RECT 2639.810 2.400 2644.670 2.680 ;
        RECT 2645.790 2.400 2650.190 2.680 ;
        RECT 2651.310 2.400 2656.170 2.680 ;
        RECT 2657.290 2.400 2662.150 2.680 ;
        RECT 2663.270 2.400 2668.130 2.680 ;
        RECT 2669.250 2.400 2674.110 2.680 ;
        RECT 2675.230 2.400 2680.090 2.680 ;
        RECT 2681.210 2.400 2685.610 2.680 ;
        RECT 2686.730 2.400 2691.590 2.680 ;
        RECT 2692.710 2.400 2697.570 2.680 ;
        RECT 2698.690 2.400 2703.550 2.680 ;
        RECT 2704.670 2.400 2709.530 2.680 ;
        RECT 2710.650 2.400 2715.510 2.680 ;
        RECT 2716.630 2.400 2721.490 2.680 ;
        RECT 2722.610 2.400 2727.010 2.680 ;
        RECT 2728.130 2.400 2732.990 2.680 ;
        RECT 2734.110 2.400 2738.970 2.680 ;
        RECT 2740.090 2.400 2744.950 2.680 ;
        RECT 2746.070 2.400 2750.930 2.680 ;
        RECT 2752.050 2.400 2756.910 2.680 ;
        RECT 2758.030 2.400 2762.890 2.680 ;
        RECT 2764.010 2.400 2768.410 2.680 ;
        RECT 2769.530 2.400 2774.390 2.680 ;
        RECT 2775.510 2.400 2780.370 2.680 ;
        RECT 2781.490 2.400 2786.350 2.680 ;
        RECT 2787.470 2.400 2792.330 2.680 ;
        RECT 2793.450 2.400 2798.310 2.680 ;
        RECT 2799.430 2.400 2803.830 2.680 ;
        RECT 2804.950 2.400 2809.810 2.680 ;
        RECT 2810.930 2.400 2815.790 2.680 ;
        RECT 2816.910 2.400 2821.770 2.680 ;
        RECT 2822.890 2.400 2827.750 2.680 ;
        RECT 2828.870 2.400 2833.730 2.680 ;
        RECT 2834.850 2.400 2839.710 2.680 ;
        RECT 2840.830 2.400 2845.230 2.680 ;
        RECT 2846.350 2.400 2851.210 2.680 ;
        RECT 2852.330 2.400 2857.190 2.680 ;
        RECT 2858.310 2.400 2863.170 2.680 ;
        RECT 2864.290 2.400 2869.150 2.680 ;
        RECT 2870.270 2.400 2875.130 2.680 ;
        RECT 2876.250 2.400 2881.110 2.680 ;
        RECT 2882.230 2.400 2886.630 2.680 ;
        RECT 2887.750 2.400 2892.610 2.680 ;
        RECT 2893.730 2.400 2898.590 2.680 ;
        RECT 2899.710 2.400 2903.890 2.680 ;
      LAYER met3 ;
        RECT 2.825 3487.020 2917.600 3502.505 ;
        RECT 2.825 3485.020 2917.200 3487.020 ;
        RECT 2.825 3420.380 2917.600 3485.020 ;
        RECT 2.825 3418.380 2917.200 3420.380 ;
        RECT 2.825 3354.420 2917.600 3418.380 ;
        RECT 2.825 3352.420 2917.200 3354.420 ;
        RECT 2.825 3287.780 2917.600 3352.420 ;
        RECT 2.825 3285.780 2917.200 3287.780 ;
        RECT 2.825 3221.140 2917.600 3285.780 ;
        RECT 2.825 3219.140 2917.200 3221.140 ;
        RECT 2.825 3155.180 2917.600 3219.140 ;
        RECT 2.825 3153.180 2917.200 3155.180 ;
        RECT 2.825 3088.540 2917.600 3153.180 ;
        RECT 2.825 3086.540 2917.200 3088.540 ;
        RECT 2.825 3021.900 2917.600 3086.540 ;
        RECT 2.825 3019.900 2917.200 3021.900 ;
        RECT 2.825 2955.940 2917.600 3019.900 ;
        RECT 2.825 2953.940 2917.200 2955.940 ;
        RECT 2.825 2889.300 2917.600 2953.940 ;
        RECT 2.825 2887.300 2917.200 2889.300 ;
        RECT 2.825 2822.660 2917.600 2887.300 ;
        RECT 2.825 2820.660 2917.200 2822.660 ;
        RECT 2.825 2756.700 2917.600 2820.660 ;
        RECT 2.825 2754.700 2917.200 2756.700 ;
        RECT 2.825 2690.060 2917.600 2754.700 ;
        RECT 2.825 2688.060 2917.200 2690.060 ;
        RECT 2.825 2623.420 2917.600 2688.060 ;
        RECT 2.825 2621.420 2917.200 2623.420 ;
        RECT 2.825 2557.460 2917.600 2621.420 ;
        RECT 2.825 2555.460 2917.200 2557.460 ;
        RECT 2.825 2490.820 2917.600 2555.460 ;
        RECT 2.825 2488.820 2917.200 2490.820 ;
        RECT 2.825 2424.180 2917.600 2488.820 ;
        RECT 2.825 2422.180 2917.200 2424.180 ;
        RECT 2.825 2358.220 2917.600 2422.180 ;
        RECT 2.825 2356.220 2917.200 2358.220 ;
        RECT 2.825 2291.580 2917.600 2356.220 ;
        RECT 2.825 2289.580 2917.200 2291.580 ;
        RECT 2.825 2224.940 2917.600 2289.580 ;
        RECT 2.825 2222.940 2917.200 2224.940 ;
        RECT 2.825 2158.980 2917.600 2222.940 ;
        RECT 2.825 2156.980 2917.200 2158.980 ;
        RECT 2.825 2092.340 2917.600 2156.980 ;
        RECT 2.825 2090.340 2917.200 2092.340 ;
        RECT 2.825 2025.700 2917.600 2090.340 ;
        RECT 2.825 2023.700 2917.200 2025.700 ;
        RECT 2.825 1959.740 2917.600 2023.700 ;
        RECT 2.825 1957.740 2917.200 1959.740 ;
        RECT 2.825 1893.100 2917.600 1957.740 ;
        RECT 2.825 1891.100 2917.200 1893.100 ;
        RECT 2.825 1826.460 2917.600 1891.100 ;
        RECT 2.825 1824.460 2917.200 1826.460 ;
        RECT 2.825 1760.500 2917.600 1824.460 ;
        RECT 2.825 1758.500 2917.200 1760.500 ;
        RECT 2.825 1693.860 2917.600 1758.500 ;
        RECT 2.825 1691.860 2917.200 1693.860 ;
        RECT 2.825 1627.220 2917.600 1691.860 ;
        RECT 2.825 1625.220 2917.200 1627.220 ;
        RECT 2.825 1561.260 2917.600 1625.220 ;
        RECT 2.825 1559.260 2917.200 1561.260 ;
        RECT 2.825 1494.620 2917.600 1559.260 ;
        RECT 2.825 1492.620 2917.200 1494.620 ;
        RECT 2.825 1427.980 2917.600 1492.620 ;
        RECT 2.825 1425.980 2917.200 1427.980 ;
        RECT 2.825 1362.020 2917.600 1425.980 ;
        RECT 2.825 1360.020 2917.200 1362.020 ;
        RECT 2.825 1295.380 2917.600 1360.020 ;
        RECT 2.825 1293.380 2917.200 1295.380 ;
        RECT 2.825 1228.740 2917.600 1293.380 ;
        RECT 2.825 1226.740 2917.200 1228.740 ;
        RECT 2.825 1162.780 2917.600 1226.740 ;
        RECT 2.825 1160.780 2917.200 1162.780 ;
        RECT 2.825 1096.140 2917.600 1160.780 ;
        RECT 2.825 1094.140 2917.200 1096.140 ;
        RECT 2.825 1029.500 2917.600 1094.140 ;
        RECT 2.825 1027.500 2917.200 1029.500 ;
        RECT 2.825 963.540 2917.600 1027.500 ;
        RECT 2.825 961.540 2917.200 963.540 ;
        RECT 2.825 896.900 2917.600 961.540 ;
        RECT 2.825 894.900 2917.200 896.900 ;
        RECT 2.825 830.260 2917.600 894.900 ;
        RECT 2.825 828.260 2917.200 830.260 ;
        RECT 2.825 764.300 2917.600 828.260 ;
        RECT 2.825 762.300 2917.200 764.300 ;
        RECT 2.825 697.660 2917.600 762.300 ;
        RECT 2.825 695.660 2917.200 697.660 ;
        RECT 2.825 631.020 2917.600 695.660 ;
        RECT 2.825 629.020 2917.200 631.020 ;
        RECT 2.825 565.060 2917.600 629.020 ;
        RECT 2.825 563.060 2917.200 565.060 ;
        RECT 2.825 498.420 2917.600 563.060 ;
        RECT 2.825 496.420 2917.200 498.420 ;
        RECT 2.825 431.780 2917.600 496.420 ;
        RECT 2.825 429.780 2917.200 431.780 ;
        RECT 2.825 365.820 2917.600 429.780 ;
        RECT 2.825 363.820 2917.200 365.820 ;
        RECT 2.825 299.180 2917.600 363.820 ;
        RECT 2.825 297.180 2917.200 299.180 ;
        RECT 2.825 232.540 2917.600 297.180 ;
        RECT 2.825 230.540 2917.200 232.540 ;
        RECT 2.825 166.580 2917.600 230.540 ;
        RECT 2.825 164.580 2917.200 166.580 ;
        RECT 2.825 99.940 2917.600 164.580 ;
        RECT 2.825 97.940 2917.200 99.940 ;
        RECT 2.825 33.980 2917.600 97.940 ;
        RECT 2.825 31.980 2917.200 33.980 ;
        RECT 2.825 3.575 2917.600 31.980 ;
      LAYER met4 ;
        RECT 43.535 4.935 45.770 2821.825 ;
        RECT 49.670 4.935 64.370 2821.825 ;
        RECT 68.270 4.935 82.970 2821.825 ;
        RECT 86.870 4.935 101.570 2821.825 ;
        RECT 105.470 4.935 120.170 2821.825 ;
        RECT 124.070 4.935 138.770 2821.825 ;
        RECT 142.670 4.935 188.570 2821.825 ;
        RECT 192.470 4.935 207.170 2821.825 ;
        RECT 211.070 4.935 225.770 2821.825 ;
        RECT 229.670 4.935 244.370 2821.825 ;
        RECT 248.270 4.935 262.970 2821.825 ;
        RECT 266.870 4.935 281.570 2821.825 ;
        RECT 285.470 4.935 300.170 2821.825 ;
        RECT 304.070 4.935 318.770 2821.825 ;
        RECT 322.670 4.935 368.570 2821.825 ;
        RECT 372.470 362.820 387.170 2821.825 ;
        RECT 391.070 362.820 405.770 2821.825 ;
        RECT 372.470 4.935 405.770 362.820 ;
        RECT 409.670 4.935 424.370 2821.825 ;
        RECT 428.270 4.935 442.970 2821.825 ;
        RECT 446.870 4.935 461.570 2821.825 ;
        RECT 465.470 4.935 480.170 2821.825 ;
        RECT 484.070 4.935 498.770 2821.825 ;
        RECT 502.670 4.935 548.570 2821.825 ;
        RECT 552.470 4.935 567.170 2821.825 ;
        RECT 571.070 4.935 585.770 2821.825 ;
        RECT 589.670 4.935 604.370 2821.825 ;
        RECT 608.270 4.935 622.970 2821.825 ;
        RECT 626.870 4.935 641.570 2821.825 ;
        RECT 645.470 4.935 660.170 2821.825 ;
        RECT 664.070 4.935 678.770 2821.825 ;
        RECT 682.670 4.935 728.570 2821.825 ;
        RECT 732.470 4.935 747.170 2821.825 ;
        RECT 751.070 4.935 765.770 2821.825 ;
        RECT 769.670 4.935 784.370 2821.825 ;
        RECT 788.270 4.935 802.970 2821.825 ;
        RECT 806.870 4.935 821.570 2821.825 ;
        RECT 825.470 4.935 840.170 2821.825 ;
        RECT 844.070 4.935 858.770 2821.825 ;
        RECT 862.670 4.935 908.570 2821.825 ;
        RECT 912.470 4.935 927.170 2821.825 ;
        RECT 931.070 4.935 945.770 2821.825 ;
        RECT 949.670 4.935 964.370 2821.825 ;
        RECT 968.270 4.935 982.970 2821.825 ;
        RECT 986.870 4.935 1001.570 2821.825 ;
        RECT 1005.470 4.935 1020.170 2821.825 ;
        RECT 1024.070 4.935 1038.770 2821.825 ;
        RECT 1042.670 4.935 1088.570 2821.825 ;
        RECT 1092.470 4.935 1107.170 2821.825 ;
        RECT 1111.070 4.935 1125.770 2821.825 ;
        RECT 1129.670 4.935 1144.370 2821.825 ;
        RECT 1148.270 4.935 1162.970 2821.825 ;
        RECT 1166.870 4.935 1181.570 2821.825 ;
        RECT 1185.470 4.935 1200.170 2821.825 ;
        RECT 1204.070 4.935 1218.770 2821.825 ;
        RECT 1222.670 4.935 1268.570 2821.825 ;
        RECT 1272.470 4.935 1287.170 2821.825 ;
        RECT 1291.070 4.935 1305.770 2821.825 ;
        RECT 1309.670 4.935 1324.370 2821.825 ;
        RECT 1328.270 4.935 1342.970 2821.825 ;
        RECT 1346.870 4.935 1361.570 2821.825 ;
        RECT 1365.470 4.935 1380.170 2821.825 ;
        RECT 1384.070 4.935 1398.770 2821.825 ;
        RECT 1402.670 4.935 1448.570 2821.825 ;
        RECT 1452.470 4.935 1467.170 2821.825 ;
        RECT 1471.070 4.935 1485.770 2821.825 ;
        RECT 1489.670 4.935 1504.370 2821.825 ;
        RECT 1508.270 4.935 1522.970 2821.825 ;
        RECT 1526.870 4.935 1541.570 2821.825 ;
        RECT 1545.470 4.935 1560.170 2821.825 ;
        RECT 1564.070 4.935 1578.770 2821.825 ;
        RECT 1582.670 4.935 1628.570 2821.825 ;
        RECT 1632.470 4.935 1647.170 2821.825 ;
        RECT 1651.070 4.935 1665.770 2821.825 ;
        RECT 1669.670 4.935 1684.370 2821.825 ;
        RECT 1688.270 4.935 1702.970 2821.825 ;
        RECT 1706.870 4.935 1721.570 2821.825 ;
        RECT 1725.470 4.935 1740.170 2821.825 ;
        RECT 1744.070 4.935 1758.770 2821.825 ;
        RECT 1762.670 4.935 1808.570 2821.825 ;
        RECT 1812.470 4.935 1827.170 2821.825 ;
        RECT 1831.070 4.935 1845.770 2821.825 ;
        RECT 1849.670 4.935 1864.370 2821.825 ;
        RECT 1868.270 4.935 1882.970 2821.825 ;
        RECT 1886.870 4.935 1901.570 2821.825 ;
        RECT 1905.470 4.935 1920.170 2821.825 ;
        RECT 1924.070 4.935 1938.770 2821.825 ;
        RECT 1942.670 4.935 1988.570 2821.825 ;
        RECT 1992.470 4.935 2007.170 2821.825 ;
        RECT 2011.070 4.935 2025.770 2821.825 ;
        RECT 2029.670 4.935 2044.370 2821.825 ;
        RECT 2048.270 4.935 2062.970 2821.825 ;
        RECT 2066.870 4.935 2081.570 2821.825 ;
        RECT 2085.470 4.935 2100.170 2821.825 ;
        RECT 2104.070 4.935 2118.770 2821.825 ;
        RECT 2122.670 4.935 2168.570 2821.825 ;
        RECT 2172.470 4.935 2187.170 2821.825 ;
        RECT 2191.070 4.935 2205.770 2821.825 ;
        RECT 2209.670 4.935 2224.370 2821.825 ;
        RECT 2228.270 4.935 2242.970 2821.825 ;
        RECT 2246.870 4.935 2261.570 2821.825 ;
        RECT 2265.470 4.935 2280.170 2821.825 ;
        RECT 2284.070 4.935 2298.770 2821.825 ;
        RECT 2302.670 4.935 2348.570 2821.825 ;
        RECT 2352.470 4.935 2367.170 2821.825 ;
        RECT 2371.070 4.935 2385.770 2821.825 ;
        RECT 2389.670 4.935 2404.370 2821.825 ;
        RECT 2408.270 4.935 2422.970 2821.825 ;
        RECT 2426.870 4.935 2441.570 2821.825 ;
        RECT 2445.470 4.935 2460.170 2821.825 ;
        RECT 2464.070 4.935 2478.770 2821.825 ;
        RECT 2482.670 4.935 2528.570 2821.825 ;
        RECT 2532.470 4.935 2547.170 2821.825 ;
        RECT 2551.070 4.935 2565.770 2821.825 ;
        RECT 2569.670 4.935 2584.370 2821.825 ;
        RECT 2588.270 4.935 2602.970 2821.825 ;
        RECT 2606.870 4.935 2621.570 2821.825 ;
        RECT 2625.470 4.935 2640.170 2821.825 ;
        RECT 2644.070 4.935 2658.770 2821.825 ;
        RECT 2662.670 4.935 2708.570 2821.825 ;
        RECT 2712.470 4.935 2727.170 2821.825 ;
        RECT 2731.070 4.935 2745.770 2821.825 ;
        RECT 2749.670 4.935 2764.370 2821.825 ;
        RECT 2768.270 4.935 2782.970 2821.825 ;
        RECT 2786.870 4.935 2801.570 2821.825 ;
        RECT 2805.470 4.935 2820.170 2821.825 ;
        RECT 2824.070 4.935 2838.770 2821.825 ;
        RECT 2842.670 4.935 2888.570 2821.825 ;
        RECT 2892.470 4.935 2902.305 2821.825 ;
  END
END user_project_wrapper
END LIBRARY

