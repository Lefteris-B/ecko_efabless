magic
tech sky130A
magscale 1 2
timestamp 1715852960
<< viali >>
rect 20913 27081 20947 27115
rect 16773 27013 16807 27047
rect 21833 27013 21867 27047
rect 3985 26945 4019 26979
rect 11069 26945 11103 26979
rect 14933 26945 14967 26979
rect 16681 26945 16715 26979
rect 16957 26945 16991 26979
rect 20821 26945 20855 26979
rect 21189 26945 21223 26979
rect 21281 26945 21315 26979
rect 1409 26877 1443 26911
rect 21005 26877 21039 26911
rect 21557 26877 21591 26911
rect 22385 26877 22419 26911
rect 21189 26809 21223 26843
rect 21373 26809 21407 26843
rect 16957 26741 16991 26775
rect 21465 26741 21499 26775
rect 16497 26537 16531 26571
rect 16681 26537 16715 26571
rect 17509 26537 17543 26571
rect 20729 26537 20763 26571
rect 22661 26537 22695 26571
rect 15853 26401 15887 26435
rect 17417 26401 17451 26435
rect 22477 26401 22511 26435
rect 9505 26333 9539 26367
rect 11437 26333 11471 26367
rect 12541 26333 12575 26367
rect 12725 26333 12759 26367
rect 15934 26333 15968 26367
rect 16037 26333 16071 26367
rect 16129 26333 16163 26367
rect 16773 26333 16807 26367
rect 18061 26333 18095 26367
rect 19441 26333 19475 26367
rect 19717 26333 19751 26367
rect 19901 26333 19935 26367
rect 19993 26333 20027 26367
rect 20545 26333 20579 26367
rect 21281 26333 21315 26367
rect 22385 26333 22419 26367
rect 22753 26333 22787 26367
rect 16313 26265 16347 26299
rect 16513 26265 16547 26299
rect 9321 26197 9355 26231
rect 10793 26197 10827 26231
rect 12633 26197 12667 26231
rect 15669 26197 15703 26231
rect 19257 26197 19291 26231
rect 21741 26197 21775 26231
rect 22477 26197 22511 26231
rect 16681 25993 16715 26027
rect 20637 25993 20671 26027
rect 21833 25993 21867 26027
rect 12449 25925 12483 25959
rect 12909 25925 12943 25959
rect 13553 25925 13587 25959
rect 15577 25925 15611 25959
rect 18880 25925 18914 25959
rect 20253 25925 20287 25959
rect 20453 25925 20487 25959
rect 20821 25925 20855 25959
rect 8217 25857 8251 25891
rect 8484 25857 8518 25891
rect 9689 25857 9723 25891
rect 9956 25857 9990 25891
rect 11345 25857 11379 25891
rect 11621 25857 11655 25891
rect 12357 25857 12391 25891
rect 12541 25857 12575 25891
rect 12679 25857 12713 25891
rect 13093 25857 13127 25891
rect 13277 25857 13311 25891
rect 13366 25857 13400 25891
rect 13461 25857 13495 25891
rect 13737 25857 13771 25891
rect 13829 25857 13863 25891
rect 14657 25857 14691 25891
rect 15117 25857 15151 25891
rect 16221 25857 16255 25891
rect 17794 25857 17828 25891
rect 20545 25857 20579 25891
rect 21097 25857 21131 25891
rect 21189 25857 21223 25891
rect 21281 25857 21315 25891
rect 21465 25857 21499 25891
rect 22946 25857 22980 25891
rect 23213 25857 23247 25891
rect 12817 25789 12851 25823
rect 14381 25789 14415 25823
rect 14473 25789 14507 25823
rect 15301 25789 15335 25823
rect 18061 25789 18095 25823
rect 18613 25789 18647 25823
rect 20913 25789 20947 25823
rect 11069 25721 11103 25755
rect 12081 25721 12115 25755
rect 15669 25721 15703 25755
rect 20085 25721 20119 25755
rect 9597 25653 9631 25687
rect 11161 25653 11195 25687
rect 11805 25653 11839 25687
rect 12173 25653 12207 25687
rect 13645 25653 13679 25687
rect 13921 25653 13955 25687
rect 14841 25653 14875 25687
rect 14933 25653 14967 25687
rect 15485 25653 15519 25687
rect 19993 25653 20027 25687
rect 20269 25653 20303 25687
rect 20821 25653 20855 25687
rect 9505 25449 9539 25483
rect 9689 25449 9723 25483
rect 9965 25449 9999 25483
rect 13737 25449 13771 25483
rect 14105 25449 14139 25483
rect 16221 25449 16255 25483
rect 17877 25449 17911 25483
rect 18981 25449 19015 25483
rect 22753 25449 22787 25483
rect 16497 25313 16531 25347
rect 18429 25313 18463 25347
rect 19073 25313 19107 25347
rect 10152 25223 10186 25257
rect 10241 25245 10275 25279
rect 10425 25245 10459 25279
rect 10517 25245 10551 25279
rect 10609 25245 10643 25279
rect 12081 25245 12115 25279
rect 12348 25245 12382 25279
rect 14289 25245 14323 25279
rect 14381 25245 14415 25279
rect 14473 25245 14507 25279
rect 14657 25245 14691 25279
rect 14749 25245 14783 25279
rect 16221 25245 16255 25279
rect 16405 25245 16439 25279
rect 16764 25245 16798 25279
rect 17969 25245 18003 25279
rect 18153 25245 18187 25279
rect 18337 25245 18371 25279
rect 18521 25245 18555 25279
rect 18827 25245 18861 25279
rect 19257 25245 19291 25279
rect 20913 25245 20947 25279
rect 21097 25245 21131 25279
rect 21373 25245 21407 25279
rect 9873 25177 9907 25211
rect 10876 25177 10910 25211
rect 13553 25177 13587 25211
rect 13769 25177 13803 25211
rect 14994 25177 15028 25211
rect 19524 25177 19558 25211
rect 21618 25177 21652 25211
rect 9673 25109 9707 25143
rect 11989 25109 12023 25143
rect 13461 25109 13495 25143
rect 13921 25109 13955 25143
rect 16129 25109 16163 25143
rect 18061 25109 18095 25143
rect 18613 25109 18647 25143
rect 20637 25109 20671 25143
rect 20729 25109 20763 25143
rect 10609 24905 10643 24939
rect 11345 24905 11379 24939
rect 13921 24905 13955 24939
rect 15761 24905 15795 24939
rect 15945 24905 15979 24939
rect 16129 24905 16163 24939
rect 17141 24905 17175 24939
rect 19809 24905 19843 24939
rect 21991 24905 22025 24939
rect 9781 24837 9815 24871
rect 11897 24837 11931 24871
rect 13093 24837 13127 24871
rect 16313 24837 16347 24871
rect 17233 24837 17267 24871
rect 18604 24837 18638 24871
rect 21281 24837 21315 24871
rect 22201 24837 22235 24871
rect 21511 24803 21545 24837
rect 9137 24769 9171 24803
rect 9597 24769 9631 24803
rect 10333 24769 10367 24803
rect 10609 24769 10643 24803
rect 10793 24769 10827 24803
rect 11161 24769 11195 24803
rect 12265 24769 12299 24803
rect 13829 24769 13863 24803
rect 14013 24769 14047 24803
rect 14648 24769 14682 24803
rect 16221 24769 16255 24803
rect 16681 24769 16715 24803
rect 16957 24769 16991 24803
rect 17509 24769 17543 24803
rect 20453 24769 20487 24803
rect 22385 24769 22419 24803
rect 9229 24701 9263 24735
rect 10517 24701 10551 24735
rect 10977 24701 11011 24735
rect 12081 24701 12115 24735
rect 12173 24701 12207 24735
rect 12449 24701 12483 24735
rect 12633 24701 12667 24735
rect 12725 24701 12759 24735
rect 12817 24701 12851 24735
rect 12909 24701 12943 24735
rect 13645 24701 13679 24735
rect 14381 24701 14415 24735
rect 16497 24701 16531 24735
rect 17233 24701 17267 24735
rect 18337 24701 18371 24735
rect 21097 24701 21131 24735
rect 9505 24633 9539 24667
rect 17417 24633 17451 24667
rect 19717 24633 19751 24667
rect 21833 24633 21867 24667
rect 22569 24633 22603 24667
rect 9965 24565 9999 24599
rect 10149 24565 10183 24599
rect 16773 24565 16807 24599
rect 20545 24565 20579 24599
rect 21465 24565 21499 24599
rect 21649 24565 21683 24599
rect 22017 24565 22051 24599
rect 9321 24361 9355 24395
rect 10057 24361 10091 24395
rect 12909 24361 12943 24395
rect 14657 24361 14691 24395
rect 16129 24361 16163 24395
rect 19073 24361 19107 24395
rect 19809 24361 19843 24395
rect 8769 24293 8803 24327
rect 12173 24293 12207 24327
rect 10425 24225 10459 24259
rect 11805 24225 11839 24259
rect 15761 24225 15795 24259
rect 19441 24225 19475 24259
rect 23213 24225 23247 24259
rect 7389 24157 7423 24191
rect 9873 24157 9907 24191
rect 10241 24157 10275 24191
rect 10517 24157 10551 24191
rect 12633 24157 12667 24191
rect 12909 24157 12943 24191
rect 14841 24157 14875 24191
rect 15945 24157 15979 24191
rect 18889 24157 18923 24191
rect 19073 24157 19107 24191
rect 19625 24157 19659 24191
rect 19717 24157 19751 24191
rect 19993 24157 20027 24191
rect 20085 24157 20119 24191
rect 20177 24157 20211 24191
rect 20269 24157 20303 24191
rect 23121 24157 23155 24191
rect 23305 24157 23339 24191
rect 23397 24157 23431 24191
rect 26157 24157 26191 24191
rect 7656 24089 7690 24123
rect 12725 24089 12759 24123
rect 19441 24089 19475 24123
rect 12265 24021 12299 24055
rect 22937 24021 22971 24055
rect 7757 23817 7791 23851
rect 9505 23817 9539 23851
rect 9689 23817 9723 23851
rect 22109 23817 22143 23851
rect 24133 23817 24167 23851
rect 7941 23681 7975 23715
rect 8033 23681 8067 23715
rect 8300 23681 8334 23715
rect 10149 23681 10183 23715
rect 10333 23681 10367 23715
rect 14473 23681 14507 23715
rect 22017 23681 22051 23715
rect 22201 23681 22235 23715
rect 22293 23681 22327 23715
rect 22385 23681 22419 23715
rect 22569 23681 22603 23715
rect 23009 23681 23043 23715
rect 24777 23681 24811 23715
rect 10241 23613 10275 23647
rect 14841 23613 14875 23647
rect 15393 23613 15427 23647
rect 19717 23613 19751 23647
rect 22753 23613 22787 23647
rect 10057 23545 10091 23579
rect 22569 23545 22603 23579
rect 9413 23477 9447 23511
rect 9689 23477 9723 23511
rect 14657 23477 14691 23511
rect 19073 23477 19107 23511
rect 24225 23477 24259 23511
rect 10149 23273 10183 23307
rect 10333 23273 10367 23307
rect 11345 23273 11379 23307
rect 13645 23273 13679 23307
rect 14473 23273 14507 23307
rect 16957 23273 16991 23307
rect 20821 23273 20855 23307
rect 11161 23205 11195 23239
rect 13737 23205 13771 23239
rect 17969 23205 18003 23239
rect 18245 23205 18279 23239
rect 9321 23137 9355 23171
rect 9413 23137 9447 23171
rect 10425 23137 10459 23171
rect 10977 23137 11011 23171
rect 13829 23137 13863 23171
rect 18613 23137 18647 23171
rect 19809 23137 19843 23171
rect 20269 23137 20303 23171
rect 21005 23137 21039 23171
rect 24777 23137 24811 23171
rect 9229 23069 9263 23103
rect 9505 23069 9539 23103
rect 9781 23069 9815 23103
rect 10701 23069 10735 23103
rect 11713 23069 11747 23103
rect 12173 23069 12207 23103
rect 12449 23069 12483 23103
rect 12633 23069 12667 23103
rect 12817 23069 12851 23103
rect 13369 23069 13403 23103
rect 13553 23069 13587 23103
rect 14197 23069 14231 23103
rect 14841 23069 14875 23103
rect 14933 23069 14967 23103
rect 15577 23069 15611 23103
rect 15945 23069 15979 23103
rect 17417 23069 17451 23103
rect 17785 23069 17819 23103
rect 17969 23069 18003 23103
rect 18153 23069 18187 23103
rect 18337 23069 18371 23103
rect 18429 23069 18463 23103
rect 20361 23069 20395 23103
rect 21649 23069 21683 23103
rect 21742 23069 21776 23103
rect 22114 23069 22148 23103
rect 22385 23069 22419 23103
rect 22569 23069 22603 23103
rect 22661 23069 22695 23103
rect 24593 23069 24627 23103
rect 24685 23069 24719 23103
rect 24869 23069 24903 23103
rect 25329 23069 25363 23103
rect 10149 23001 10183 23035
rect 10793 23001 10827 23035
rect 11345 23001 11379 23035
rect 17141 23001 17175 23035
rect 21557 23001 21591 23035
rect 21925 23001 21959 23035
rect 22017 23001 22051 23035
rect 22928 23001 22962 23035
rect 9689 22933 9723 22967
rect 10609 22933 10643 22967
rect 11989 22933 12023 22967
rect 15025 22933 15059 22967
rect 16589 22933 16623 22967
rect 16773 22933 16807 22967
rect 16941 22933 16975 22967
rect 17509 22933 17543 22967
rect 19257 22933 19291 22967
rect 20453 22933 20487 22967
rect 22293 22933 22327 22967
rect 22477 22933 22511 22967
rect 24041 22933 24075 22967
rect 24409 22933 24443 22967
rect 25145 22933 25179 22967
rect 9965 22729 9999 22763
rect 11345 22729 11379 22763
rect 13093 22729 13127 22763
rect 15117 22729 15151 22763
rect 15209 22729 15243 22763
rect 15853 22729 15887 22763
rect 16497 22729 16531 22763
rect 21097 22729 21131 22763
rect 23305 22729 23339 22763
rect 23581 22729 23615 22763
rect 23673 22729 23707 22763
rect 24317 22729 24351 22763
rect 25973 22729 26007 22763
rect 10701 22661 10735 22695
rect 11888 22661 11922 22695
rect 17018 22661 17052 22695
rect 23055 22661 23089 22695
rect 23857 22661 23891 22695
rect 8585 22593 8619 22627
rect 8852 22593 8886 22627
rect 10241 22593 10275 22627
rect 10425 22593 10459 22627
rect 11161 22593 11195 22627
rect 11621 22593 11655 22627
rect 13277 22593 13311 22627
rect 13369 22593 13403 22627
rect 13553 22593 13587 22627
rect 13645 22593 13679 22627
rect 14004 22593 14038 22627
rect 15485 22593 15519 22627
rect 15945 22593 15979 22627
rect 16313 22593 16347 22627
rect 18245 22593 18279 22627
rect 18512 22593 18546 22627
rect 19717 22593 19751 22627
rect 19973 22593 20007 22627
rect 21373 22593 21407 22627
rect 21465 22593 21499 22627
rect 22477 22593 22511 22627
rect 22753 22593 22787 22627
rect 22845 22593 22879 22627
rect 22937 22593 22971 22627
rect 23489 22593 23523 22627
rect 24133 22593 24167 22627
rect 24225 22593 24259 22627
rect 24501 22593 24535 22627
rect 24849 22593 24883 22627
rect 10977 22525 11011 22559
rect 13737 22525 13771 22559
rect 16773 22525 16807 22559
rect 22569 22525 22603 22559
rect 23213 22525 23247 22559
rect 24593 22525 24627 22559
rect 15577 22457 15611 22491
rect 10057 22389 10091 22423
rect 10609 22389 10643 22423
rect 13001 22389 13035 22423
rect 15669 22389 15703 22423
rect 18153 22389 18187 22423
rect 19625 22389 19659 22423
rect 21189 22389 21223 22423
rect 21833 22389 21867 22423
rect 23949 22389 23983 22423
rect 9321 22185 9355 22219
rect 13737 22185 13771 22219
rect 14105 22185 14139 22219
rect 16129 22185 16163 22219
rect 16221 22185 16255 22219
rect 16405 22185 16439 22219
rect 19809 22185 19843 22219
rect 19901 22185 19935 22219
rect 24409 22185 24443 22219
rect 18245 22117 18279 22151
rect 22661 22117 22695 22151
rect 13001 22049 13035 22083
rect 14749 22049 14783 22083
rect 18337 22049 18371 22083
rect 21281 22049 21315 22083
rect 22109 22049 22143 22083
rect 22937 22049 22971 22083
rect 23029 22049 23063 22083
rect 25789 22049 25823 22083
rect 9413 21981 9447 22015
rect 13093 21981 13127 22015
rect 14289 21981 14323 22015
rect 14473 21981 14507 22015
rect 14565 21981 14599 22015
rect 16865 21981 16899 22015
rect 19625 21981 19659 22015
rect 21014 21981 21048 22015
rect 22845 21981 22879 22015
rect 23857 21981 23891 22015
rect 24041 21981 24075 22015
rect 24593 21981 24627 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 25237 21981 25271 22015
rect 12734 21913 12768 21947
rect 14994 21913 15028 21947
rect 16389 21913 16423 21947
rect 16589 21913 16623 21947
rect 17132 21913 17166 21947
rect 21373 21913 21407 21947
rect 23949 21913 23983 21947
rect 11621 21845 11655 21879
rect 18981 21845 19015 21879
rect 12265 21641 12299 21675
rect 15853 21641 15887 21675
rect 16037 21641 16071 21675
rect 17325 21641 17359 21675
rect 17601 21641 17635 21675
rect 17693 21641 17727 21675
rect 17785 21641 17819 21675
rect 18153 21641 18187 21675
rect 21465 21641 21499 21675
rect 25513 21641 25547 21675
rect 17049 21573 17083 21607
rect 18429 21573 18463 21607
rect 18613 21573 18647 21607
rect 19901 21573 19935 21607
rect 23029 21573 23063 21607
rect 7665 21505 7699 21539
rect 12173 21505 12207 21539
rect 12357 21505 12391 21539
rect 14473 21505 14507 21539
rect 14740 21505 14774 21539
rect 16129 21505 16163 21539
rect 16681 21505 16715 21539
rect 16773 21505 16807 21539
rect 17325 21505 17359 21539
rect 18061 21505 18095 21539
rect 18245 21505 18279 21539
rect 18337 21505 18371 21539
rect 20269 21505 20303 21539
rect 21373 21505 21407 21539
rect 21557 21505 21591 21539
rect 22017 21505 22051 21539
rect 22293 21505 22327 21539
rect 22477 21505 22511 21539
rect 22569 21505 22603 21539
rect 22661 21505 22695 21539
rect 22845 21505 22879 21539
rect 23949 21505 23983 21539
rect 24225 21505 24259 21539
rect 24409 21505 24443 21539
rect 24777 21505 24811 21539
rect 25697 21505 25731 21539
rect 25789 21505 25823 21539
rect 7941 21437 7975 21471
rect 23581 21437 23615 21471
rect 25329 21437 25363 21471
rect 17233 21369 17267 21403
rect 17969 21369 18003 21403
rect 18613 21369 18647 21403
rect 9413 21301 9447 21335
rect 17417 21301 17451 21335
rect 21833 21301 21867 21335
rect 22845 21301 22879 21335
rect 23765 21301 23799 21335
rect 18337 21097 18371 21131
rect 22385 21097 22419 21131
rect 25789 21097 25823 21131
rect 16773 21029 16807 21063
rect 17233 21029 17267 21063
rect 15485 20961 15519 20995
rect 24409 20961 24443 20995
rect 8033 20893 8067 20927
rect 8217 20893 8251 20927
rect 8493 20893 8527 20927
rect 8769 20893 8803 20927
rect 9505 20893 9539 20927
rect 10241 20893 10275 20927
rect 10793 20893 10827 20927
rect 11069 20893 11103 20927
rect 16313 20893 16347 20927
rect 16497 20893 16531 20927
rect 16773 20893 16807 20927
rect 16865 20893 16899 20927
rect 17785 20893 17819 20927
rect 18245 20893 18279 20927
rect 18613 20893 18647 20927
rect 21373 20893 21407 20927
rect 22569 20893 22603 20927
rect 22661 20893 22695 20927
rect 22845 20893 22879 20927
rect 22937 20893 22971 20927
rect 23029 20893 23063 20927
rect 23397 20893 23431 20927
rect 23765 20893 23799 20927
rect 24665 20893 24699 20927
rect 8125 20825 8159 20859
rect 11345 20825 11379 20859
rect 16957 20825 16991 20859
rect 17141 20825 17175 20859
rect 22201 20825 22235 20859
rect 8309 20757 8343 20791
rect 8677 20757 8711 20791
rect 8953 20757 8987 20791
rect 9689 20757 9723 20791
rect 10977 20757 11011 20791
rect 12817 20757 12851 20791
rect 16589 20757 16623 20791
rect 17042 20757 17076 20791
rect 18337 20757 18371 20791
rect 18429 20757 18463 20791
rect 23305 20757 23339 20791
rect 11529 20553 11563 20587
rect 11989 20553 12023 20587
rect 18521 20553 18555 20587
rect 21005 20553 21039 20587
rect 23949 20553 23983 20587
rect 24935 20553 24969 20587
rect 10701 20485 10735 20519
rect 16681 20485 16715 20519
rect 22078 20485 22112 20519
rect 23581 20485 23615 20519
rect 24041 20485 24075 20519
rect 25145 20485 25179 20519
rect 7389 20417 7423 20451
rect 7573 20417 7607 20451
rect 7665 20417 7699 20451
rect 7757 20417 7791 20451
rect 8033 20417 8067 20451
rect 9873 20417 9907 20451
rect 11897 20417 11931 20451
rect 13185 20417 13219 20451
rect 13829 20417 13863 20451
rect 14013 20417 14047 20451
rect 15117 20417 15151 20451
rect 15301 20417 15335 20451
rect 15485 20417 15519 20451
rect 15577 20417 15611 20451
rect 16957 20417 16991 20451
rect 17417 20417 17451 20451
rect 17601 20417 17635 20451
rect 17877 20417 17911 20451
rect 19165 20417 19199 20451
rect 20637 20417 20671 20451
rect 20821 20417 20855 20451
rect 21097 20417 21131 20451
rect 23305 20417 23339 20451
rect 23398 20417 23432 20451
rect 23673 20417 23707 20451
rect 23811 20417 23845 20451
rect 8309 20349 8343 20383
rect 12173 20349 12207 20383
rect 13093 20349 13127 20383
rect 16865 20349 16899 20383
rect 17325 20349 17359 20383
rect 21833 20349 21867 20383
rect 24593 20349 24627 20383
rect 7941 20281 7975 20315
rect 13645 20281 13679 20315
rect 18613 20281 18647 20315
rect 23213 20281 23247 20315
rect 9781 20213 9815 20247
rect 13553 20213 13587 20247
rect 15761 20213 15795 20247
rect 16957 20213 16991 20247
rect 17785 20213 17819 20247
rect 20361 20213 20395 20247
rect 20821 20213 20855 20247
rect 24777 20213 24811 20247
rect 24961 20213 24995 20247
rect 8033 20009 8067 20043
rect 9045 20009 9079 20043
rect 9597 20009 9631 20043
rect 15117 20009 15151 20043
rect 17141 20009 17175 20043
rect 18797 20009 18831 20043
rect 21097 20009 21131 20043
rect 23581 20009 23615 20043
rect 16957 19941 16991 19975
rect 21005 19941 21039 19975
rect 14841 19873 14875 19907
rect 15669 19873 15703 19907
rect 19625 19873 19659 19907
rect 21649 19873 21683 19907
rect 22201 19873 22235 19907
rect 7481 19805 7515 19839
rect 7573 19805 7607 19839
rect 8217 19805 8251 19839
rect 8401 19805 8435 19839
rect 8585 19805 8619 19839
rect 8953 19805 8987 19839
rect 9128 19805 9162 19839
rect 9229 19805 9263 19839
rect 9413 19805 9447 19839
rect 9505 19805 9539 19839
rect 11069 19805 11103 19839
rect 13553 19805 13587 19839
rect 14657 19805 14691 19839
rect 15853 19805 15887 19839
rect 17417 19805 17451 19839
rect 17684 19805 17718 19839
rect 19349 19805 19383 19839
rect 19533 19805 19567 19839
rect 8309 19737 8343 19771
rect 11345 19737 11379 19771
rect 16589 19737 16623 19771
rect 17325 19737 17359 19771
rect 19441 19737 19475 19771
rect 19870 19737 19904 19771
rect 22468 19737 22502 19771
rect 7297 19669 7331 19703
rect 7941 19669 7975 19703
rect 9321 19669 9355 19703
rect 12817 19669 12851 19703
rect 13001 19669 13035 19703
rect 14289 19669 14323 19703
rect 14749 19669 14783 19703
rect 17125 19669 17159 19703
rect 7389 19465 7423 19499
rect 8125 19465 8159 19499
rect 9045 19465 9079 19499
rect 9689 19465 9723 19499
rect 12633 19465 12667 19499
rect 18337 19465 18371 19499
rect 22753 19465 22787 19499
rect 9229 19397 9263 19431
rect 11529 19397 11563 19431
rect 11897 19397 11931 19431
rect 17132 19397 17166 19431
rect 21005 19397 21039 19431
rect 22477 19397 22511 19431
rect 1777 19329 1811 19363
rect 6377 19329 6411 19363
rect 8309 19329 8343 19363
rect 8493 19329 8527 19363
rect 8769 19329 8803 19363
rect 9137 19329 9171 19363
rect 9689 19329 9723 19363
rect 9873 19329 9907 19363
rect 9965 19329 9999 19363
rect 10241 19329 10275 19363
rect 10517 19329 10551 19363
rect 10609 19329 10643 19363
rect 11161 19329 11195 19363
rect 11345 19329 11379 19363
rect 11713 19329 11747 19363
rect 11805 19329 11839 19363
rect 12015 19329 12049 19363
rect 12265 19329 12299 19363
rect 12449 19329 12483 19363
rect 14381 19329 14415 19363
rect 19073 19329 19107 19363
rect 21281 19329 21315 19363
rect 22753 19329 22787 19363
rect 8033 19261 8067 19295
rect 10149 19261 10183 19295
rect 10977 19261 11011 19295
rect 12173 19261 12207 19295
rect 14105 19261 14139 19295
rect 15945 19261 15979 19295
rect 16221 19261 16255 19295
rect 16865 19261 16899 19295
rect 18889 19261 18923 19295
rect 19349 19261 19383 19295
rect 22661 19261 22695 19295
rect 9413 19193 9447 19227
rect 10425 19193 10459 19227
rect 18245 19193 18279 19227
rect 19533 19193 19567 19227
rect 1501 19125 1535 19159
rect 6561 19125 6595 19159
rect 8493 19125 8527 19159
rect 8861 19125 8895 19159
rect 10149 19125 10183 19159
rect 12265 19125 12299 19159
rect 14473 19125 14507 19159
rect 19165 19125 19199 19159
rect 19257 19125 19291 19159
rect 7941 18921 7975 18955
rect 12541 18921 12575 18955
rect 14473 18921 14507 18955
rect 18429 18921 18463 18955
rect 7849 18853 7883 18887
rect 20361 18853 20395 18887
rect 6101 18785 6135 18819
rect 8401 18785 8435 18819
rect 8493 18785 8527 18819
rect 13461 18785 13495 18819
rect 13737 18785 13771 18819
rect 14105 18785 14139 18819
rect 15945 18785 15979 18819
rect 9229 18717 9263 18751
rect 9321 18717 9355 18751
rect 9413 18717 9447 18751
rect 9689 18717 9723 18751
rect 9781 18717 9815 18751
rect 10425 18717 10459 18751
rect 11989 18717 12023 18751
rect 12357 18717 12391 18751
rect 13185 18717 13219 18751
rect 13553 18717 13587 18751
rect 13645 18717 13679 18751
rect 14289 18717 14323 18751
rect 14381 18717 14415 18751
rect 16221 18717 16255 18751
rect 17049 18717 17083 18751
rect 17316 18717 17350 18751
rect 20177 18717 20211 18751
rect 20453 18717 20487 18751
rect 22845 18717 22879 18751
rect 6377 18649 6411 18683
rect 9531 18649 9565 18683
rect 10517 18649 10551 18683
rect 11253 18649 11287 18683
rect 12173 18649 12207 18683
rect 12265 18649 12299 18683
rect 12633 18649 12667 18683
rect 8309 18581 8343 18615
rect 9045 18581 9079 18615
rect 13921 18581 13955 18615
rect 14105 18581 14139 18615
rect 19993 18581 20027 18615
rect 23029 18581 23063 18615
rect 2145 18377 2179 18411
rect 8125 18377 8159 18411
rect 8217 18377 8251 18411
rect 12173 18377 12207 18411
rect 15117 18377 15151 18411
rect 6653 18309 6687 18343
rect 8953 18309 8987 18343
rect 15301 18309 15335 18343
rect 19441 18309 19475 18343
rect 23397 18309 23431 18343
rect 2329 18241 2363 18275
rect 8401 18241 8435 18275
rect 8677 18241 8711 18275
rect 10517 18241 10551 18275
rect 10609 18241 10643 18275
rect 10793 18241 10827 18275
rect 10893 18241 10927 18275
rect 11253 18241 11287 18275
rect 11345 18241 11379 18275
rect 12081 18241 12115 18275
rect 12173 18241 12207 18275
rect 12357 18241 12391 18275
rect 13093 18241 13127 18275
rect 13369 18241 13403 18275
rect 13829 18241 13863 18275
rect 14473 18241 14507 18275
rect 15209 18241 15243 18275
rect 19165 18241 19199 18275
rect 22753 18241 22787 18275
rect 23121 18241 23155 18275
rect 6377 18173 6411 18207
rect 8585 18173 8619 18207
rect 11805 18173 11839 18207
rect 13185 18173 13219 18207
rect 13277 18173 13311 18207
rect 13645 18173 13679 18207
rect 23029 18173 23063 18207
rect 25145 18173 25179 18207
rect 10425 18105 10459 18139
rect 11069 18037 11103 18071
rect 11529 18037 11563 18071
rect 11989 18037 12023 18071
rect 13553 18037 13587 18071
rect 14013 18037 14047 18071
rect 20913 18037 20947 18071
rect 22569 18037 22603 18071
rect 22937 18037 22971 18071
rect 8125 17833 8159 17867
rect 8401 17833 8435 17867
rect 9137 17833 9171 17867
rect 12357 17833 12391 17867
rect 22201 17833 22235 17867
rect 23213 17833 23247 17867
rect 12541 17765 12575 17799
rect 5733 17697 5767 17731
rect 10425 17697 10459 17731
rect 22109 17697 22143 17731
rect 23857 17697 23891 17731
rect 24409 17697 24443 17731
rect 6469 17629 6503 17663
rect 8401 17629 8435 17663
rect 8585 17629 8619 17663
rect 8953 17629 8987 17663
rect 9137 17629 9171 17663
rect 10149 17629 10183 17663
rect 10793 17629 10827 17663
rect 10977 17629 11011 17663
rect 11253 17629 11287 17663
rect 11345 17629 11379 17663
rect 12081 17629 12115 17663
rect 12173 17629 12207 17663
rect 14565 17629 14599 17663
rect 18153 17629 18187 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 18705 17629 18739 17663
rect 19809 17629 19843 17663
rect 22753 17629 22787 17663
rect 22937 17629 22971 17663
rect 23121 17629 23155 17663
rect 24225 17629 24259 17663
rect 5457 17561 5491 17595
rect 5917 17561 5951 17595
rect 12725 17561 12759 17595
rect 20085 17561 20119 17595
rect 21833 17561 21867 17595
rect 24685 17561 24719 17595
rect 5089 17493 5123 17527
rect 5549 17493 5583 17527
rect 9965 17493 9999 17527
rect 11805 17493 11839 17527
rect 14841 17493 14875 17527
rect 17509 17493 17543 17527
rect 18613 17493 18647 17527
rect 19257 17493 19291 17527
rect 22937 17493 22971 17527
rect 23581 17493 23615 17527
rect 23673 17493 23707 17527
rect 24133 17493 24167 17527
rect 26157 17493 26191 17527
rect 11621 17289 11655 17323
rect 12449 17289 12483 17323
rect 13737 17289 13771 17323
rect 18429 17289 18463 17323
rect 18889 17289 18923 17323
rect 20729 17289 20763 17323
rect 21925 17289 21959 17323
rect 22753 17289 22787 17323
rect 25053 17289 25087 17323
rect 16313 17221 16347 17255
rect 16957 17221 16991 17255
rect 19257 17221 19291 17255
rect 6193 17153 6227 17187
rect 11529 17153 11563 17187
rect 12173 17153 12207 17187
rect 12265 17153 12299 17187
rect 12541 17153 12575 17187
rect 12725 17153 12759 17187
rect 13921 17153 13955 17187
rect 14013 17153 14047 17187
rect 14197 17153 14231 17187
rect 15209 17153 15243 17187
rect 16129 17153 16163 17187
rect 16221 17153 16255 17187
rect 18613 17153 18647 17187
rect 21373 17153 21407 17187
rect 22109 17153 22143 17187
rect 22201 17153 22235 17187
rect 22293 17153 22327 17187
rect 22411 17153 22445 17187
rect 22661 17153 22695 17187
rect 23305 17153 23339 17187
rect 25421 17153 25455 17187
rect 2421 17085 2455 17119
rect 2697 17085 2731 17119
rect 4169 17085 4203 17119
rect 4905 17085 4939 17119
rect 5457 17085 5491 17119
rect 6469 17085 6503 17119
rect 10609 17085 10643 17119
rect 15025 17085 15059 17119
rect 15485 17085 15519 17119
rect 16681 17085 16715 17119
rect 18889 17085 18923 17119
rect 18981 17085 19015 17119
rect 22569 17085 22603 17119
rect 23121 17085 23155 17119
rect 23581 17085 23615 17119
rect 12633 17017 12667 17051
rect 14013 17017 14047 17051
rect 4261 16949 4295 16983
rect 7113 16949 7147 16983
rect 11253 16949 11287 16983
rect 14381 16949 14415 16983
rect 15301 16949 15335 16983
rect 18705 16949 18739 16983
rect 20821 16949 20855 16983
rect 22937 16949 22971 16983
rect 25973 16949 26007 16983
rect 3249 16745 3283 16779
rect 8045 16745 8079 16779
rect 16484 16745 16518 16779
rect 18889 16745 18923 16779
rect 20361 16745 20395 16779
rect 21281 16745 21315 16779
rect 21649 16745 21683 16779
rect 23121 16745 23155 16779
rect 24225 16745 24259 16779
rect 25145 16745 25179 16779
rect 12173 16677 12207 16711
rect 18797 16677 18831 16711
rect 21097 16677 21131 16711
rect 21833 16677 21867 16711
rect 22109 16677 22143 16711
rect 4721 16609 4755 16643
rect 8309 16609 8343 16643
rect 9597 16609 9631 16643
rect 10425 16609 10459 16643
rect 12265 16609 12299 16643
rect 13921 16609 13955 16643
rect 14105 16609 14139 16643
rect 15577 16609 15611 16643
rect 15853 16609 15887 16643
rect 16221 16609 16255 16643
rect 17969 16609 18003 16643
rect 18153 16609 18187 16643
rect 22201 16609 22235 16643
rect 22329 16609 22363 16643
rect 22661 16609 22695 16643
rect 25053 16609 25087 16643
rect 25789 16609 25823 16643
rect 3433 16541 3467 16575
rect 3985 16541 4019 16575
rect 4445 16541 4479 16575
rect 12357 16541 12391 16575
rect 12541 16541 12575 16575
rect 12909 16541 12943 16575
rect 13001 16541 13035 16575
rect 18889 16541 18923 16575
rect 19073 16541 19107 16575
rect 19257 16541 19291 16575
rect 19993 16541 20027 16575
rect 20177 16541 20211 16575
rect 20821 16541 20855 16575
rect 21097 16541 21131 16575
rect 21189 16541 21223 16575
rect 22017 16541 22051 16575
rect 22477 16541 22511 16575
rect 23029 16541 23063 16575
rect 23305 16541 23339 16575
rect 23765 16541 23799 16575
rect 24409 16541 24443 16575
rect 25329 16541 25363 16575
rect 25881 16541 25915 16575
rect 4169 16473 4203 16507
rect 4353 16473 4387 16507
rect 4997 16473 5031 16507
rect 10701 16473 10735 16507
rect 22845 16473 22879 16507
rect 23397 16473 23431 16507
rect 23489 16473 23523 16507
rect 23607 16473 23641 16507
rect 23857 16473 23891 16507
rect 24041 16473 24075 16507
rect 25421 16473 25455 16507
rect 25514 16473 25548 16507
rect 25651 16473 25685 16507
rect 25973 16473 26007 16507
rect 4629 16405 4663 16439
rect 6469 16405 6503 16439
rect 6561 16405 6595 16439
rect 8953 16405 8987 16439
rect 12725 16405 12759 16439
rect 13277 16405 13311 16439
rect 19901 16405 19935 16439
rect 20913 16405 20947 16439
rect 5641 16201 5675 16235
rect 6009 16201 6043 16235
rect 9597 16201 9631 16235
rect 18429 16201 18463 16235
rect 19625 16201 19659 16235
rect 19809 16201 19843 16235
rect 19993 16201 20027 16235
rect 23305 16201 23339 16235
rect 25053 16201 25087 16235
rect 6377 16133 6411 16167
rect 7113 16133 7147 16167
rect 7941 16133 7975 16167
rect 25329 16133 25363 16167
rect 25941 16133 25975 16167
rect 26157 16133 26191 16167
rect 5733 16065 5767 16099
rect 7573 16065 7607 16099
rect 7665 16065 7699 16099
rect 11345 16065 11379 16099
rect 12541 16065 12575 16099
rect 15761 16065 15795 16099
rect 16405 16065 16439 16099
rect 16681 16065 16715 16099
rect 19073 16065 19107 16099
rect 19257 16065 19291 16099
rect 19349 16065 19383 16099
rect 19901 16065 19935 16099
rect 20177 16065 20211 16099
rect 23121 16065 23155 16099
rect 23305 16065 23339 16099
rect 24593 16065 24627 16099
rect 24869 16065 24903 16099
rect 25421 16065 25455 16099
rect 25513 16065 25547 16099
rect 1593 15997 1627 16031
rect 1869 15997 1903 16031
rect 3617 15997 3651 16031
rect 3893 15997 3927 16031
rect 4169 15997 4203 16031
rect 6009 15997 6043 16031
rect 11069 15997 11103 16031
rect 12909 15997 12943 16031
rect 13553 15997 13587 16031
rect 13829 15997 13863 16031
rect 15853 15997 15887 16031
rect 15945 15997 15979 16031
rect 16957 15997 16991 16031
rect 24685 15997 24719 16031
rect 24777 15997 24811 16031
rect 5825 15929 5859 15963
rect 7389 15929 7423 15963
rect 9413 15929 9447 15963
rect 15393 15929 15427 15963
rect 16221 15929 16255 15963
rect 25145 15929 25179 15963
rect 11989 15861 12023 15895
rect 13461 15861 13495 15895
rect 15301 15861 15335 15895
rect 18521 15861 18555 15895
rect 19441 15861 19475 15895
rect 25697 15861 25731 15895
rect 25789 15861 25823 15895
rect 25973 15861 26007 15895
rect 2145 15657 2179 15691
rect 3065 15657 3099 15691
rect 3433 15657 3467 15691
rect 6285 15657 6319 15691
rect 13001 15657 13035 15691
rect 13737 15657 13771 15691
rect 15853 15657 15887 15691
rect 21281 15657 21315 15691
rect 16773 15589 16807 15623
rect 16957 15589 16991 15623
rect 5457 15521 5491 15555
rect 6745 15521 6779 15555
rect 8493 15521 8527 15555
rect 8953 15521 8987 15555
rect 9689 15521 9723 15555
rect 10425 15521 10459 15555
rect 12173 15521 12207 15555
rect 12817 15521 12851 15555
rect 14105 15521 14139 15555
rect 14381 15521 14415 15555
rect 17601 15521 17635 15555
rect 19533 15521 19567 15555
rect 22477 15521 22511 15555
rect 22753 15521 22787 15555
rect 1409 15453 1443 15487
rect 2329 15453 2363 15487
rect 3157 15453 3191 15487
rect 3617 15453 3651 15487
rect 5273 15453 5307 15487
rect 5365 15453 5399 15487
rect 6377 15453 6411 15487
rect 6469 15453 6503 15487
rect 6653 15453 6687 15487
rect 13185 15453 13219 15487
rect 13461 15453 13495 15487
rect 13921 15453 13955 15487
rect 16589 15453 16623 15487
rect 18613 15453 18647 15487
rect 18705 15453 18739 15487
rect 19257 15453 19291 15487
rect 21189 15453 21223 15487
rect 22385 15453 22419 15487
rect 24685 15453 24719 15487
rect 24961 15453 24995 15487
rect 26065 15453 26099 15487
rect 6561 15385 6595 15419
rect 7021 15385 7055 15419
rect 10701 15385 10735 15419
rect 17325 15385 17359 15419
rect 1593 15317 1627 15351
rect 4905 15317 4939 15351
rect 9597 15317 9631 15351
rect 10333 15317 10367 15351
rect 12265 15317 12299 15351
rect 13369 15317 13403 15351
rect 17417 15317 17451 15351
rect 17969 15317 18003 15351
rect 18797 15317 18831 15351
rect 21005 15317 21039 15351
rect 24501 15317 24535 15351
rect 24869 15317 24903 15351
rect 25421 15317 25455 15351
rect 6561 15113 6595 15147
rect 9229 15113 9263 15147
rect 10057 15113 10091 15147
rect 10425 15113 10459 15147
rect 10885 15113 10919 15147
rect 11529 15113 11563 15147
rect 11897 15113 11931 15147
rect 24225 15113 24259 15147
rect 26065 15113 26099 15147
rect 19901 15045 19935 15079
rect 23121 15045 23155 15079
rect 23857 15045 23891 15079
rect 24593 15045 24627 15079
rect 6653 14977 6687 15011
rect 7389 14977 7423 15011
rect 9965 14977 9999 15011
rect 10241 14977 10275 15011
rect 10517 14977 10551 15011
rect 11069 14977 11103 15011
rect 12357 14977 12391 15011
rect 12541 14977 12575 15011
rect 13829 14977 13863 15011
rect 17141 14977 17175 15011
rect 19349 14977 19383 15011
rect 22385 14977 22419 15011
rect 23397 14977 23431 15011
rect 23765 14977 23799 15011
rect 24041 14977 24075 15011
rect 1593 14909 1627 14943
rect 1869 14909 1903 14943
rect 3617 14909 3651 14943
rect 7665 14909 7699 14943
rect 9781 14909 9815 14943
rect 11989 14909 12023 14943
rect 12081 14909 12115 14943
rect 17417 14909 17451 14943
rect 18889 14909 18923 14943
rect 19625 14909 19659 14943
rect 23029 14909 23063 14943
rect 23305 14909 23339 14943
rect 24317 14909 24351 14943
rect 19533 14841 19567 14875
rect 9137 14773 9171 14807
rect 10609 14773 10643 14807
rect 12357 14773 12391 14807
rect 15117 14773 15151 14807
rect 21373 14773 21407 14807
rect 23121 14773 23155 14807
rect 23581 14773 23615 14807
rect 2329 14569 2363 14603
rect 7757 14569 7791 14603
rect 10241 14569 10275 14603
rect 12344 14569 12378 14603
rect 14933 14569 14967 14603
rect 17601 14569 17635 14603
rect 20177 14569 20211 14603
rect 22845 14569 22879 14603
rect 23857 14569 23891 14603
rect 8033 14501 8067 14535
rect 10609 14501 10643 14535
rect 14565 14501 14599 14535
rect 18705 14501 18739 14535
rect 23397 14501 23431 14535
rect 2973 14433 3007 14467
rect 8585 14433 8619 14467
rect 12081 14433 12115 14467
rect 14841 14433 14875 14467
rect 20821 14433 20855 14467
rect 22293 14433 22327 14467
rect 22477 14433 22511 14467
rect 23029 14433 23063 14467
rect 24961 14433 24995 14467
rect 2145 14365 2179 14399
rect 2237 14365 2271 14399
rect 3341 14365 3375 14399
rect 3617 14365 3651 14399
rect 5365 14365 5399 14399
rect 5549 14365 5583 14399
rect 6745 14365 6779 14399
rect 7941 14365 7975 14399
rect 9505 14365 9539 14399
rect 10241 14365 10275 14399
rect 10333 14365 10367 14399
rect 14933 14365 14967 14399
rect 16129 14365 16163 14399
rect 16589 14365 16623 14399
rect 17509 14365 17543 14399
rect 18245 14365 18279 14399
rect 18337 14365 18371 14399
rect 18521 14365 18555 14399
rect 18613 14365 18647 14399
rect 18797 14365 18831 14399
rect 19257 14365 19291 14399
rect 19441 14365 19475 14399
rect 20637 14365 20671 14399
rect 21557 14365 21591 14399
rect 22661 14365 22695 14399
rect 23213 14365 23247 14399
rect 23765 14365 23799 14399
rect 23857 14365 23891 14399
rect 24133 14365 24167 14399
rect 25237 14365 25271 14399
rect 25421 14365 25455 14399
rect 1961 14297 1995 14331
rect 3525 14297 3559 14331
rect 9781 14297 9815 14331
rect 20545 14297 20579 14331
rect 21005 14297 21039 14331
rect 23949 14297 23983 14331
rect 24869 14297 24903 14331
rect 2237 14229 2271 14263
rect 2697 14229 2731 14263
rect 2789 14229 2823 14263
rect 3157 14229 3191 14263
rect 5365 14229 5399 14263
rect 7389 14229 7423 14263
rect 8401 14229 8435 14263
rect 8493 14229 8527 14263
rect 8953 14229 8987 14263
rect 10057 14229 10091 14263
rect 13829 14229 13863 14263
rect 15577 14229 15611 14263
rect 16681 14229 16715 14263
rect 16865 14229 16899 14263
rect 19349 14229 19383 14263
rect 21741 14229 21775 14263
rect 23581 14229 23615 14263
rect 24409 14229 24443 14263
rect 24777 14229 24811 14263
rect 25605 14229 25639 14263
rect 2329 14025 2363 14059
rect 3433 14025 3467 14059
rect 6009 14025 6043 14059
rect 15945 14025 15979 14059
rect 16405 14025 16439 14059
rect 24133 14025 24167 14059
rect 2605 13957 2639 13991
rect 3617 13957 3651 13991
rect 4813 13957 4847 13991
rect 5273 13957 5307 13991
rect 8677 13957 8711 13991
rect 13461 13957 13495 13991
rect 2513 13889 2547 13923
rect 2697 13889 2731 13923
rect 2835 13889 2869 13923
rect 3249 13889 3283 13923
rect 3341 13889 3375 13923
rect 4537 13889 4571 13923
rect 5089 13889 5123 13923
rect 5181 13889 5215 13923
rect 5391 13889 5425 13923
rect 5549 13889 5583 13923
rect 5825 13889 5859 13923
rect 6101 13889 6135 13923
rect 8953 13889 8987 13923
rect 9137 13889 9171 13923
rect 11529 13889 11563 13923
rect 11713 13889 11747 13923
rect 13093 13889 13127 13923
rect 13277 13889 13311 13923
rect 13369 13889 13403 13923
rect 14197 13889 14231 13923
rect 16221 13889 16255 13923
rect 16497 13889 16531 13923
rect 19349 13889 19383 13923
rect 22201 13889 22235 13923
rect 22385 13889 22419 13923
rect 23489 13889 23523 13923
rect 23581 13889 23615 13923
rect 24041 13889 24075 13923
rect 24225 13889 24259 13923
rect 24777 13889 24811 13923
rect 24869 13889 24903 13923
rect 25053 13889 25087 13923
rect 2973 13821 3007 13855
rect 4813 13821 4847 13855
rect 14105 13821 14139 13855
rect 14473 13821 14507 13855
rect 16037 13821 16071 13855
rect 16681 13821 16715 13855
rect 19073 13821 19107 13855
rect 19717 13821 19751 13855
rect 20085 13821 20119 13855
rect 24685 13821 24719 13855
rect 10885 13753 10919 13787
rect 22293 13753 22327 13787
rect 3065 13685 3099 13719
rect 4629 13685 4663 13719
rect 4905 13685 4939 13719
rect 5641 13685 5675 13719
rect 7205 13685 7239 13719
rect 9394 13685 9428 13719
rect 11621 13685 11655 13719
rect 12909 13685 12943 13719
rect 17325 13685 17359 13719
rect 17601 13685 17635 13719
rect 21511 13685 21545 13719
rect 23213 13685 23247 13719
rect 23581 13685 23615 13719
rect 25053 13685 25087 13719
rect 3249 13481 3283 13515
rect 7205 13481 7239 13515
rect 8033 13481 8067 13515
rect 8953 13481 8987 13515
rect 14565 13481 14599 13515
rect 15393 13481 15427 13515
rect 18245 13481 18279 13515
rect 18337 13481 18371 13515
rect 20453 13481 20487 13515
rect 23857 13481 23891 13515
rect 25697 13481 25731 13515
rect 3157 13413 3191 13447
rect 8309 13413 8343 13447
rect 9689 13413 9723 13447
rect 25421 13413 25455 13447
rect 25513 13413 25547 13447
rect 1409 13345 1443 13379
rect 4721 13345 4755 13379
rect 4997 13345 5031 13379
rect 6745 13345 6779 13379
rect 8401 13345 8435 13379
rect 9597 13345 9631 13379
rect 10333 13345 10367 13379
rect 11345 13345 11379 13379
rect 11713 13345 11747 13379
rect 13277 13345 13311 13379
rect 15715 13345 15749 13379
rect 17141 13345 17175 13379
rect 17509 13345 17543 13379
rect 18981 13345 19015 13379
rect 3433 13277 3467 13311
rect 3617 13277 3651 13311
rect 4445 13277 4479 13311
rect 8217 13277 8251 13311
rect 8493 13277 8527 13311
rect 10609 13277 10643 13311
rect 15209 13277 15243 13311
rect 15485 13277 15519 13311
rect 17601 13277 17635 13311
rect 19441 13277 19475 13311
rect 19809 13277 19843 13311
rect 20361 13277 20395 13311
rect 20545 13277 20579 13311
rect 21097 13277 21131 13311
rect 23489 13277 23523 13311
rect 24593 13277 24627 13311
rect 24961 13277 24995 13311
rect 25053 13277 25087 13311
rect 26157 13277 26191 13311
rect 1685 13209 1719 13243
rect 6837 13209 6871 13243
rect 7021 13209 7055 13243
rect 19533 13209 19567 13243
rect 19625 13209 19659 13243
rect 24041 13209 24075 13243
rect 24225 13209 24259 13243
rect 24685 13209 24719 13243
rect 24777 13209 24811 13243
rect 25237 13209 25271 13243
rect 25676 13209 25710 13243
rect 25881 13209 25915 13243
rect 3801 13141 3835 13175
rect 11253 13141 11287 13175
rect 13139 13141 13173 13175
rect 13921 13141 13955 13175
rect 19257 13141 19291 13175
rect 21005 13141 21039 13175
rect 23305 13141 23339 13175
rect 24409 13141 24443 13175
rect 25973 13141 26007 13175
rect 2329 12937 2363 12971
rect 3065 12937 3099 12971
rect 7573 12937 7607 12971
rect 9045 12937 9079 12971
rect 9321 12937 9355 12971
rect 15439 12937 15473 12971
rect 25329 12937 25363 12971
rect 2605 12869 2639 12903
rect 2835 12869 2869 12903
rect 21557 12869 21591 12903
rect 23949 12869 23983 12903
rect 24041 12869 24075 12903
rect 24179 12869 24213 12903
rect 25513 12869 25547 12903
rect 2513 12801 2547 12835
rect 2697 12801 2731 12835
rect 3801 12801 3835 12835
rect 4787 12801 4821 12835
rect 4905 12801 4939 12835
rect 4997 12801 5031 12835
rect 5089 12801 5123 12835
rect 5549 12801 5583 12835
rect 6377 12801 6411 12835
rect 6653 12801 6687 12835
rect 8953 12801 8987 12835
rect 9137 12801 9171 12835
rect 14013 12801 14047 12835
rect 16865 12801 16899 12835
rect 20177 12801 20211 12835
rect 20453 12801 20487 12835
rect 20913 12801 20947 12835
rect 21189 12801 21223 12835
rect 21373 12801 21407 12835
rect 21465 12801 21499 12835
rect 21649 12801 21683 12835
rect 22109 12801 22143 12835
rect 23213 12801 23247 12835
rect 23581 12801 23615 12835
rect 23857 12801 23891 12835
rect 25237 12801 25271 12835
rect 25421 12801 25455 12835
rect 26157 12801 26191 12835
rect 2973 12733 3007 12767
rect 3249 12733 3283 12767
rect 3341 12733 3375 12767
rect 3433 12733 3467 12767
rect 3525 12733 3559 12767
rect 4629 12733 4663 12767
rect 5457 12733 5491 12767
rect 5917 12733 5951 12767
rect 6469 12733 6503 12767
rect 8125 12733 8159 12767
rect 10793 12733 10827 12767
rect 11069 12733 11103 12767
rect 11621 12733 11655 12767
rect 11897 12733 11931 12767
rect 13645 12733 13679 12767
rect 17141 12733 17175 12767
rect 20637 12733 20671 12767
rect 24317 12733 24351 12767
rect 24409 12733 24443 12767
rect 24961 12733 24995 12767
rect 3893 12665 3927 12699
rect 18613 12665 18647 12699
rect 5273 12597 5307 12631
rect 6377 12597 6411 12631
rect 6837 12597 6871 12631
rect 13369 12597 13403 12631
rect 20269 12597 20303 12631
rect 20729 12597 20763 12631
rect 21925 12597 21959 12631
rect 23673 12597 23707 12631
rect 4997 12393 5031 12427
rect 6285 12393 6319 12427
rect 12265 12393 12299 12427
rect 13737 12393 13771 12427
rect 14565 12393 14599 12427
rect 24225 12393 24259 12427
rect 26157 12393 26191 12427
rect 5273 12325 5307 12359
rect 6469 12325 6503 12359
rect 3985 12257 4019 12291
rect 4997 12257 5031 12291
rect 9229 12257 9263 12291
rect 12633 12257 12667 12291
rect 12817 12257 12851 12291
rect 19441 12257 19475 12291
rect 20545 12257 20579 12291
rect 22477 12257 22511 12291
rect 24409 12257 24443 12291
rect 3893 12189 3927 12223
rect 4721 12189 4755 12223
rect 5365 12189 5399 12223
rect 5549 12189 5583 12223
rect 5733 12189 5767 12223
rect 6101 12189 6135 12223
rect 6285 12189 6319 12223
rect 6561 12189 6595 12223
rect 6929 12189 6963 12223
rect 7113 12189 7147 12223
rect 8493 12189 8527 12223
rect 8677 12189 8711 12223
rect 9597 12189 9631 12223
rect 11713 12189 11747 12223
rect 12449 12189 12483 12223
rect 12725 12189 12759 12223
rect 13001 12189 13035 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 13737 12189 13771 12223
rect 14749 12189 14783 12223
rect 14841 12189 14875 12223
rect 14933 12189 14967 12223
rect 15117 12189 15151 12223
rect 19257 12189 19291 12223
rect 19533 12189 19567 12223
rect 19625 12189 19659 12223
rect 19717 12189 19751 12223
rect 20269 12189 20303 12223
rect 20453 12189 20487 12223
rect 5825 12121 5859 12155
rect 11023 12121 11057 12155
rect 20821 12121 20855 12155
rect 22753 12121 22787 12155
rect 24685 12121 24719 12155
rect 6745 12053 6779 12087
rect 7021 12053 7055 12087
rect 8585 12053 8619 12087
rect 11161 12053 11195 12087
rect 13921 12053 13955 12087
rect 19901 12053 19935 12087
rect 20361 12053 20395 12087
rect 22293 12053 22327 12087
rect 9229 11849 9263 11883
rect 10057 11849 10091 11883
rect 11161 11849 11195 11883
rect 12909 11849 12943 11883
rect 17785 11849 17819 11883
rect 20085 11849 20119 11883
rect 20545 11849 20579 11883
rect 24409 11849 24443 11883
rect 2881 11781 2915 11815
rect 3985 11781 4019 11815
rect 4169 11781 4203 11815
rect 9689 11781 9723 11815
rect 18705 11781 18739 11815
rect 20453 11781 20487 11815
rect 2789 11713 2823 11747
rect 2973 11713 3007 11747
rect 3157 11713 3191 11747
rect 3249 11713 3283 11747
rect 3893 11713 3927 11747
rect 4445 11713 4479 11747
rect 4813 11713 4847 11747
rect 4997 11713 5031 11747
rect 5549 11713 5583 11747
rect 5733 11713 5767 11747
rect 5825 11713 5859 11747
rect 6009 11713 6043 11747
rect 7021 11713 7055 11747
rect 8953 11713 8987 11747
rect 9597 11713 9631 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 10977 11713 11011 11747
rect 11253 11713 11287 11747
rect 12817 11713 12851 11747
rect 13001 11713 13035 11747
rect 13829 11713 13863 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 14381 11713 14415 11747
rect 14841 11713 14875 11747
rect 14933 11713 14967 11747
rect 15025 11713 15059 11747
rect 15209 11713 15243 11747
rect 15301 11713 15335 11747
rect 15393 11713 15427 11747
rect 15577 11713 15611 11747
rect 15669 11713 15703 11747
rect 15847 11713 15881 11747
rect 15935 11713 15969 11747
rect 16129 11713 16163 11747
rect 17693 11713 17727 11747
rect 17877 11713 17911 11747
rect 17969 11713 18003 11747
rect 19625 11713 19659 11747
rect 19717 11713 19751 11747
rect 19901 11713 19935 11747
rect 21189 11713 21223 11747
rect 22661 11713 22695 11747
rect 5917 11645 5951 11679
rect 6653 11645 6687 11679
rect 10701 11645 10735 11679
rect 10793 11645 10827 11679
rect 14197 11645 14231 11679
rect 20729 11645 20763 11679
rect 22937 11645 22971 11679
rect 4353 11577 4387 11611
rect 9413 11577 9447 11611
rect 21097 11577 21131 11611
rect 2605 11509 2639 11543
rect 4629 11509 4663 11543
rect 4997 11509 5031 11543
rect 5365 11509 5399 11543
rect 8447 11509 8481 11543
rect 14565 11509 14599 11543
rect 14657 11509 14691 11543
rect 15393 11509 15427 11543
rect 15669 11509 15703 11543
rect 16037 11509 16071 11543
rect 18981 11509 19015 11543
rect 19717 11509 19751 11543
rect 1672 11305 1706 11339
rect 3157 11305 3191 11339
rect 3985 11305 4019 11339
rect 4629 11305 4663 11339
rect 4813 11305 4847 11339
rect 6009 11305 6043 11339
rect 14565 11305 14599 11339
rect 15945 11305 15979 11339
rect 16405 11305 16439 11339
rect 5549 11237 5583 11271
rect 14657 11237 14691 11271
rect 1409 11169 1443 11203
rect 3249 11169 3283 11203
rect 6469 11169 6503 11203
rect 7849 11169 7883 11203
rect 8769 11169 8803 11203
rect 9413 11169 9447 11203
rect 9505 11169 9539 11203
rect 17601 11169 17635 11203
rect 17877 11169 17911 11203
rect 19257 11169 19291 11203
rect 19533 11169 19567 11203
rect 21281 11169 21315 11203
rect 22477 11169 22511 11203
rect 3433 11101 3467 11135
rect 4997 11101 5031 11135
rect 5181 11101 5215 11135
rect 5365 11101 5399 11135
rect 6377 11101 6411 11135
rect 6561 11101 6595 11135
rect 8033 11101 8067 11135
rect 8493 11101 8527 11135
rect 8677 11101 8711 11135
rect 9321 11101 9355 11135
rect 14381 11101 14415 11135
rect 14565 11101 14599 11135
rect 14795 11101 14829 11135
rect 15208 11101 15242 11135
rect 15301 11101 15335 11135
rect 15761 11101 15795 11135
rect 16221 11101 16255 11135
rect 17509 11101 17543 11135
rect 18245 11101 18279 11135
rect 18521 11101 18555 11135
rect 18705 11101 18739 11135
rect 21649 11101 21683 11135
rect 3617 11033 3651 11067
rect 3953 11033 3987 11067
rect 4169 11033 4203 11067
rect 4445 11033 4479 11067
rect 5273 11033 5307 11067
rect 5641 11033 5675 11067
rect 5825 11033 5859 11067
rect 8217 11033 8251 11067
rect 14933 11033 14967 11067
rect 15025 11033 15059 11067
rect 15577 11033 15611 11067
rect 16037 11033 16071 11067
rect 16497 11033 16531 11067
rect 16681 11033 16715 11067
rect 18613 11033 18647 11067
rect 3801 10965 3835 10999
rect 4645 10965 4679 10999
rect 8309 10965 8343 10999
rect 8953 10965 8987 10999
rect 15393 10965 15427 10999
rect 2605 10761 2639 10795
rect 2973 10761 3007 10795
rect 5549 10761 5583 10795
rect 6929 10761 6963 10795
rect 7389 10761 7423 10795
rect 9781 10761 9815 10795
rect 14657 10761 14691 10795
rect 14749 10761 14783 10795
rect 15117 10761 15151 10795
rect 3065 10693 3099 10727
rect 4353 10693 4387 10727
rect 4583 10693 4617 10727
rect 6561 10693 6595 10727
rect 8309 10693 8343 10727
rect 12357 10693 12391 10727
rect 15393 10693 15427 10727
rect 16773 10693 16807 10727
rect 17877 10693 17911 10727
rect 19625 10693 19659 10727
rect 20545 10693 20579 10727
rect 21833 10693 21867 10727
rect 2329 10625 2363 10659
rect 3709 10625 3743 10659
rect 3801 10625 3835 10659
rect 3893 10625 3927 10659
rect 4262 10647 4296 10681
rect 4445 10625 4479 10659
rect 5365 10625 5399 10659
rect 6377 10625 6411 10659
rect 7297 10625 7331 10659
rect 8033 10625 8067 10659
rect 11161 10625 11195 10659
rect 12173 10625 12207 10659
rect 12449 10625 12483 10659
rect 15296 10625 15330 10659
rect 15485 10625 15519 10659
rect 15613 10625 15647 10659
rect 15761 10625 15795 10659
rect 16405 10625 16439 10659
rect 16681 10625 16715 10659
rect 16865 10625 16899 10659
rect 16957 10625 16991 10659
rect 17601 10625 17635 10659
rect 19717 10625 19751 10659
rect 19901 10625 19935 10659
rect 20269 10625 20303 10659
rect 3249 10557 3283 10591
rect 4721 10557 4755 10591
rect 4813 10557 4847 10591
rect 6193 10557 6227 10591
rect 7573 10557 7607 10591
rect 14841 10557 14875 10591
rect 16129 10557 16163 10591
rect 22569 10557 22603 10591
rect 6745 10489 6779 10523
rect 2145 10421 2179 10455
rect 4077 10421 4111 10455
rect 10977 10421 11011 10455
rect 12173 10421 12207 10455
rect 14289 10421 14323 10455
rect 15853 10421 15887 10455
rect 16313 10421 16347 10455
rect 17049 10421 17083 10455
rect 19809 10421 19843 10455
rect 1764 10217 1798 10251
rect 3249 10217 3283 10251
rect 5168 10217 5202 10251
rect 6653 10217 6687 10251
rect 15577 10217 15611 10251
rect 15945 10217 15979 10251
rect 16497 10217 16531 10251
rect 18521 10217 18555 10251
rect 23489 10217 23523 10251
rect 18889 10149 18923 10183
rect 1501 10081 1535 10115
rect 4537 10081 4571 10115
rect 4905 10081 4939 10115
rect 9413 10081 9447 10115
rect 9689 10081 9723 10115
rect 11253 10081 11287 10115
rect 18153 10081 18187 10115
rect 20913 10081 20947 10115
rect 7481 10013 7515 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 8033 10013 8067 10047
rect 13093 10013 13127 10047
rect 13277 10013 13311 10047
rect 15393 10013 15427 10047
rect 16037 10013 16071 10047
rect 16221 10013 16255 10047
rect 16865 10013 16899 10047
rect 18337 10013 18371 10047
rect 18613 10013 18647 10047
rect 18705 10013 18739 10047
rect 19809 10013 19843 10047
rect 19993 10013 20027 10047
rect 20177 10013 20211 10047
rect 23213 10013 23247 10047
rect 24593 10013 24627 10047
rect 24866 9991 24900 10025
rect 25513 10013 25547 10047
rect 11529 9945 11563 9979
rect 16451 9945 16485 9979
rect 18889 9945 18923 9979
rect 19257 9945 19291 9979
rect 21189 9945 21223 9979
rect 22937 9945 22971 9979
rect 23305 9945 23339 9979
rect 3985 9877 4019 9911
rect 7297 9877 7331 9911
rect 7665 9877 7699 9911
rect 7941 9877 7975 9911
rect 11161 9877 11195 9911
rect 13001 9877 13035 9911
rect 13185 9877 13219 9911
rect 15209 9877 15243 9911
rect 20085 9877 20119 9911
rect 23029 9877 23063 9911
rect 23505 9877 23539 9911
rect 23673 9877 23707 9911
rect 24409 9877 24443 9911
rect 24777 9877 24811 9911
rect 25329 9877 25363 9911
rect 8033 9673 8067 9707
rect 13829 9673 13863 9707
rect 21097 9673 21131 9707
rect 25237 9673 25271 9707
rect 11161 9605 11195 9639
rect 15761 9605 15795 9639
rect 22845 9605 22879 9639
rect 25329 9605 25363 9639
rect 3525 9537 3559 9571
rect 7573 9537 7607 9571
rect 8125 9537 8159 9571
rect 10057 9537 10091 9571
rect 10425 9537 10459 9571
rect 11529 9537 11563 9571
rect 13888 9537 13922 9571
rect 15853 9537 15887 9571
rect 20821 9537 20855 9571
rect 21005 9537 21039 9571
rect 21281 9537 21315 9571
rect 22017 9537 22051 9571
rect 24777 9537 24811 9571
rect 24869 9537 24903 9571
rect 3801 9469 3835 9503
rect 7389 9469 7423 9503
rect 9689 9469 9723 9503
rect 11805 9469 11839 9503
rect 13369 9469 13403 9503
rect 15945 9469 15979 9503
rect 17601 9469 17635 9503
rect 17877 9469 17911 9503
rect 19625 9469 19659 9503
rect 20913 9469 20947 9503
rect 21557 9469 21591 9503
rect 22201 9469 22235 9503
rect 22569 9469 22603 9503
rect 24685 9469 24719 9503
rect 25881 9469 25915 9503
rect 5273 9401 5307 9435
rect 13277 9401 13311 9435
rect 14013 9401 14047 9435
rect 15393 9401 15427 9435
rect 7757 9333 7791 9367
rect 8263 9333 8297 9367
rect 13461 9333 13495 9367
rect 21465 9333 21499 9367
rect 21833 9333 21867 9367
rect 24317 9333 24351 9367
rect 3985 9129 4019 9163
rect 10149 9129 10183 9163
rect 12449 9129 12483 9163
rect 15485 9129 15519 9163
rect 18797 9129 18831 9163
rect 22155 9129 22189 9163
rect 23305 9129 23339 9163
rect 8033 9061 8067 9095
rect 23213 9061 23247 9095
rect 7205 8993 7239 9027
rect 8125 8993 8159 9027
rect 10793 8993 10827 9027
rect 14197 8993 14231 9027
rect 14381 8993 14415 9027
rect 16129 8993 16163 9027
rect 22661 8993 22695 9027
rect 23949 8993 23983 9027
rect 24685 8993 24719 9027
rect 3525 8925 3559 8959
rect 4445 8925 4479 8959
rect 4537 8925 4571 8959
rect 4629 8925 4663 8959
rect 4813 8925 4847 8959
rect 6469 8925 6503 8959
rect 6745 8925 6779 8959
rect 7481 8925 7515 8959
rect 7849 8925 7883 8959
rect 8677 8925 8711 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 9413 8925 9447 8959
rect 9505 8925 9539 8959
rect 11069 8925 11103 8959
rect 11253 8925 11287 8959
rect 12081 8925 12115 8959
rect 13277 8925 13311 8959
rect 15853 8925 15887 8959
rect 18705 8925 18739 8959
rect 18797 8925 18831 8959
rect 18981 8925 19015 8959
rect 20361 8925 20395 8959
rect 20729 8925 20763 8959
rect 22937 8925 22971 8959
rect 23029 8925 23063 8959
rect 23673 8925 23707 8959
rect 24409 8925 24443 8959
rect 3953 8857 3987 8891
rect 4169 8857 4203 8891
rect 6193 8857 6227 8891
rect 7665 8857 7699 8891
rect 7757 8857 7791 8891
rect 9045 8857 9079 8891
rect 12633 8857 12667 8891
rect 17877 8857 17911 8891
rect 2973 8789 3007 8823
rect 3801 8789 3835 8823
rect 4261 8789 4295 8823
rect 10241 8789 10275 8823
rect 11437 8789 11471 8823
rect 11529 8789 11563 8823
rect 12265 8789 12299 8823
rect 12433 8789 12467 8823
rect 12725 8789 12759 8823
rect 14473 8789 14507 8823
rect 14841 8789 14875 8823
rect 15945 8789 15979 8823
rect 22845 8789 22879 8823
rect 23765 8789 23799 8823
rect 26157 8789 26191 8823
rect 4353 8585 4387 8619
rect 7941 8585 7975 8619
rect 10977 8585 11011 8619
rect 11989 8585 12023 8619
rect 13277 8585 13311 8619
rect 14933 8585 14967 8619
rect 19993 8585 20027 8619
rect 25605 8585 25639 8619
rect 4103 8517 4137 8551
rect 5457 8517 5491 8551
rect 6193 8517 6227 8551
rect 7297 8517 7331 8551
rect 11621 8517 11655 8551
rect 15853 8517 15887 8551
rect 16037 8517 16071 8551
rect 20913 8517 20947 8551
rect 23581 8517 23615 8551
rect 24133 8517 24167 8551
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 3985 8449 4019 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 7849 8449 7883 8483
rect 9689 8449 9723 8483
rect 10885 8449 10919 8483
rect 11161 8449 11195 8483
rect 11897 8449 11931 8483
rect 12173 8449 12207 8483
rect 12265 8449 12299 8483
rect 12449 8449 12483 8483
rect 12633 8455 12667 8489
rect 12725 8439 12759 8473
rect 13093 8449 13127 8483
rect 15117 8449 15151 8483
rect 15209 8449 15243 8483
rect 15393 8449 15427 8483
rect 15485 8449 15519 8483
rect 16129 8449 16163 8483
rect 16313 8449 16347 8483
rect 16681 8449 16715 8483
rect 17233 8449 17267 8483
rect 19993 8449 20027 8483
rect 20361 8449 20395 8483
rect 20821 8449 20855 8483
rect 21005 8449 21039 8483
rect 21833 8449 21867 8483
rect 22937 8449 22971 8483
rect 23121 8449 23155 8483
rect 23213 8449 23247 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 4261 8381 4295 8415
rect 4997 8381 5031 8415
rect 6561 8381 6595 8415
rect 9413 8381 9447 8415
rect 10793 8381 10827 8415
rect 11345 8381 11379 8415
rect 11805 8381 11839 8415
rect 19717 8381 19751 8415
rect 22385 8381 22419 8415
rect 23857 8381 23891 8415
rect 3617 8313 3651 8347
rect 11897 8313 11931 8347
rect 12357 8313 12391 8347
rect 19901 8313 19935 8347
rect 20545 8313 20579 8347
rect 23029 8313 23063 8347
rect 3157 8245 3191 8279
rect 7389 8245 7423 8279
rect 12817 8245 12851 8279
rect 15669 8245 15703 8279
rect 16221 8245 16255 8279
rect 23581 8245 23615 8279
rect 23765 8245 23799 8279
rect 3985 8041 4019 8075
rect 23305 8041 23339 8075
rect 23581 8041 23615 8075
rect 10057 7973 10091 8007
rect 14841 7973 14875 8007
rect 2145 7905 2179 7939
rect 4077 7905 4111 7939
rect 4813 7905 4847 7939
rect 6745 7905 6779 7939
rect 8769 7905 8803 7939
rect 10701 7905 10735 7939
rect 15485 7905 15519 7939
rect 19901 7905 19935 7939
rect 20637 7905 20671 7939
rect 24041 7905 24075 7939
rect 1869 7837 1903 7871
rect 3801 7837 3835 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 5181 7837 5215 7871
rect 11897 7837 11931 7871
rect 12633 7837 12667 7871
rect 13001 7837 13035 7871
rect 14657 7837 14691 7871
rect 15025 7837 15059 7871
rect 15301 7837 15335 7871
rect 15393 7837 15427 7871
rect 18797 7837 18831 7871
rect 18981 7837 19015 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 23029 7837 23063 7871
rect 23213 7837 23247 7871
rect 23397 7837 23431 7871
rect 23765 7837 23799 7871
rect 23857 7837 23891 7871
rect 23949 7837 23983 7871
rect 7021 7769 7055 7803
rect 11161 7769 11195 7803
rect 15117 7769 15151 7803
rect 15761 7769 15795 7803
rect 20913 7769 20947 7803
rect 3617 7701 3651 7735
rect 6607 7701 6641 7735
rect 12081 7701 12115 7735
rect 12817 7701 12851 7735
rect 14565 7701 14599 7735
rect 15215 7701 15249 7735
rect 17233 7701 17267 7735
rect 18889 7701 18923 7735
rect 19257 7701 19291 7735
rect 20545 7701 20579 7735
rect 22385 7701 22419 7735
rect 22477 7701 22511 7735
rect 2145 7497 2179 7531
rect 3065 7497 3099 7531
rect 10609 7497 10643 7531
rect 11989 7497 12023 7531
rect 16083 7497 16117 7531
rect 17601 7497 17635 7531
rect 19625 7497 19659 7531
rect 20361 7497 20395 7531
rect 20729 7497 20763 7531
rect 20821 7497 20855 7531
rect 23305 7497 23339 7531
rect 24317 7497 24351 7531
rect 3893 7429 3927 7463
rect 4445 7429 4479 7463
rect 12725 7429 12759 7463
rect 20085 7429 20119 7463
rect 24133 7429 24167 7463
rect 24409 7429 24443 7463
rect 2329 7361 2363 7395
rect 3157 7361 3191 7395
rect 4169 7361 4203 7395
rect 6009 7361 6043 7395
rect 6193 7361 6227 7395
rect 7389 7361 7423 7395
rect 10517 7361 10551 7395
rect 12081 7361 12115 7395
rect 17233 7361 17267 7395
rect 19901 7361 19935 7395
rect 20177 7361 20211 7395
rect 21189 7361 21223 7395
rect 21373 7361 21407 7395
rect 22937 7361 22971 7395
rect 23213 7361 23247 7395
rect 23397 7361 23431 7395
rect 23673 7361 23707 7395
rect 23857 7361 23891 7395
rect 23949 7361 23983 7395
rect 24593 7361 24627 7395
rect 24777 7361 24811 7395
rect 25053 7361 25087 7395
rect 25237 7361 25271 7395
rect 3341 7293 3375 7327
rect 6101 7293 6135 7327
rect 7941 7293 7975 7327
rect 10057 7293 10091 7327
rect 10333 7293 10367 7327
rect 12265 7293 12299 7327
rect 12449 7293 12483 7327
rect 14289 7293 14323 7327
rect 14657 7293 14691 7327
rect 17877 7293 17911 7327
rect 18153 7293 18187 7327
rect 19717 7293 19751 7327
rect 21005 7293 21039 7327
rect 22753 7293 22787 7327
rect 2697 7225 2731 7259
rect 17785 7225 17819 7259
rect 23121 7225 23155 7259
rect 3617 7157 3651 7191
rect 5917 7157 5951 7191
rect 8585 7157 8619 7191
rect 11621 7157 11655 7191
rect 14197 7157 14231 7191
rect 17601 7157 17635 7191
rect 21557 7157 21591 7191
rect 23857 7157 23891 7191
rect 24869 7157 24903 7191
rect 25053 7157 25087 7191
rect 10504 6953 10538 6987
rect 11989 6953 12023 6987
rect 16129 6953 16163 6987
rect 23305 6953 23339 6987
rect 23765 6953 23799 6987
rect 26157 6953 26191 6987
rect 3801 6885 3835 6919
rect 4721 6885 4755 6919
rect 8033 6885 8067 6919
rect 15669 6885 15703 6919
rect 23489 6885 23523 6919
rect 23857 6885 23891 6919
rect 3249 6817 3283 6851
rect 5733 6817 5767 6851
rect 9505 6817 9539 6851
rect 10241 6817 10275 6851
rect 12081 6817 12115 6851
rect 14657 6817 14691 6851
rect 14933 6817 14967 6851
rect 19073 6817 19107 6851
rect 19993 6817 20027 6851
rect 20177 6817 20211 6851
rect 21557 6817 21591 6851
rect 22109 6817 22143 6851
rect 23121 6817 23155 6851
rect 23949 6817 23983 6851
rect 4353 6749 4387 6783
rect 4556 6749 4590 6783
rect 4688 6749 4722 6783
rect 4997 6749 5031 6783
rect 5365 6749 5399 6783
rect 5549 6749 5583 6783
rect 7849 6749 7883 6783
rect 8217 6749 8251 6783
rect 14565 6749 14599 6783
rect 15577 6749 15611 6783
rect 16037 6749 16071 6783
rect 16221 6749 16255 6783
rect 17325 6749 17359 6783
rect 21649 6749 21683 6783
rect 21925 6749 21959 6783
rect 23397 6749 23431 6783
rect 24225 6749 24259 6783
rect 24409 6749 24443 6783
rect 3433 6681 3467 6715
rect 3617 6681 3651 6715
rect 8769 6681 8803 6715
rect 9321 6681 9355 6715
rect 12357 6681 12391 6715
rect 15853 6681 15887 6715
rect 17601 6681 17635 6715
rect 20913 6681 20947 6715
rect 24685 6681 24719 6715
rect 8953 6613 8987 6647
rect 9413 6613 9447 6647
rect 13829 6613 13863 6647
rect 14105 6613 14139 6647
rect 14473 6613 14507 6647
rect 19441 6613 19475 6647
rect 20821 6613 20855 6647
rect 21741 6613 21775 6647
rect 22845 6613 22879 6647
rect 24133 6613 24167 6647
rect 3157 6409 3191 6443
rect 3617 6409 3651 6443
rect 4169 6409 4203 6443
rect 4353 6409 4387 6443
rect 5917 6409 5951 6443
rect 6009 6409 6043 6443
rect 8861 6409 8895 6443
rect 10701 6409 10735 6443
rect 11161 6409 11195 6443
rect 14841 6409 14875 6443
rect 18889 6409 18923 6443
rect 21189 6409 21223 6443
rect 21833 6409 21867 6443
rect 22569 6409 22603 6443
rect 24225 6409 24259 6443
rect 4721 6341 4755 6375
rect 4997 6341 5031 6375
rect 19717 6341 19751 6375
rect 21373 6341 21407 6375
rect 24593 6341 24627 6375
rect 25513 6341 25547 6375
rect 4491 6307 4525 6341
rect 3433 6273 3467 6307
rect 3709 6273 3743 6307
rect 4077 6273 4111 6307
rect 4261 6273 4295 6307
rect 4813 6273 4847 6307
rect 5457 6273 5491 6307
rect 5733 6273 5767 6307
rect 6009 6273 6043 6307
rect 6193 6273 6227 6307
rect 6377 6273 6411 6307
rect 11345 6273 11379 6307
rect 11529 6273 11563 6307
rect 14197 6273 14231 6307
rect 19349 6273 19383 6307
rect 19441 6273 19475 6307
rect 21557 6273 21591 6307
rect 21649 6273 21683 6307
rect 22753 6273 22787 6307
rect 22845 6273 22879 6307
rect 23029 6273 23063 6307
rect 23121 6273 23155 6307
rect 23489 6273 23523 6307
rect 23765 6273 23799 6307
rect 24409 6273 24443 6307
rect 24501 6273 24535 6307
rect 24777 6273 24811 6307
rect 25237 6273 25271 6307
rect 26065 6273 26099 6307
rect 1409 6205 1443 6239
rect 1685 6205 1719 6239
rect 3249 6205 3283 6239
rect 5181 6205 5215 6239
rect 5549 6205 5583 6239
rect 7113 6205 7147 6239
rect 7389 6205 7423 6239
rect 8953 6205 8987 6239
rect 9229 6205 9263 6239
rect 11805 6205 11839 6239
rect 13921 6205 13955 6239
rect 16221 6205 16255 6239
rect 22385 6205 22419 6239
rect 24869 6205 24903 6239
rect 25145 6205 25179 6239
rect 21649 6137 21683 6171
rect 4537 6069 4571 6103
rect 5733 6069 5767 6103
rect 6561 6069 6595 6103
rect 13277 6069 13311 6103
rect 13369 6069 13403 6103
rect 15577 6069 15611 6103
rect 19257 6069 19291 6103
rect 23213 6069 23247 6103
rect 23489 6069 23523 6103
rect 3433 5865 3467 5899
rect 3801 5865 3835 5899
rect 3985 5865 4019 5899
rect 5457 5865 5491 5899
rect 5825 5865 5859 5899
rect 9873 5865 9907 5899
rect 11621 5865 11655 5899
rect 21741 5865 21775 5899
rect 22753 5865 22787 5899
rect 24961 5865 24995 5899
rect 13461 5797 13495 5831
rect 14657 5797 14691 5831
rect 21373 5797 21407 5831
rect 21925 5797 21959 5831
rect 23121 5797 23155 5831
rect 6101 5729 6135 5763
rect 8401 5729 8435 5763
rect 19625 5729 19659 5763
rect 24777 5729 24811 5763
rect 3157 5661 3191 5695
rect 5089 5661 5123 5695
rect 5457 5661 5491 5695
rect 5641 5661 5675 5695
rect 6193 5661 6227 5695
rect 9505 5661 9539 5695
rect 9689 5661 9723 5695
rect 9873 5661 9907 5695
rect 11437 5661 11471 5695
rect 11897 5661 11931 5695
rect 12081 5661 12115 5695
rect 13645 5661 13679 5695
rect 14197 5661 14231 5695
rect 17233 5661 17267 5695
rect 17417 5661 17451 5695
rect 17509 5661 17543 5695
rect 21465 5661 21499 5695
rect 22753 5661 22787 5695
rect 22937 5661 22971 5695
rect 23213 5661 23247 5695
rect 25053 5661 25087 5695
rect 3249 5593 3283 5627
rect 3465 5593 3499 5627
rect 4169 5593 4203 5627
rect 8125 5593 8159 5627
rect 8953 5593 8987 5627
rect 12265 5593 12299 5627
rect 16957 5593 16991 5627
rect 19901 5593 19935 5627
rect 3065 5525 3099 5559
rect 3617 5525 3651 5559
rect 3959 5525 3993 5559
rect 5273 5525 5307 5559
rect 6653 5525 6687 5559
rect 14381 5525 14415 5559
rect 15485 5525 15519 5559
rect 17693 5525 17727 5559
rect 23397 5525 23431 5559
rect 24501 5525 24535 5559
rect 3157 5321 3191 5355
rect 4353 5321 4387 5355
rect 5641 5321 5675 5355
rect 8309 5321 8343 5355
rect 14933 5321 14967 5355
rect 16681 5321 16715 5355
rect 19993 5321 20027 5355
rect 22569 5321 22603 5355
rect 24317 5321 24351 5355
rect 3985 5253 4019 5287
rect 12357 5253 12391 5287
rect 16497 5253 16531 5287
rect 17049 5253 17083 5287
rect 17601 5253 17635 5287
rect 22109 5253 22143 5287
rect 22201 5253 22235 5287
rect 24225 5253 24259 5287
rect 24501 5253 24535 5287
rect 1409 5185 1443 5219
rect 3617 5185 3651 5219
rect 4261 5185 4295 5219
rect 5089 5185 5123 5219
rect 7113 5185 7147 5219
rect 7941 5185 7975 5219
rect 8125 5185 8159 5219
rect 8769 5185 8803 5219
rect 12541 5185 12575 5219
rect 12633 5185 12667 5219
rect 12725 5185 12759 5219
rect 13369 5185 13403 5219
rect 13461 5185 13495 5219
rect 13645 5185 13679 5219
rect 15117 5185 15151 5219
rect 15209 5185 15243 5219
rect 15393 5185 15427 5219
rect 15485 5185 15519 5219
rect 15577 5185 15611 5219
rect 15761 5185 15795 5219
rect 16865 5185 16899 5219
rect 17141 5185 17175 5219
rect 20177 5185 20211 5219
rect 22017 5185 22051 5219
rect 22319 5185 22353 5219
rect 22753 5185 22787 5219
rect 22937 5185 22971 5219
rect 23029 5185 23063 5219
rect 23213 5185 23247 5219
rect 24133 5185 24167 5219
rect 1685 5117 1719 5151
rect 3525 5117 3559 5151
rect 3893 5117 3927 5151
rect 5365 5117 5399 5151
rect 7757 5117 7791 5151
rect 7849 5117 7883 5151
rect 13001 5117 13035 5151
rect 15945 5117 15979 5151
rect 17325 5117 17359 5151
rect 22477 5117 22511 5151
rect 3341 5049 3375 5083
rect 8585 5049 8619 5083
rect 5181 4981 5215 5015
rect 12633 4981 12667 5015
rect 13001 4981 13035 5015
rect 13277 4981 13311 5015
rect 13829 4981 13863 5015
rect 15669 4981 15703 5015
rect 19073 4981 19107 5015
rect 21833 4981 21867 5015
rect 23397 4981 23431 5015
rect 23949 4981 23983 5015
rect 26157 4981 26191 5015
rect 2789 4777 2823 4811
rect 4445 4777 4479 4811
rect 4905 4777 4939 4811
rect 5641 4777 5675 4811
rect 9689 4777 9723 4811
rect 10057 4777 10091 4811
rect 13645 4777 13679 4811
rect 14749 4777 14783 4811
rect 15669 4777 15703 4811
rect 15853 4777 15887 4811
rect 16129 4777 16163 4811
rect 17417 4777 17451 4811
rect 22845 4777 22879 4811
rect 3341 4709 3375 4743
rect 16313 4709 16347 4743
rect 17785 4709 17819 4743
rect 17969 4709 18003 4743
rect 2881 4641 2915 4675
rect 3801 4641 3835 4675
rect 7573 4641 7607 4675
rect 7665 4641 7699 4675
rect 8677 4641 8711 4675
rect 12817 4641 12851 4675
rect 13001 4641 13035 4675
rect 16957 4641 16991 4675
rect 17325 4641 17359 4675
rect 17877 4641 17911 4675
rect 20637 4641 20671 4675
rect 22661 4641 22695 4675
rect 25237 4641 25271 4675
rect 2605 4573 2639 4607
rect 2697 4573 2731 4607
rect 2973 4573 3007 4607
rect 3157 4573 3191 4607
rect 3985 4573 4019 4607
rect 4169 4573 4203 4607
rect 5089 4573 5123 4607
rect 5273 4573 5307 4607
rect 5549 4573 5583 4607
rect 6009 4573 6043 4607
rect 6653 4573 6687 4607
rect 7297 4573 7331 4607
rect 7757 4573 7791 4607
rect 7849 4573 7883 4607
rect 8493 4573 8527 4607
rect 8953 4573 8987 4607
rect 9873 4573 9907 4607
rect 10057 4573 10091 4607
rect 13185 4573 13219 4607
rect 13277 4573 13311 4607
rect 13461 4573 13495 4607
rect 13737 4573 13771 4607
rect 13921 4573 13955 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 14381 4573 14415 4607
rect 14493 4573 14527 4607
rect 15117 4573 15151 4607
rect 15209 4573 15243 4607
rect 15393 4573 15427 4607
rect 15945 4573 15979 4607
rect 16037 4573 16071 4607
rect 16405 4573 16439 4607
rect 16865 4573 16899 4607
rect 17049 4573 17083 4607
rect 17141 4573 17175 4607
rect 17601 4573 17635 4607
rect 18153 4573 18187 4607
rect 18429 4573 18463 4607
rect 19441 4573 19475 4607
rect 19533 4573 19567 4607
rect 19809 4573 19843 4607
rect 22753 4575 22787 4609
rect 22937 4573 22971 4607
rect 23305 4573 23339 4607
rect 23581 4573 23615 4607
rect 25329 4573 25363 4607
rect 4629 4505 4663 4539
rect 5181 4505 5215 4539
rect 5411 4505 5445 4539
rect 5825 4505 5859 4539
rect 7205 4505 7239 4539
rect 8401 4505 8435 4539
rect 9597 4505 9631 4539
rect 12725 4505 12759 4539
rect 14841 4505 14875 4539
rect 15485 4505 15519 4539
rect 16313 4505 16347 4539
rect 18521 4505 18555 4539
rect 18705 4505 18739 4539
rect 19901 4505 19935 4539
rect 20913 4505 20947 4539
rect 4261 4437 4295 4471
rect 4429 4437 4463 4471
rect 6101 4437 6135 4471
rect 7389 4437 7423 4471
rect 8033 4437 8067 4471
rect 12357 4437 12391 4471
rect 13737 4437 13771 4471
rect 15025 4437 15059 4471
rect 15690 4437 15724 4471
rect 16497 4437 16531 4471
rect 18337 4437 18371 4471
rect 18889 4437 18923 4471
rect 19349 4437 19383 4471
rect 19625 4437 19659 4471
rect 23121 4437 23155 4471
rect 23489 4437 23523 4471
rect 24593 4437 24627 4471
rect 25421 4437 25455 4471
rect 3065 4233 3099 4267
rect 5733 4233 5767 4267
rect 6101 4233 6135 4267
rect 6377 4233 6411 4267
rect 7481 4233 7515 4267
rect 8309 4233 8343 4267
rect 10517 4233 10551 4267
rect 17325 4233 17359 4267
rect 19717 4233 19751 4267
rect 22293 4233 22327 4267
rect 25513 4233 25547 4267
rect 4011 4165 4045 4199
rect 5273 4165 5307 4199
rect 9781 4165 9815 4199
rect 14355 4165 14389 4199
rect 14473 4165 14507 4199
rect 14565 4165 14599 4199
rect 17785 4165 17819 4199
rect 19901 4165 19935 4199
rect 22201 4165 22235 4199
rect 22937 4165 22971 4199
rect 23029 4165 23063 4199
rect 23489 4165 23523 4199
rect 3157 4097 3191 4131
rect 3710 4087 3744 4121
rect 3802 4097 3836 4131
rect 3893 4097 3927 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 5483 4097 5517 4131
rect 5917 4097 5951 4131
rect 6193 4097 6227 4131
rect 6652 4119 6686 4153
rect 7665 4097 7699 4131
rect 10333 4097 10367 4131
rect 10609 4097 10643 4131
rect 10701 4097 10735 4131
rect 10885 4097 10919 4131
rect 14657 4097 14691 4131
rect 16313 4097 16347 4131
rect 16681 4097 16715 4131
rect 16865 4097 16899 4131
rect 16957 4097 16991 4131
rect 17509 4097 17543 4131
rect 17601 4097 17635 4131
rect 18061 4097 18095 4131
rect 18337 4097 18371 4131
rect 19809 4097 19843 4131
rect 20361 4097 20395 4131
rect 22862 4087 22896 4121
rect 23147 4097 23181 4131
rect 23397 4097 23431 4131
rect 23673 4097 23707 4131
rect 23765 4097 23799 4131
rect 3249 4029 3283 4063
rect 4169 4029 4203 4063
rect 4261 4029 4295 4063
rect 4813 4029 4847 4063
rect 5641 4029 5675 4063
rect 6377 4029 6411 4063
rect 6837 4029 6871 4063
rect 10057 4029 10091 4063
rect 10793 4029 10827 4063
rect 11529 4029 11563 4063
rect 13277 4029 13311 4063
rect 13553 4029 13587 4063
rect 14197 4029 14231 4063
rect 14841 4029 14875 4063
rect 15485 4029 15519 4063
rect 15853 4029 15887 4063
rect 15945 4029 15979 4063
rect 16037 4029 16071 4063
rect 16129 4029 16163 4063
rect 18245 4029 18279 4063
rect 19349 4029 19383 4063
rect 19533 4029 19567 4063
rect 22477 4029 22511 4063
rect 23305 4029 23339 4063
rect 24041 4029 24075 4063
rect 14933 3961 14967 3995
rect 18153 3961 18187 3995
rect 23397 3961 23431 3995
rect 2697 3893 2731 3927
rect 3525 3893 3559 3927
rect 4997 3893 5031 3927
rect 6561 3893 6595 3927
rect 8217 3893 8251 3927
rect 10149 3893 10183 3927
rect 15669 3893 15703 3927
rect 16405 3893 16439 3927
rect 16681 3893 16715 3927
rect 17141 3893 17175 3927
rect 17785 3893 17819 3927
rect 18521 3893 18555 3927
rect 18797 3893 18831 3927
rect 20085 3893 20119 3927
rect 20177 3893 20211 3927
rect 21833 3893 21867 3927
rect 22661 3893 22695 3927
rect 3249 3689 3283 3723
rect 4169 3689 4203 3723
rect 4984 3689 5018 3723
rect 6469 3689 6503 3723
rect 8769 3689 8803 3723
rect 16313 3689 16347 3723
rect 19993 3689 20027 3723
rect 24225 3689 24259 3723
rect 13921 3621 13955 3655
rect 24409 3621 24443 3655
rect 7021 3553 7055 3587
rect 9137 3553 9171 3587
rect 10701 3553 10735 3587
rect 12725 3553 12759 3587
rect 14565 3553 14599 3587
rect 16957 3553 16991 3587
rect 17325 3553 17359 3587
rect 19349 3553 19383 3587
rect 20637 3553 20671 3587
rect 20913 3553 20947 3587
rect 22661 3553 22695 3587
rect 23581 3553 23615 3587
rect 24961 3553 24995 3587
rect 25605 3553 25639 3587
rect 1501 3485 1535 3519
rect 4353 3485 4387 3519
rect 4629 3485 4663 3519
rect 4721 3485 4755 3519
rect 10425 3485 10459 3519
rect 13185 3485 13219 3519
rect 13277 3485 13311 3519
rect 19533 3485 19567 3519
rect 19625 3485 19659 3519
rect 23719 3485 23753 3519
rect 23857 3485 23891 3519
rect 24041 3485 24075 3519
rect 25329 3485 25363 3519
rect 25421 3485 25455 3519
rect 25513 3485 25547 3519
rect 1777 3417 1811 3451
rect 7297 3417 7331 3451
rect 9873 3417 9907 3451
rect 10977 3417 11011 3451
rect 13001 3417 13035 3451
rect 14105 3417 14139 3451
rect 14289 3417 14323 3451
rect 14841 3417 14875 3451
rect 17601 3417 17635 3451
rect 23949 3417 23983 3451
rect 4537 3349 4571 3383
rect 9781 3349 9815 3383
rect 12817 3349 12851 3383
rect 14473 3349 14507 3383
rect 16405 3349 16439 3383
rect 19073 3349 19107 3383
rect 25145 3349 25179 3383
rect 2145 3145 2179 3179
rect 4537 3145 4571 3179
rect 4905 3145 4939 3179
rect 6377 3145 6411 3179
rect 8217 3145 8251 3179
rect 8585 3145 8619 3179
rect 10701 3145 10735 3179
rect 11161 3145 11195 3179
rect 14289 3145 14323 3179
rect 16681 3145 16715 3179
rect 17785 3145 17819 3179
rect 21281 3145 21315 3179
rect 3065 3077 3099 3111
rect 7849 3077 7883 3111
rect 13967 3077 14001 3111
rect 15025 3077 15059 3111
rect 15143 3077 15177 3111
rect 20085 3077 20119 3111
rect 22477 3077 22511 3111
rect 24225 3077 24259 3111
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 4721 3009 4755 3043
rect 4905 3009 4939 3043
rect 8125 3009 8159 3043
rect 8401 3009 8435 3043
rect 8677 3009 8711 3043
rect 8769 3009 8803 3043
rect 10609 3009 10643 3043
rect 11345 3009 11379 3043
rect 11529 3009 11563 3043
rect 13645 3009 13679 3043
rect 13737 3009 13771 3043
rect 13829 3009 13863 3043
rect 14105 3009 14139 3043
rect 14381 3009 14415 3043
rect 14841 3009 14875 3043
rect 14933 3009 14967 3043
rect 15301 3009 15335 3043
rect 15853 3009 15887 3043
rect 16037 3009 16071 3043
rect 17049 3009 17083 3043
rect 17141 3009 17175 3043
rect 20361 3009 20395 3043
rect 21465 3009 21499 3043
rect 9045 2941 9079 2975
rect 10517 2941 10551 2975
rect 11805 2941 11839 2975
rect 13461 2941 13495 2975
rect 16957 2941 16991 2975
rect 18337 2941 18371 2975
rect 22201 2941 22235 2975
rect 13277 2873 13311 2907
rect 14657 2873 14691 2907
rect 18613 2873 18647 2907
rect 16037 2805 16071 2839
rect 17049 2805 17083 2839
rect 17325 2805 17359 2839
rect 9137 2601 9171 2635
rect 14565 2601 14599 2635
rect 17877 2601 17911 2635
rect 14381 2533 14415 2567
rect 9781 2465 9815 2499
rect 18521 2465 18555 2499
rect 10425 2397 10459 2431
rect 14105 2397 14139 2431
rect 18061 2397 18095 2431
rect 18153 2397 18187 2431
rect 18245 2397 18279 2431
rect 25789 2397 25823 2431
rect 18363 2329 18397 2363
rect 18705 2329 18739 2363
rect 26157 2329 26191 2363
rect 18797 2261 18831 2295
<< metal1 >>
rect 1104 27226 26656 27248
rect 1104 27174 7298 27226
rect 7350 27174 7362 27226
rect 7414 27174 7426 27226
rect 7478 27174 7490 27226
rect 7542 27174 7554 27226
rect 7606 27174 13646 27226
rect 13698 27174 13710 27226
rect 13762 27174 13774 27226
rect 13826 27174 13838 27226
rect 13890 27174 13902 27226
rect 13954 27174 19994 27226
rect 20046 27174 20058 27226
rect 20110 27174 20122 27226
rect 20174 27174 20186 27226
rect 20238 27174 20250 27226
rect 20302 27174 26342 27226
rect 26394 27174 26406 27226
rect 26458 27174 26470 27226
rect 26522 27174 26534 27226
rect 26586 27174 26598 27226
rect 26650 27174 26656 27226
rect 1104 27152 26656 27174
rect 20901 27115 20959 27121
rect 20901 27081 20913 27115
rect 20947 27112 20959 27115
rect 21174 27112 21180 27124
rect 20947 27084 21180 27112
rect 20947 27081 20959 27084
rect 20901 27075 20959 27081
rect 21174 27072 21180 27084
rect 21232 27072 21238 27124
rect 16761 27047 16819 27053
rect 16761 27013 16773 27047
rect 16807 27044 16819 27047
rect 17494 27044 17500 27056
rect 16807 27016 17500 27044
rect 16807 27013 16819 27016
rect 16761 27007 16819 27013
rect 17494 27004 17500 27016
rect 17552 27004 17558 27056
rect 21821 27047 21879 27053
rect 21821 27044 21833 27047
rect 21192 27016 21833 27044
rect 3878 26936 3884 26988
rect 3936 26976 3942 26988
rect 3973 26979 4031 26985
rect 3973 26976 3985 26979
rect 3936 26948 3985 26976
rect 3936 26936 3942 26948
rect 3973 26945 3985 26948
rect 4019 26945 4031 26979
rect 3973 26939 4031 26945
rect 11054 26936 11060 26988
rect 11112 26936 11118 26988
rect 14826 26936 14832 26988
rect 14884 26976 14890 26988
rect 14921 26979 14979 26985
rect 14921 26976 14933 26979
rect 14884 26948 14933 26976
rect 14884 26936 14890 26948
rect 14921 26945 14933 26948
rect 14967 26945 14979 26979
rect 14921 26939 14979 26945
rect 16574 26936 16580 26988
rect 16632 26976 16638 26988
rect 16669 26979 16727 26985
rect 16669 26976 16681 26979
rect 16632 26948 16681 26976
rect 16632 26936 16638 26948
rect 16669 26945 16681 26948
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 16945 26979 17003 26985
rect 16945 26945 16957 26979
rect 16991 26976 17003 26979
rect 17218 26976 17224 26988
rect 16991 26948 17224 26976
rect 16991 26945 17003 26948
rect 16945 26939 17003 26945
rect 17218 26936 17224 26948
rect 17276 26936 17282 26988
rect 20809 26979 20867 26985
rect 20809 26945 20821 26979
rect 20855 26976 20867 26979
rect 21082 26976 21088 26988
rect 20855 26948 21088 26976
rect 20855 26945 20867 26948
rect 20809 26939 20867 26945
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 21192 26985 21220 27016
rect 21821 27013 21833 27016
rect 21867 27013 21879 27047
rect 21821 27007 21879 27013
rect 21177 26979 21235 26985
rect 21177 26945 21189 26979
rect 21223 26945 21235 26979
rect 21177 26939 21235 26945
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26976 21327 26979
rect 21315 26948 21496 26976
rect 21315 26945 21327 26948
rect 21269 26939 21327 26945
rect 21468 26920 21496 26948
rect 934 26868 940 26920
rect 992 26908 998 26920
rect 1397 26911 1455 26917
rect 1397 26908 1409 26911
rect 992 26880 1409 26908
rect 992 26868 998 26880
rect 1397 26877 1409 26880
rect 1443 26877 1455 26911
rect 1397 26871 1455 26877
rect 20990 26868 20996 26920
rect 21048 26868 21054 26920
rect 21450 26868 21456 26920
rect 21508 26868 21514 26920
rect 21545 26911 21603 26917
rect 21545 26877 21557 26911
rect 21591 26908 21603 26911
rect 21634 26908 21640 26920
rect 21591 26880 21640 26908
rect 21591 26877 21603 26880
rect 21545 26871 21603 26877
rect 21634 26868 21640 26880
rect 21692 26868 21698 26920
rect 21818 26868 21824 26920
rect 21876 26908 21882 26920
rect 22373 26911 22431 26917
rect 22373 26908 22385 26911
rect 21876 26880 22385 26908
rect 21876 26868 21882 26880
rect 22373 26877 22385 26880
rect 22419 26877 22431 26911
rect 22373 26871 22431 26877
rect 21177 26843 21235 26849
rect 21177 26809 21189 26843
rect 21223 26840 21235 26843
rect 21361 26843 21419 26849
rect 21361 26840 21373 26843
rect 21223 26812 21373 26840
rect 21223 26809 21235 26812
rect 21177 26803 21235 26809
rect 21361 26809 21373 26812
rect 21407 26809 21419 26843
rect 22554 26840 22560 26852
rect 21361 26803 21419 26809
rect 21468 26812 22560 26840
rect 16666 26732 16672 26784
rect 16724 26772 16730 26784
rect 21468 26781 21496 26812
rect 22554 26800 22560 26812
rect 22612 26800 22618 26852
rect 16945 26775 17003 26781
rect 16945 26772 16957 26775
rect 16724 26744 16957 26772
rect 16724 26732 16730 26744
rect 16945 26741 16957 26744
rect 16991 26741 17003 26775
rect 16945 26735 17003 26741
rect 21453 26775 21511 26781
rect 21453 26741 21465 26775
rect 21499 26741 21511 26775
rect 21453 26735 21511 26741
rect 1104 26682 26496 26704
rect 1104 26630 4124 26682
rect 4176 26630 4188 26682
rect 4240 26630 4252 26682
rect 4304 26630 4316 26682
rect 4368 26630 4380 26682
rect 4432 26630 10472 26682
rect 10524 26630 10536 26682
rect 10588 26630 10600 26682
rect 10652 26630 10664 26682
rect 10716 26630 10728 26682
rect 10780 26630 16820 26682
rect 16872 26630 16884 26682
rect 16936 26630 16948 26682
rect 17000 26630 17012 26682
rect 17064 26630 17076 26682
rect 17128 26630 23168 26682
rect 23220 26630 23232 26682
rect 23284 26630 23296 26682
rect 23348 26630 23360 26682
rect 23412 26630 23424 26682
rect 23476 26630 26496 26682
rect 1104 26608 26496 26630
rect 16485 26571 16543 26577
rect 16485 26537 16497 26571
rect 16531 26537 16543 26571
rect 16485 26531 16543 26537
rect 15841 26435 15899 26441
rect 15841 26401 15853 26435
rect 15887 26432 15899 26435
rect 16206 26432 16212 26444
rect 15887 26404 16212 26432
rect 15887 26401 15899 26404
rect 15841 26395 15899 26401
rect 16206 26392 16212 26404
rect 16264 26432 16270 26444
rect 16500 26432 16528 26531
rect 16574 26528 16580 26580
rect 16632 26568 16638 26580
rect 16669 26571 16727 26577
rect 16669 26568 16681 26571
rect 16632 26540 16681 26568
rect 16632 26528 16638 26540
rect 16669 26537 16681 26540
rect 16715 26568 16727 26571
rect 17402 26568 17408 26580
rect 16715 26540 17408 26568
rect 16715 26537 16727 26540
rect 16669 26531 16727 26537
rect 17402 26528 17408 26540
rect 17460 26528 17466 26580
rect 17494 26528 17500 26580
rect 17552 26528 17558 26580
rect 20717 26571 20775 26577
rect 20717 26537 20729 26571
rect 20763 26568 20775 26571
rect 20990 26568 20996 26580
rect 20763 26540 20996 26568
rect 20763 26537 20775 26540
rect 20717 26531 20775 26537
rect 20990 26528 20996 26540
rect 21048 26528 21054 26580
rect 21450 26528 21456 26580
rect 21508 26568 21514 26580
rect 22649 26571 22707 26577
rect 22649 26568 22661 26571
rect 21508 26540 22661 26568
rect 21508 26528 21514 26540
rect 22649 26537 22661 26540
rect 22695 26537 22707 26571
rect 22649 26531 22707 26537
rect 16264 26404 16528 26432
rect 16264 26392 16270 26404
rect 16574 26392 16580 26444
rect 16632 26432 16638 26444
rect 17405 26435 17463 26441
rect 17405 26432 17417 26435
rect 16632 26404 17417 26432
rect 16632 26392 16638 26404
rect 17405 26401 17417 26404
rect 17451 26401 17463 26435
rect 17405 26395 17463 26401
rect 22094 26392 22100 26444
rect 22152 26432 22158 26444
rect 22465 26435 22523 26441
rect 22465 26432 22477 26435
rect 22152 26404 22477 26432
rect 22152 26392 22158 26404
rect 22465 26401 22477 26404
rect 22511 26401 22523 26435
rect 22465 26395 22523 26401
rect 9490 26324 9496 26376
rect 9548 26324 9554 26376
rect 11422 26324 11428 26376
rect 11480 26324 11486 26376
rect 12526 26324 12532 26376
rect 12584 26324 12590 26376
rect 12713 26367 12771 26373
rect 12713 26333 12725 26367
rect 12759 26364 12771 26367
rect 12894 26364 12900 26376
rect 12759 26336 12900 26364
rect 12759 26333 12771 26336
rect 12713 26327 12771 26333
rect 12894 26324 12900 26336
rect 12952 26324 12958 26376
rect 15922 26367 15980 26373
rect 15922 26364 15934 26367
rect 15856 26336 15934 26364
rect 15856 26296 15884 26336
rect 15922 26333 15934 26336
rect 15968 26333 15980 26367
rect 15922 26327 15980 26333
rect 16022 26324 16028 26376
rect 16080 26324 16086 26376
rect 16114 26324 16120 26376
rect 16172 26324 16178 26376
rect 16758 26364 16764 26376
rect 16316 26336 16764 26364
rect 16316 26305 16344 26336
rect 16758 26324 16764 26336
rect 16816 26324 16822 26376
rect 18046 26324 18052 26376
rect 18104 26324 18110 26376
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26364 19487 26367
rect 19610 26364 19616 26376
rect 19475 26336 19616 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 19610 26324 19616 26336
rect 19668 26324 19674 26376
rect 19702 26324 19708 26376
rect 19760 26324 19766 26376
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 19981 26367 20039 26373
rect 19981 26364 19993 26367
rect 19935 26336 19993 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 19981 26333 19993 26336
rect 20027 26333 20039 26367
rect 19981 26327 20039 26333
rect 20533 26367 20591 26373
rect 20533 26333 20545 26367
rect 20579 26364 20591 26367
rect 21266 26364 21272 26376
rect 20579 26336 21272 26364
rect 20579 26333 20591 26336
rect 20533 26327 20591 26333
rect 16301 26299 16359 26305
rect 16301 26296 16313 26299
rect 15856 26268 16313 26296
rect 16301 26265 16313 26268
rect 16347 26265 16359 26299
rect 16301 26259 16359 26265
rect 16482 26256 16488 26308
rect 16540 26305 16546 26308
rect 16540 26299 16559 26305
rect 16547 26265 16559 26299
rect 20548 26296 20576 26327
rect 21266 26324 21272 26336
rect 21324 26324 21330 26376
rect 22370 26324 22376 26376
rect 22428 26324 22434 26376
rect 22741 26367 22799 26373
rect 22741 26333 22753 26367
rect 22787 26333 22799 26367
rect 22741 26327 22799 26333
rect 22756 26296 22784 26327
rect 16540 26259 16559 26265
rect 19904 26268 20576 26296
rect 22066 26268 22784 26296
rect 16540 26256 16546 26259
rect 19904 26240 19932 26268
rect 9306 26188 9312 26240
rect 9364 26188 9370 26240
rect 10318 26188 10324 26240
rect 10376 26228 10382 26240
rect 10781 26231 10839 26237
rect 10781 26228 10793 26231
rect 10376 26200 10793 26228
rect 10376 26188 10382 26200
rect 10781 26197 10793 26200
rect 10827 26197 10839 26231
rect 10781 26191 10839 26197
rect 12618 26188 12624 26240
rect 12676 26188 12682 26240
rect 15654 26188 15660 26240
rect 15712 26188 15718 26240
rect 19242 26188 19248 26240
rect 19300 26188 19306 26240
rect 19886 26188 19892 26240
rect 19944 26188 19950 26240
rect 21726 26188 21732 26240
rect 21784 26228 21790 26240
rect 22066 26228 22094 26268
rect 21784 26200 22094 26228
rect 21784 26188 21790 26200
rect 22462 26188 22468 26240
rect 22520 26188 22526 26240
rect 1104 26138 26656 26160
rect 1104 26086 7298 26138
rect 7350 26086 7362 26138
rect 7414 26086 7426 26138
rect 7478 26086 7490 26138
rect 7542 26086 7554 26138
rect 7606 26086 13646 26138
rect 13698 26086 13710 26138
rect 13762 26086 13774 26138
rect 13826 26086 13838 26138
rect 13890 26086 13902 26138
rect 13954 26086 19994 26138
rect 20046 26086 20058 26138
rect 20110 26086 20122 26138
rect 20174 26086 20186 26138
rect 20238 26086 20250 26138
rect 20302 26086 26342 26138
rect 26394 26086 26406 26138
rect 26458 26086 26470 26138
rect 26522 26086 26534 26138
rect 26586 26086 26598 26138
rect 26650 26086 26656 26138
rect 1104 26064 26656 26086
rect 15930 26024 15936 26036
rect 13832 25996 15936 26024
rect 12437 25959 12495 25965
rect 8220 25928 10732 25956
rect 8110 25848 8116 25900
rect 8168 25888 8174 25900
rect 8220 25897 8248 25928
rect 8205 25891 8263 25897
rect 8205 25888 8217 25891
rect 8168 25860 8217 25888
rect 8168 25848 8174 25860
rect 8205 25857 8217 25860
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 8472 25891 8530 25897
rect 8472 25857 8484 25891
rect 8518 25888 8530 25891
rect 9306 25888 9312 25900
rect 8518 25860 9312 25888
rect 8518 25857 8530 25860
rect 8472 25851 8530 25857
rect 9306 25848 9312 25860
rect 9364 25848 9370 25900
rect 9692 25897 9720 25928
rect 9950 25897 9956 25900
rect 9677 25891 9735 25897
rect 9677 25857 9689 25891
rect 9723 25857 9735 25891
rect 9677 25851 9735 25857
rect 9944 25851 9956 25897
rect 9950 25848 9956 25851
rect 10008 25848 10014 25900
rect 10704 25820 10732 25928
rect 10980 25928 11652 25956
rect 10980 25900 11008 25928
rect 10962 25848 10968 25900
rect 11020 25848 11026 25900
rect 11330 25848 11336 25900
rect 11388 25848 11394 25900
rect 11624 25897 11652 25928
rect 12437 25925 12449 25959
rect 12483 25956 12495 25959
rect 12897 25959 12955 25965
rect 12897 25956 12909 25959
rect 12483 25928 12909 25956
rect 12483 25925 12495 25928
rect 12437 25919 12495 25925
rect 12897 25925 12909 25928
rect 12943 25925 12955 25959
rect 12897 25919 12955 25925
rect 13096 25928 13492 25956
rect 11609 25891 11667 25897
rect 11609 25857 11621 25891
rect 11655 25857 11667 25891
rect 11609 25851 11667 25857
rect 12342 25848 12348 25900
rect 12400 25848 12406 25900
rect 13096 25897 13124 25928
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25857 12587 25891
rect 12667 25891 12725 25897
rect 12667 25888 12679 25891
rect 12529 25851 12587 25857
rect 12662 25857 12679 25888
rect 12713 25857 12725 25891
rect 12662 25851 12725 25857
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25857 13139 25891
rect 13081 25851 13139 25857
rect 13265 25891 13323 25897
rect 13265 25857 13277 25891
rect 13311 25857 13323 25891
rect 13265 25851 13323 25857
rect 11238 25820 11244 25832
rect 10704 25792 11244 25820
rect 11238 25780 11244 25792
rect 11296 25780 11302 25832
rect 12250 25780 12256 25832
rect 12308 25820 12314 25832
rect 12545 25820 12573 25851
rect 12308 25792 12573 25820
rect 12308 25780 12314 25792
rect 11057 25755 11115 25761
rect 11057 25721 11069 25755
rect 11103 25752 11115 25755
rect 11422 25752 11428 25764
rect 11103 25724 11428 25752
rect 11103 25721 11115 25724
rect 11057 25715 11115 25721
rect 11422 25712 11428 25724
rect 11480 25752 11486 25764
rect 12069 25755 12127 25761
rect 11480 25724 11836 25752
rect 11480 25712 11486 25724
rect 11808 25696 11836 25724
rect 12069 25721 12081 25755
rect 12115 25752 12127 25755
rect 12434 25752 12440 25764
rect 12115 25724 12440 25752
rect 12115 25721 12127 25724
rect 12069 25715 12127 25721
rect 12434 25712 12440 25724
rect 12492 25752 12498 25764
rect 12662 25752 12690 25851
rect 12805 25823 12863 25829
rect 12805 25789 12817 25823
rect 12851 25820 12863 25823
rect 13096 25820 13124 25851
rect 12851 25792 13124 25820
rect 12851 25789 12863 25792
rect 12805 25783 12863 25789
rect 12492 25724 12690 25752
rect 12492 25712 12498 25724
rect 9585 25687 9643 25693
rect 9585 25653 9597 25687
rect 9631 25684 9643 25687
rect 9858 25684 9864 25696
rect 9631 25656 9864 25684
rect 9631 25653 9643 25656
rect 9585 25647 9643 25653
rect 9858 25644 9864 25656
rect 9916 25644 9922 25696
rect 11146 25644 11152 25696
rect 11204 25644 11210 25696
rect 11790 25644 11796 25696
rect 11848 25644 11854 25696
rect 11974 25644 11980 25696
rect 12032 25684 12038 25696
rect 12161 25687 12219 25693
rect 12161 25684 12173 25687
rect 12032 25656 12173 25684
rect 12032 25644 12038 25656
rect 12161 25653 12173 25656
rect 12207 25653 12219 25687
rect 12161 25647 12219 25653
rect 12250 25644 12256 25696
rect 12308 25684 12314 25696
rect 12820 25684 12848 25783
rect 13280 25752 13308 25851
rect 13354 25848 13360 25900
rect 13412 25848 13418 25900
rect 13464 25897 13492 25928
rect 13538 25916 13544 25968
rect 13596 25916 13602 25968
rect 13832 25897 13860 25996
rect 15930 25984 15936 25996
rect 15988 25984 15994 26036
rect 16669 26027 16727 26033
rect 16669 25993 16681 26027
rect 16715 26024 16727 26027
rect 16758 26024 16764 26036
rect 16715 25996 16764 26024
rect 16715 25993 16727 25996
rect 16669 25987 16727 25993
rect 14550 25916 14556 25968
rect 14608 25956 14614 25968
rect 15565 25959 15623 25965
rect 15565 25956 15577 25959
rect 14608 25928 15577 25956
rect 14608 25916 14614 25928
rect 15565 25925 15577 25928
rect 15611 25956 15623 25959
rect 15746 25956 15752 25968
rect 15611 25928 15752 25956
rect 15611 25925 15623 25928
rect 15565 25919 15623 25925
rect 15746 25916 15752 25928
rect 15804 25956 15810 25968
rect 16114 25956 16120 25968
rect 15804 25928 16120 25956
rect 15804 25916 15810 25928
rect 16114 25916 16120 25928
rect 16172 25916 16178 25968
rect 13449 25891 13507 25897
rect 13449 25857 13461 25891
rect 13495 25857 13507 25891
rect 13449 25851 13507 25857
rect 13725 25891 13783 25897
rect 13725 25857 13737 25891
rect 13771 25888 13783 25891
rect 13817 25891 13875 25897
rect 13817 25888 13829 25891
rect 13771 25860 13829 25888
rect 13771 25857 13783 25860
rect 13725 25851 13783 25857
rect 13817 25857 13829 25860
rect 13863 25857 13875 25891
rect 13817 25851 13875 25857
rect 14645 25891 14703 25897
rect 14645 25857 14657 25891
rect 14691 25888 14703 25891
rect 15010 25888 15016 25900
rect 14691 25860 15016 25888
rect 14691 25857 14703 25860
rect 14645 25851 14703 25857
rect 13369 25820 13397 25848
rect 13740 25820 13768 25851
rect 15010 25848 15016 25860
rect 15068 25848 15074 25900
rect 15105 25891 15163 25897
rect 15105 25857 15117 25891
rect 15151 25888 15163 25891
rect 16022 25888 16028 25900
rect 15151 25860 16028 25888
rect 15151 25857 15163 25860
rect 15105 25851 15163 25857
rect 16022 25848 16028 25860
rect 16080 25848 16086 25900
rect 16206 25848 16212 25900
rect 16264 25848 16270 25900
rect 13369 25792 13768 25820
rect 14369 25823 14427 25829
rect 14369 25789 14381 25823
rect 14415 25789 14427 25823
rect 14369 25783 14427 25789
rect 13538 25752 13544 25764
rect 13280 25724 13544 25752
rect 13538 25712 13544 25724
rect 13596 25712 13602 25764
rect 14384 25752 14412 25783
rect 14458 25780 14464 25832
rect 14516 25780 14522 25832
rect 15289 25823 15347 25829
rect 15289 25789 15301 25823
rect 15335 25820 15347 25823
rect 16224 25820 16252 25848
rect 15335 25792 16252 25820
rect 15335 25789 15347 25792
rect 15289 25783 15347 25789
rect 15657 25755 15715 25761
rect 15657 25752 15669 25755
rect 14384 25724 15669 25752
rect 15657 25721 15669 25724
rect 15703 25721 15715 25755
rect 15657 25715 15715 25721
rect 12308 25656 12848 25684
rect 12308 25644 12314 25656
rect 13630 25644 13636 25696
rect 13688 25644 13694 25696
rect 13909 25687 13967 25693
rect 13909 25653 13921 25687
rect 13955 25684 13967 25687
rect 14274 25684 14280 25696
rect 13955 25656 14280 25684
rect 13955 25653 13967 25656
rect 13909 25647 13967 25653
rect 14274 25644 14280 25656
rect 14332 25644 14338 25696
rect 14826 25644 14832 25696
rect 14884 25644 14890 25696
rect 14918 25644 14924 25696
rect 14976 25644 14982 25696
rect 15473 25687 15531 25693
rect 15473 25653 15485 25687
rect 15519 25684 15531 25687
rect 16390 25684 16396 25696
rect 15519 25656 16396 25684
rect 15519 25653 15531 25656
rect 15473 25647 15531 25653
rect 16390 25644 16396 25656
rect 16448 25684 16454 25696
rect 16684 25684 16712 25987
rect 16758 25984 16764 25996
rect 16816 25984 16822 26036
rect 20625 26027 20683 26033
rect 20625 25993 20637 26027
rect 20671 26024 20683 26027
rect 21726 26024 21732 26036
rect 20671 25996 21732 26024
rect 20671 25993 20683 25996
rect 20625 25987 20683 25993
rect 21726 25984 21732 25996
rect 21784 25984 21790 26036
rect 21818 25984 21824 26036
rect 21876 25984 21882 26036
rect 18868 25959 18926 25965
rect 18868 25925 18880 25959
rect 18914 25956 18926 25959
rect 19242 25956 19248 25968
rect 18914 25928 19248 25956
rect 18914 25925 18926 25928
rect 18868 25919 18926 25925
rect 19242 25916 19248 25928
rect 19300 25916 19306 25968
rect 20241 25959 20299 25965
rect 20241 25925 20253 25959
rect 20287 25956 20299 25959
rect 20441 25959 20499 25965
rect 20441 25956 20453 25959
rect 20287 25925 20300 25956
rect 20241 25919 20300 25925
rect 17494 25848 17500 25900
rect 17552 25888 17558 25900
rect 17782 25891 17840 25897
rect 17782 25888 17794 25891
rect 17552 25860 17794 25888
rect 17552 25848 17558 25860
rect 17782 25857 17794 25860
rect 17828 25857 17840 25891
rect 19150 25888 19156 25900
rect 17782 25851 17840 25857
rect 18616 25860 19156 25888
rect 18616 25829 18644 25860
rect 19150 25848 19156 25860
rect 19208 25848 19214 25900
rect 18049 25823 18107 25829
rect 18049 25789 18061 25823
rect 18095 25820 18107 25823
rect 18601 25823 18659 25829
rect 18601 25820 18613 25823
rect 18095 25792 18613 25820
rect 18095 25789 18107 25792
rect 18049 25783 18107 25789
rect 18601 25789 18613 25792
rect 18647 25789 18659 25823
rect 20272 25820 20300 25919
rect 20364 25928 20453 25956
rect 20364 25900 20392 25928
rect 20441 25925 20453 25928
rect 20487 25925 20499 25959
rect 20441 25919 20499 25925
rect 20809 25959 20867 25965
rect 20809 25925 20821 25959
rect 20855 25956 20867 25959
rect 22462 25956 22468 25968
rect 20855 25928 22468 25956
rect 20855 25925 20867 25928
rect 20809 25919 20867 25925
rect 22462 25916 22468 25928
rect 22520 25916 22526 25968
rect 22554 25916 22560 25968
rect 22612 25916 22618 25968
rect 22738 25916 22744 25968
rect 22796 25956 22802 25968
rect 22796 25928 23244 25956
rect 22796 25916 22802 25928
rect 20346 25848 20352 25900
rect 20404 25848 20410 25900
rect 20533 25891 20591 25897
rect 20533 25857 20545 25891
rect 20579 25888 20591 25891
rect 20579 25860 20944 25888
rect 20579 25857 20591 25860
rect 20533 25851 20591 25857
rect 20806 25820 20812 25832
rect 20272 25792 20812 25820
rect 18601 25783 18659 25789
rect 20806 25780 20812 25792
rect 20864 25780 20870 25832
rect 20916 25829 20944 25860
rect 21082 25848 21088 25900
rect 21140 25848 21146 25900
rect 21174 25848 21180 25900
rect 21232 25848 21238 25900
rect 21266 25848 21272 25900
rect 21324 25848 21330 25900
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25888 21511 25891
rect 21818 25888 21824 25900
rect 21499 25860 21824 25888
rect 21499 25857 21511 25860
rect 21453 25851 21511 25857
rect 21818 25848 21824 25860
rect 21876 25848 21882 25900
rect 22572 25888 22600 25916
rect 23216 25897 23244 25928
rect 22934 25891 22992 25897
rect 22934 25888 22946 25891
rect 22572 25860 22946 25888
rect 22934 25857 22946 25860
rect 22980 25857 22992 25891
rect 22934 25851 22992 25857
rect 23201 25891 23259 25897
rect 23201 25857 23213 25891
rect 23247 25857 23259 25891
rect 23201 25851 23259 25857
rect 20901 25823 20959 25829
rect 20901 25789 20913 25823
rect 20947 25820 20959 25823
rect 20947 25792 21496 25820
rect 20947 25789 20959 25792
rect 20901 25783 20959 25789
rect 21468 25764 21496 25792
rect 20073 25755 20131 25761
rect 20073 25752 20085 25755
rect 19720 25724 20085 25752
rect 19720 25696 19748 25724
rect 20073 25721 20085 25724
rect 20119 25721 20131 25755
rect 20073 25715 20131 25721
rect 20272 25724 21128 25752
rect 16448 25656 16712 25684
rect 16448 25644 16454 25656
rect 19702 25644 19708 25696
rect 19760 25644 19766 25696
rect 19886 25644 19892 25696
rect 19944 25684 19950 25696
rect 20272 25693 20300 25724
rect 21100 25696 21128 25724
rect 21450 25712 21456 25764
rect 21508 25712 21514 25764
rect 19981 25687 20039 25693
rect 19981 25684 19993 25687
rect 19944 25656 19993 25684
rect 19944 25644 19950 25656
rect 19981 25653 19993 25656
rect 20027 25653 20039 25687
rect 19981 25647 20039 25653
rect 20257 25687 20315 25693
rect 20257 25653 20269 25687
rect 20303 25653 20315 25687
rect 20257 25647 20315 25653
rect 20806 25644 20812 25696
rect 20864 25644 20870 25696
rect 21082 25644 21088 25696
rect 21140 25644 21146 25696
rect 1104 25594 26496 25616
rect 1104 25542 4124 25594
rect 4176 25542 4188 25594
rect 4240 25542 4252 25594
rect 4304 25542 4316 25594
rect 4368 25542 4380 25594
rect 4432 25542 10472 25594
rect 10524 25542 10536 25594
rect 10588 25542 10600 25594
rect 10652 25542 10664 25594
rect 10716 25542 10728 25594
rect 10780 25542 16820 25594
rect 16872 25542 16884 25594
rect 16936 25542 16948 25594
rect 17000 25542 17012 25594
rect 17064 25542 17076 25594
rect 17128 25542 23168 25594
rect 23220 25542 23232 25594
rect 23284 25542 23296 25594
rect 23348 25542 23360 25594
rect 23412 25542 23424 25594
rect 23476 25542 26496 25594
rect 1104 25520 26496 25542
rect 9490 25440 9496 25492
rect 9548 25440 9554 25492
rect 9677 25483 9735 25489
rect 9677 25449 9689 25483
rect 9723 25480 9735 25483
rect 9766 25480 9772 25492
rect 9723 25452 9772 25480
rect 9723 25449 9735 25452
rect 9677 25443 9735 25449
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 9950 25440 9956 25492
rect 10008 25440 10014 25492
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 13725 25483 13783 25489
rect 12492 25452 13676 25480
rect 12492 25440 12498 25452
rect 13648 25412 13676 25452
rect 13725 25449 13737 25483
rect 13771 25480 13783 25483
rect 14093 25483 14151 25489
rect 14093 25480 14105 25483
rect 13771 25452 14105 25480
rect 13771 25449 13783 25452
rect 13725 25443 13783 25449
rect 14093 25449 14105 25452
rect 14139 25449 14151 25483
rect 14093 25443 14151 25449
rect 14274 25440 14280 25492
rect 14332 25480 14338 25492
rect 14332 25452 14688 25480
rect 14332 25440 14338 25452
rect 13648 25384 14320 25412
rect 14182 25344 14188 25356
rect 13556 25316 14188 25344
rect 10140 25257 10198 25263
rect 10140 25223 10152 25257
rect 10186 25223 10198 25257
rect 10226 25236 10232 25288
rect 10284 25236 10290 25288
rect 10410 25236 10416 25288
rect 10468 25236 10474 25288
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25245 10563 25279
rect 10505 25239 10563 25245
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25276 10655 25279
rect 11238 25276 11244 25288
rect 10643 25248 11244 25276
rect 10643 25245 10655 25248
rect 10597 25239 10655 25245
rect 10140 25220 10198 25223
rect 9858 25168 9864 25220
rect 9916 25168 9922 25220
rect 10134 25168 10140 25220
rect 10192 25168 10198 25220
rect 10318 25168 10324 25220
rect 10376 25208 10382 25220
rect 10520 25208 10548 25239
rect 11238 25236 11244 25248
rect 11296 25276 11302 25288
rect 12069 25279 12127 25285
rect 12069 25276 12081 25279
rect 11296 25248 12081 25276
rect 11296 25236 11302 25248
rect 12069 25245 12081 25248
rect 12115 25245 12127 25279
rect 12069 25239 12127 25245
rect 12336 25279 12394 25285
rect 12336 25245 12348 25279
rect 12382 25276 12394 25279
rect 12618 25276 12624 25288
rect 12382 25248 12624 25276
rect 12382 25245 12394 25248
rect 12336 25239 12394 25245
rect 12618 25236 12624 25248
rect 12676 25236 12682 25288
rect 10376 25180 10548 25208
rect 10864 25211 10922 25217
rect 10376 25168 10382 25180
rect 10864 25177 10876 25211
rect 10910 25208 10922 25211
rect 11146 25208 11152 25220
rect 10910 25180 11152 25208
rect 10910 25177 10922 25180
rect 10864 25171 10922 25177
rect 11146 25168 11152 25180
rect 11204 25168 11210 25220
rect 13556 25217 13584 25316
rect 14182 25304 14188 25316
rect 14240 25304 14246 25356
rect 14292 25288 14320 25384
rect 14550 25372 14556 25424
rect 14608 25372 14614 25424
rect 14568 25344 14596 25372
rect 14384 25316 14596 25344
rect 14274 25236 14280 25288
rect 14332 25236 14338 25288
rect 14384 25285 14412 25316
rect 14369 25279 14427 25285
rect 14369 25245 14381 25279
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 14458 25236 14464 25288
rect 14516 25236 14522 25288
rect 14660 25285 14688 25452
rect 15010 25440 15016 25492
rect 15068 25480 15074 25492
rect 16209 25483 16267 25489
rect 16209 25480 16221 25483
rect 15068 25452 16221 25480
rect 15068 25440 15074 25452
rect 16209 25449 16221 25452
rect 16255 25449 16267 25483
rect 17865 25483 17923 25489
rect 17865 25480 17877 25483
rect 16209 25443 16267 25449
rect 16316 25452 17877 25480
rect 16022 25372 16028 25424
rect 16080 25412 16086 25424
rect 16316 25412 16344 25452
rect 17865 25449 17877 25452
rect 17911 25480 17923 25483
rect 18046 25480 18052 25492
rect 17911 25452 18052 25480
rect 17911 25449 17923 25452
rect 17865 25443 17923 25449
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 18969 25483 19027 25489
rect 18969 25449 18981 25483
rect 19015 25480 19027 25483
rect 20714 25480 20720 25492
rect 19015 25452 20720 25480
rect 19015 25449 19027 25452
rect 18969 25443 19027 25449
rect 20714 25440 20720 25452
rect 20772 25440 20778 25492
rect 20806 25440 20812 25492
rect 20864 25440 20870 25492
rect 22370 25440 22376 25492
rect 22428 25480 22434 25492
rect 22741 25483 22799 25489
rect 22741 25480 22753 25483
rect 22428 25452 22753 25480
rect 22428 25440 22434 25452
rect 22741 25449 22753 25452
rect 22787 25449 22799 25483
rect 22741 25443 22799 25449
rect 16080 25384 16344 25412
rect 18340 25384 19012 25412
rect 16080 25372 16086 25384
rect 16485 25347 16543 25353
rect 16485 25344 16497 25347
rect 15764 25316 16497 25344
rect 14645 25279 14703 25285
rect 14645 25245 14657 25279
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 14734 25236 14740 25288
rect 14792 25276 14798 25288
rect 15764 25276 15792 25316
rect 16485 25313 16497 25316
rect 16531 25313 16543 25347
rect 16485 25307 16543 25313
rect 14792 25248 15792 25276
rect 14792 25236 14798 25248
rect 16114 25236 16120 25288
rect 16172 25276 16178 25288
rect 16209 25279 16267 25285
rect 16209 25276 16221 25279
rect 16172 25248 16221 25276
rect 16172 25236 16178 25248
rect 16209 25245 16221 25248
rect 16255 25245 16267 25279
rect 16209 25239 16267 25245
rect 16298 25236 16304 25288
rect 16356 25276 16362 25288
rect 16393 25279 16451 25285
rect 16393 25276 16405 25279
rect 16356 25248 16405 25276
rect 16356 25236 16362 25248
rect 16393 25245 16405 25248
rect 16439 25245 16451 25279
rect 16393 25239 16451 25245
rect 16752 25279 16810 25285
rect 16752 25245 16764 25279
rect 16798 25245 16810 25279
rect 16752 25239 16810 25245
rect 13541 25211 13599 25217
rect 13541 25208 13553 25211
rect 11900 25180 13553 25208
rect 9661 25143 9719 25149
rect 9661 25109 9673 25143
rect 9707 25140 9719 25143
rect 10594 25140 10600 25152
rect 9707 25112 10600 25140
rect 9707 25109 9719 25112
rect 9661 25103 9719 25109
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 10778 25100 10784 25152
rect 10836 25140 10842 25152
rect 11900 25140 11928 25180
rect 13541 25177 13553 25180
rect 13587 25177 13599 25211
rect 13541 25171 13599 25177
rect 13757 25211 13815 25217
rect 13757 25177 13769 25211
rect 13803 25208 13815 25211
rect 13803 25180 14320 25208
rect 13803 25177 13815 25180
rect 13757 25171 13815 25177
rect 10836 25112 11928 25140
rect 11977 25143 12035 25149
rect 10836 25100 10842 25112
rect 11977 25109 11989 25143
rect 12023 25140 12035 25143
rect 12250 25140 12256 25152
rect 12023 25112 12256 25140
rect 12023 25109 12035 25112
rect 11977 25103 12035 25109
rect 12250 25100 12256 25112
rect 12308 25100 12314 25152
rect 13446 25100 13452 25152
rect 13504 25100 13510 25152
rect 13909 25143 13967 25149
rect 13909 25109 13921 25143
rect 13955 25140 13967 25143
rect 13998 25140 14004 25152
rect 13955 25112 14004 25140
rect 13955 25109 13967 25112
rect 13909 25103 13967 25109
rect 13998 25100 14004 25112
rect 14056 25100 14062 25152
rect 14292 25140 14320 25180
rect 14826 25168 14832 25220
rect 14884 25208 14890 25220
rect 14982 25211 15040 25217
rect 14982 25208 14994 25211
rect 14884 25180 14994 25208
rect 14884 25168 14890 25180
rect 14982 25177 14994 25180
rect 15028 25177 15040 25211
rect 14982 25171 15040 25177
rect 15654 25168 15660 25220
rect 15712 25168 15718 25220
rect 15672 25140 15700 25168
rect 14292 25112 15700 25140
rect 16117 25143 16175 25149
rect 16117 25109 16129 25143
rect 16163 25140 16175 25143
rect 16206 25140 16212 25152
rect 16163 25112 16212 25140
rect 16163 25109 16175 25112
rect 16117 25103 16175 25109
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 16408 25140 16436 25239
rect 16666 25168 16672 25220
rect 16724 25208 16730 25220
rect 16776 25208 16804 25239
rect 17310 25236 17316 25288
rect 17368 25276 17374 25288
rect 18340 25285 18368 25384
rect 18417 25347 18475 25353
rect 18417 25313 18429 25347
rect 18463 25344 18475 25347
rect 18463 25316 18828 25344
rect 18463 25313 18475 25316
rect 18417 25307 18475 25313
rect 18800 25285 18828 25316
rect 17957 25279 18015 25285
rect 17957 25276 17969 25279
rect 17368 25248 17969 25276
rect 17368 25236 17374 25248
rect 17957 25245 17969 25248
rect 18003 25245 18015 25279
rect 17957 25239 18015 25245
rect 18141 25279 18199 25285
rect 18141 25245 18153 25279
rect 18187 25276 18199 25279
rect 18325 25279 18383 25285
rect 18325 25276 18337 25279
rect 18187 25248 18337 25276
rect 18187 25245 18199 25248
rect 18141 25239 18199 25245
rect 18325 25245 18337 25248
rect 18371 25245 18383 25279
rect 18325 25239 18383 25245
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25245 18567 25279
rect 18800 25279 18873 25285
rect 18800 25248 18827 25279
rect 18509 25239 18567 25245
rect 18815 25245 18827 25248
rect 18861 25245 18873 25279
rect 18815 25239 18873 25245
rect 18156 25208 18184 25239
rect 16724 25180 16804 25208
rect 17972 25180 18184 25208
rect 18524 25208 18552 25239
rect 18984 25208 19012 25384
rect 19061 25347 19119 25353
rect 19061 25313 19073 25347
rect 19107 25344 19119 25347
rect 19107 25316 19380 25344
rect 19107 25313 19119 25316
rect 19061 25307 19119 25313
rect 19352 25288 19380 25316
rect 19150 25236 19156 25288
rect 19208 25276 19214 25288
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 19208 25248 19257 25276
rect 19208 25236 19214 25248
rect 19245 25245 19257 25248
rect 19291 25245 19303 25279
rect 19245 25239 19303 25245
rect 19334 25236 19340 25288
rect 19392 25236 19398 25288
rect 20622 25276 20628 25288
rect 19444 25248 20628 25276
rect 19444 25208 19472 25248
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 19518 25217 19524 25220
rect 18524 25180 18736 25208
rect 18984 25180 19472 25208
rect 16724 25168 16730 25180
rect 17972 25140 18000 25180
rect 16408 25112 18000 25140
rect 18046 25100 18052 25152
rect 18104 25100 18110 25152
rect 18598 25100 18604 25152
rect 18656 25100 18662 25152
rect 18708 25140 18736 25180
rect 19512 25171 19524 25217
rect 19518 25168 19524 25171
rect 19576 25168 19582 25220
rect 19794 25168 19800 25220
rect 19852 25208 19858 25220
rect 20824 25208 20852 25440
rect 20898 25236 20904 25288
rect 20956 25236 20962 25288
rect 21082 25236 21088 25288
rect 21140 25236 21146 25288
rect 21361 25279 21419 25285
rect 21361 25245 21373 25279
rect 21407 25276 21419 25279
rect 22738 25276 22744 25288
rect 21407 25248 22744 25276
rect 21407 25245 21419 25248
rect 21361 25239 21419 25245
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 21606 25211 21664 25217
rect 21606 25208 21618 25211
rect 19852 25180 20760 25208
rect 20824 25180 21618 25208
rect 19852 25168 19858 25180
rect 19812 25140 19840 25168
rect 18708 25112 19840 25140
rect 20346 25100 20352 25152
rect 20404 25140 20410 25152
rect 20732 25149 20760 25180
rect 21606 25177 21618 25180
rect 21652 25177 21664 25211
rect 21606 25171 21664 25177
rect 20625 25143 20683 25149
rect 20625 25140 20637 25143
rect 20404 25112 20637 25140
rect 20404 25100 20410 25112
rect 20625 25109 20637 25112
rect 20671 25109 20683 25143
rect 20625 25103 20683 25109
rect 20717 25143 20775 25149
rect 20717 25109 20729 25143
rect 20763 25140 20775 25143
rect 20990 25140 20996 25152
rect 20763 25112 20996 25140
rect 20763 25109 20775 25112
rect 20717 25103 20775 25109
rect 20990 25100 20996 25112
rect 21048 25100 21054 25152
rect 1104 25050 26656 25072
rect 1104 24998 7298 25050
rect 7350 24998 7362 25050
rect 7414 24998 7426 25050
rect 7478 24998 7490 25050
rect 7542 24998 7554 25050
rect 7606 24998 13646 25050
rect 13698 24998 13710 25050
rect 13762 24998 13774 25050
rect 13826 24998 13838 25050
rect 13890 24998 13902 25050
rect 13954 24998 19994 25050
rect 20046 24998 20058 25050
rect 20110 24998 20122 25050
rect 20174 24998 20186 25050
rect 20238 24998 20250 25050
rect 20302 24998 26342 25050
rect 26394 24998 26406 25050
rect 26458 24998 26470 25050
rect 26522 24998 26534 25050
rect 26586 24998 26598 25050
rect 26650 24998 26656 25050
rect 1104 24976 26656 24998
rect 10594 24896 10600 24948
rect 10652 24896 10658 24948
rect 11330 24896 11336 24948
rect 11388 24896 11394 24948
rect 12618 24896 12624 24948
rect 12676 24936 12682 24948
rect 13354 24936 13360 24948
rect 12676 24908 13360 24936
rect 12676 24896 12682 24908
rect 13354 24896 13360 24908
rect 13412 24896 13418 24948
rect 13909 24939 13967 24945
rect 13909 24905 13921 24939
rect 13955 24936 13967 24939
rect 14458 24936 14464 24948
rect 13955 24908 14464 24936
rect 13955 24905 13967 24908
rect 13909 24899 13967 24905
rect 14458 24896 14464 24908
rect 14516 24896 14522 24948
rect 14918 24896 14924 24948
rect 14976 24896 14982 24948
rect 15746 24896 15752 24948
rect 15804 24896 15810 24948
rect 15930 24896 15936 24948
rect 15988 24896 15994 24948
rect 16022 24896 16028 24948
rect 16080 24896 16086 24948
rect 16117 24939 16175 24945
rect 16117 24905 16129 24939
rect 16163 24936 16175 24939
rect 16206 24936 16212 24948
rect 16163 24908 16212 24936
rect 16163 24905 16175 24908
rect 16117 24899 16175 24905
rect 16206 24896 16212 24908
rect 16264 24896 16270 24948
rect 16390 24896 16396 24948
rect 16448 24896 16454 24948
rect 17129 24939 17187 24945
rect 17129 24905 17141 24939
rect 17175 24936 17187 24939
rect 17494 24936 17500 24948
rect 17175 24908 17500 24936
rect 17175 24905 17187 24908
rect 17129 24899 17187 24905
rect 17494 24896 17500 24908
rect 17552 24896 17558 24948
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19797 24939 19855 24945
rect 19797 24936 19809 24939
rect 19392 24908 19809 24936
rect 19392 24896 19398 24908
rect 19797 24905 19809 24908
rect 19843 24905 19855 24939
rect 19797 24899 19855 24905
rect 21082 24896 21088 24948
rect 21140 24936 21146 24948
rect 21979 24939 22037 24945
rect 21979 24936 21991 24939
rect 21140 24908 21991 24936
rect 21140 24896 21146 24908
rect 9769 24871 9827 24877
rect 9769 24837 9781 24871
rect 9815 24868 9827 24871
rect 9858 24868 9864 24880
rect 9815 24840 9864 24868
rect 9815 24837 9827 24840
rect 9769 24831 9827 24837
rect 9858 24828 9864 24840
rect 9916 24828 9922 24880
rect 10226 24828 10232 24880
rect 10284 24868 10290 24880
rect 11885 24871 11943 24877
rect 11885 24868 11897 24871
rect 10284 24840 11897 24868
rect 10284 24828 10290 24840
rect 9122 24760 9128 24812
rect 9180 24760 9186 24812
rect 9582 24760 9588 24812
rect 9640 24760 9646 24812
rect 9217 24735 9275 24741
rect 9217 24701 9229 24735
rect 9263 24732 9275 24735
rect 9674 24732 9680 24744
rect 9263 24704 9680 24732
rect 9263 24701 9275 24704
rect 9217 24695 9275 24701
rect 9674 24692 9680 24704
rect 9732 24692 9738 24744
rect 9876 24732 9904 24828
rect 10796 24809 10824 24840
rect 11885 24837 11897 24840
rect 11931 24868 11943 24871
rect 11931 24840 12434 24868
rect 11931 24837 11943 24840
rect 11885 24831 11943 24837
rect 10321 24803 10379 24809
rect 10321 24769 10333 24803
rect 10367 24800 10379 24803
rect 10597 24803 10655 24809
rect 10597 24800 10609 24803
rect 10367 24772 10609 24800
rect 10367 24769 10379 24772
rect 10321 24763 10379 24769
rect 10597 24769 10609 24772
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 11149 24803 11207 24809
rect 11149 24769 11161 24803
rect 11195 24800 11207 24803
rect 11974 24800 11980 24812
rect 11195 24772 11980 24800
rect 11195 24769 11207 24772
rect 11149 24763 11207 24769
rect 10226 24732 10232 24744
rect 9876 24704 10232 24732
rect 10226 24692 10232 24704
rect 10284 24732 10290 24744
rect 10505 24735 10563 24741
rect 10505 24732 10517 24735
rect 10284 24704 10517 24732
rect 10284 24692 10290 24704
rect 10505 24701 10517 24704
rect 10551 24701 10563 24735
rect 10505 24695 10563 24701
rect 9493 24667 9551 24673
rect 9493 24633 9505 24667
rect 9539 24664 9551 24667
rect 10042 24664 10048 24676
rect 9539 24636 10048 24664
rect 9539 24633 9551 24636
rect 9493 24627 9551 24633
rect 10042 24624 10048 24636
rect 10100 24624 10106 24676
rect 10612 24664 10640 24763
rect 11974 24760 11980 24772
rect 12032 24760 12038 24812
rect 12250 24760 12256 24812
rect 12308 24760 12314 24812
rect 12406 24800 12434 24840
rect 13078 24828 13084 24880
rect 13136 24828 13142 24880
rect 14936 24868 14964 24896
rect 13924 24840 14964 24868
rect 13817 24803 13875 24809
rect 13817 24800 13829 24803
rect 12406 24772 13829 24800
rect 13817 24769 13829 24772
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 10870 24692 10876 24744
rect 10928 24732 10934 24744
rect 10965 24735 11023 24741
rect 10965 24732 10977 24735
rect 10928 24704 10977 24732
rect 10928 24692 10934 24704
rect 10965 24701 10977 24704
rect 11011 24701 11023 24735
rect 10965 24695 11023 24701
rect 12069 24735 12127 24741
rect 12069 24701 12081 24735
rect 12115 24701 12127 24735
rect 12069 24695 12127 24701
rect 12161 24735 12219 24741
rect 12161 24701 12173 24735
rect 12207 24701 12219 24735
rect 12161 24695 12219 24701
rect 12437 24735 12495 24741
rect 12437 24701 12449 24735
rect 12483 24732 12495 24735
rect 12526 24732 12532 24744
rect 12483 24704 12532 24732
rect 12483 24701 12495 24704
rect 12437 24695 12495 24701
rect 10612 24636 11192 24664
rect 11164 24608 11192 24636
rect 9950 24556 9956 24608
rect 10008 24556 10014 24608
rect 10134 24556 10140 24608
rect 10192 24596 10198 24608
rect 10962 24596 10968 24608
rect 10192 24568 10968 24596
rect 10192 24556 10198 24568
rect 10962 24556 10968 24568
rect 11020 24556 11026 24608
rect 11146 24556 11152 24608
rect 11204 24556 11210 24608
rect 12084 24596 12112 24695
rect 12176 24664 12204 24695
rect 12526 24692 12532 24704
rect 12584 24692 12590 24744
rect 12618 24692 12624 24744
rect 12676 24692 12682 24744
rect 12710 24692 12716 24744
rect 12768 24692 12774 24744
rect 12805 24735 12863 24741
rect 12805 24701 12817 24735
rect 12851 24701 12863 24735
rect 12805 24695 12863 24701
rect 12897 24735 12955 24741
rect 12897 24701 12909 24735
rect 12943 24732 12955 24735
rect 13354 24732 13360 24744
rect 12943 24704 13360 24732
rect 12943 24701 12955 24704
rect 12897 24695 12955 24701
rect 12820 24664 12848 24695
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 13633 24735 13691 24741
rect 13633 24701 13645 24735
rect 13679 24701 13691 24735
rect 13633 24695 13691 24701
rect 13446 24664 13452 24676
rect 12176 24636 13452 24664
rect 13446 24624 13452 24636
rect 13504 24664 13510 24676
rect 13648 24664 13676 24695
rect 13504 24636 13676 24664
rect 13504 24624 13510 24636
rect 13924 24596 13952 24840
rect 14001 24803 14059 24809
rect 14001 24769 14013 24803
rect 14047 24800 14059 24803
rect 14274 24800 14280 24812
rect 14047 24772 14280 24800
rect 14047 24769 14059 24772
rect 14001 24763 14059 24769
rect 14274 24760 14280 24772
rect 14332 24760 14338 24812
rect 14642 24809 14648 24812
rect 14636 24763 14648 24809
rect 14642 24760 14648 24763
rect 14700 24760 14706 24812
rect 14369 24735 14427 24741
rect 14369 24701 14381 24735
rect 14415 24701 14427 24735
rect 15764 24732 15792 24896
rect 16040 24868 16068 24896
rect 16301 24871 16359 24877
rect 16301 24868 16313 24871
rect 16040 24840 16313 24868
rect 16301 24837 16313 24840
rect 16347 24837 16359 24871
rect 16301 24831 16359 24837
rect 16209 24803 16267 24809
rect 16209 24769 16221 24803
rect 16255 24800 16267 24803
rect 16408 24800 16436 24896
rect 17218 24828 17224 24880
rect 17276 24828 17282 24880
rect 18598 24877 18604 24880
rect 18592 24868 18604 24877
rect 18559 24840 18604 24868
rect 18592 24831 18604 24840
rect 18598 24828 18604 24831
rect 18656 24828 18662 24880
rect 19886 24828 19892 24880
rect 19944 24868 19950 24880
rect 21269 24871 21327 24877
rect 21269 24868 21281 24871
rect 19944 24840 21281 24868
rect 19944 24828 19950 24840
rect 21269 24837 21281 24840
rect 21315 24837 21327 24871
rect 21269 24831 21327 24837
rect 16255 24772 16436 24800
rect 16255 24769 16267 24772
rect 16209 24763 16267 24769
rect 16574 24760 16580 24812
rect 16632 24800 16638 24812
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 16632 24772 16681 24800
rect 16632 24760 16638 24772
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 16945 24803 17003 24809
rect 16945 24769 16957 24803
rect 16991 24800 17003 24803
rect 17497 24803 17555 24809
rect 16991 24772 17448 24800
rect 16991 24769 17003 24772
rect 16945 24763 17003 24769
rect 16485 24735 16543 24741
rect 16485 24732 16497 24735
rect 15764 24704 16497 24732
rect 14369 24695 14427 24701
rect 16485 24701 16497 24704
rect 16531 24701 16543 24735
rect 16485 24695 16543 24701
rect 17221 24735 17279 24741
rect 17221 24701 17233 24735
rect 17267 24701 17279 24735
rect 17420 24732 17448 24772
rect 17497 24769 17509 24803
rect 17543 24800 17555 24803
rect 17586 24800 17592 24812
rect 17543 24772 17592 24800
rect 17543 24769 17555 24772
rect 17497 24763 17555 24769
rect 17586 24760 17592 24772
rect 17644 24760 17650 24812
rect 18046 24760 18052 24812
rect 18104 24760 18110 24812
rect 19150 24800 19156 24812
rect 18340 24772 19156 24800
rect 18064 24732 18092 24760
rect 18340 24744 18368 24772
rect 19150 24760 19156 24772
rect 19208 24760 19214 24812
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24800 20499 24803
rect 21376 24800 21404 24908
rect 21979 24905 21991 24908
rect 22025 24905 22037 24939
rect 22370 24936 22376 24948
rect 21979 24899 22037 24905
rect 22204 24908 22376 24936
rect 22204 24877 22232 24908
rect 22370 24896 22376 24908
rect 22428 24896 22434 24948
rect 22189 24871 22247 24877
rect 20487 24772 21404 24800
rect 21499 24837 21557 24843
rect 21499 24803 21511 24837
rect 21545 24834 21557 24837
rect 22189 24837 22201 24871
rect 22235 24837 22247 24871
rect 21545 24806 21680 24834
rect 22189 24831 22247 24837
rect 21545 24803 21557 24806
rect 21499 24797 21557 24803
rect 20487 24769 20499 24772
rect 20441 24763 20499 24769
rect 17420 24704 18092 24732
rect 17221 24695 17279 24701
rect 12084 24568 13952 24596
rect 14384 24596 14412 24695
rect 14734 24596 14740 24608
rect 14384 24568 14740 24596
rect 14734 24556 14740 24568
rect 14792 24556 14798 24608
rect 16114 24556 16120 24608
rect 16172 24596 16178 24608
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16172 24568 16773 24596
rect 16172 24556 16178 24568
rect 16761 24565 16773 24568
rect 16807 24565 16819 24599
rect 17236 24596 17264 24695
rect 18322 24692 18328 24744
rect 18380 24692 18386 24744
rect 17402 24624 17408 24676
rect 17460 24624 17466 24676
rect 19705 24667 19763 24673
rect 19705 24633 19717 24667
rect 19751 24664 19763 24667
rect 20456 24664 20484 24763
rect 20530 24692 20536 24744
rect 20588 24732 20594 24744
rect 21085 24735 21143 24741
rect 21085 24732 21097 24735
rect 20588 24704 21097 24732
rect 20588 24692 20594 24704
rect 21085 24701 21097 24704
rect 21131 24732 21143 24735
rect 21174 24732 21180 24744
rect 21131 24704 21180 24732
rect 21131 24701 21143 24704
rect 21085 24695 21143 24701
rect 19751 24636 20484 24664
rect 19751 24633 19763 24636
rect 19705 24627 19763 24633
rect 18138 24596 18144 24608
rect 17236 24568 18144 24596
rect 16761 24559 16819 24565
rect 18138 24556 18144 24568
rect 18196 24556 18202 24608
rect 20530 24556 20536 24608
rect 20588 24556 20594 24608
rect 21100 24596 21128 24695
rect 21174 24692 21180 24704
rect 21232 24692 21238 24744
rect 21652 24664 21680 24806
rect 22373 24803 22431 24809
rect 22373 24800 22385 24803
rect 21928 24772 22385 24800
rect 21821 24667 21879 24673
rect 21821 24664 21833 24667
rect 21652 24636 21833 24664
rect 21821 24633 21833 24636
rect 21867 24633 21879 24667
rect 21821 24627 21879 24633
rect 21453 24599 21511 24605
rect 21453 24596 21465 24599
rect 21100 24568 21465 24596
rect 21453 24565 21465 24568
rect 21499 24565 21511 24599
rect 21453 24559 21511 24565
rect 21637 24599 21695 24605
rect 21637 24565 21649 24599
rect 21683 24596 21695 24599
rect 21928 24596 21956 24772
rect 22373 24769 22385 24772
rect 22419 24769 22431 24803
rect 22373 24763 22431 24769
rect 22278 24624 22284 24676
rect 22336 24664 22342 24676
rect 22557 24667 22615 24673
rect 22557 24664 22569 24667
rect 22336 24636 22569 24664
rect 22336 24624 22342 24636
rect 22557 24633 22569 24636
rect 22603 24664 22615 24667
rect 23014 24664 23020 24676
rect 22603 24636 23020 24664
rect 22603 24633 22615 24636
rect 22557 24627 22615 24633
rect 23014 24624 23020 24636
rect 23072 24624 23078 24676
rect 21683 24568 21956 24596
rect 21683 24565 21695 24568
rect 21637 24559 21695 24565
rect 22002 24556 22008 24608
rect 22060 24556 22066 24608
rect 1104 24506 26496 24528
rect 1104 24454 4124 24506
rect 4176 24454 4188 24506
rect 4240 24454 4252 24506
rect 4304 24454 4316 24506
rect 4368 24454 4380 24506
rect 4432 24454 10472 24506
rect 10524 24454 10536 24506
rect 10588 24454 10600 24506
rect 10652 24454 10664 24506
rect 10716 24454 10728 24506
rect 10780 24454 16820 24506
rect 16872 24454 16884 24506
rect 16936 24454 16948 24506
rect 17000 24454 17012 24506
rect 17064 24454 17076 24506
rect 17128 24454 23168 24506
rect 23220 24454 23232 24506
rect 23284 24454 23296 24506
rect 23348 24454 23360 24506
rect 23412 24454 23424 24506
rect 23476 24454 26496 24506
rect 1104 24432 26496 24454
rect 9122 24352 9128 24404
rect 9180 24392 9186 24404
rect 9309 24395 9367 24401
rect 9309 24392 9321 24395
rect 9180 24364 9321 24392
rect 9180 24352 9186 24364
rect 9309 24361 9321 24364
rect 9355 24361 9367 24395
rect 9309 24355 9367 24361
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 10045 24395 10103 24401
rect 10045 24392 10057 24395
rect 9732 24364 10057 24392
rect 9732 24352 9738 24364
rect 10045 24361 10057 24364
rect 10091 24392 10103 24395
rect 10134 24392 10140 24404
rect 10091 24364 10140 24392
rect 10091 24361 10103 24364
rect 10045 24355 10103 24361
rect 10134 24352 10140 24364
rect 10192 24352 10198 24404
rect 12894 24352 12900 24404
rect 12952 24352 12958 24404
rect 13078 24352 13084 24404
rect 13136 24352 13142 24404
rect 13354 24352 13360 24404
rect 13412 24352 13418 24404
rect 14642 24352 14648 24404
rect 14700 24352 14706 24404
rect 16114 24352 16120 24404
rect 16172 24352 16178 24404
rect 19061 24395 19119 24401
rect 19061 24361 19073 24395
rect 19107 24392 19119 24395
rect 19518 24392 19524 24404
rect 19107 24364 19524 24392
rect 19107 24361 19119 24364
rect 19061 24355 19119 24361
rect 19518 24352 19524 24364
rect 19576 24352 19582 24404
rect 19610 24352 19616 24404
rect 19668 24392 19674 24404
rect 19797 24395 19855 24401
rect 19797 24392 19809 24395
rect 19668 24364 19809 24392
rect 19668 24352 19674 24364
rect 19797 24361 19809 24364
rect 19843 24361 19855 24395
rect 19797 24355 19855 24361
rect 20530 24352 20536 24404
rect 20588 24352 20594 24404
rect 8757 24327 8815 24333
rect 8757 24293 8769 24327
rect 8803 24324 8815 24327
rect 9582 24324 9588 24336
rect 8803 24296 9588 24324
rect 8803 24293 8815 24296
rect 8757 24287 8815 24293
rect 9582 24284 9588 24296
rect 9640 24284 9646 24336
rect 9766 24284 9772 24336
rect 9824 24324 9830 24336
rect 10870 24324 10876 24336
rect 9824 24296 10876 24324
rect 9824 24284 9830 24296
rect 10870 24284 10876 24296
rect 10928 24284 10934 24336
rect 10962 24284 10968 24336
rect 11020 24324 11026 24336
rect 12161 24327 12219 24333
rect 12161 24324 12173 24327
rect 11020 24296 12173 24324
rect 11020 24284 11026 24296
rect 12161 24293 12173 24296
rect 12207 24324 12219 24327
rect 12526 24324 12532 24336
rect 12207 24296 12532 24324
rect 12207 24293 12219 24296
rect 12161 24287 12219 24293
rect 12526 24284 12532 24296
rect 12584 24284 12590 24336
rect 9600 24256 9628 24284
rect 10413 24259 10471 24265
rect 9600 24228 10364 24256
rect 7377 24191 7435 24197
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 8110 24188 8116 24200
rect 7423 24160 8116 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 8110 24148 8116 24160
rect 8168 24148 8174 24200
rect 9398 24148 9404 24200
rect 9456 24188 9462 24200
rect 9861 24191 9919 24197
rect 9861 24188 9873 24191
rect 9456 24160 9873 24188
rect 9456 24148 9462 24160
rect 9861 24157 9873 24160
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 10226 24148 10232 24200
rect 10284 24148 10290 24200
rect 10336 24188 10364 24228
rect 10413 24225 10425 24259
rect 10459 24256 10471 24259
rect 10459 24228 11192 24256
rect 10459 24225 10471 24228
rect 10413 24219 10471 24225
rect 11164 24200 11192 24228
rect 11790 24216 11796 24268
rect 11848 24216 11854 24268
rect 10505 24191 10563 24197
rect 10505 24188 10517 24191
rect 10336 24160 10517 24188
rect 10505 24157 10517 24160
rect 10551 24157 10563 24191
rect 10505 24151 10563 24157
rect 11146 24148 11152 24200
rect 11204 24148 11210 24200
rect 12618 24148 12624 24200
rect 12676 24148 12682 24200
rect 12897 24191 12955 24197
rect 12897 24157 12909 24191
rect 12943 24188 12955 24191
rect 13096 24188 13124 24352
rect 13372 24324 13400 24352
rect 16298 24324 16304 24336
rect 13372 24296 16304 24324
rect 16298 24284 16304 24296
rect 16356 24284 16362 24336
rect 19702 24324 19708 24336
rect 18892 24296 19708 24324
rect 13998 24216 14004 24268
rect 14056 24216 14062 24268
rect 15749 24259 15807 24265
rect 15749 24225 15761 24259
rect 15795 24256 15807 24259
rect 16206 24256 16212 24268
rect 15795 24228 16212 24256
rect 15795 24225 15807 24228
rect 15749 24219 15807 24225
rect 16206 24216 16212 24228
rect 16264 24216 16270 24268
rect 16482 24216 16488 24268
rect 16540 24216 16546 24268
rect 12943 24160 13124 24188
rect 14016 24188 14044 24216
rect 14829 24191 14887 24197
rect 14829 24188 14841 24191
rect 14016 24160 14841 24188
rect 12943 24157 12955 24160
rect 12897 24151 12955 24157
rect 14829 24157 14841 24160
rect 14875 24157 14887 24191
rect 14829 24151 14887 24157
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 16500 24188 16528 24216
rect 18892 24197 18920 24296
rect 19702 24284 19708 24296
rect 19760 24284 19766 24336
rect 19429 24259 19487 24265
rect 19429 24225 19441 24259
rect 19475 24256 19487 24259
rect 19518 24256 19524 24268
rect 19475 24228 19524 24256
rect 19475 24225 19487 24228
rect 19429 24219 19487 24225
rect 19518 24216 19524 24228
rect 19576 24216 19582 24268
rect 20548 24256 20576 24352
rect 19720 24228 20576 24256
rect 19720 24197 19748 24228
rect 20622 24216 20628 24268
rect 20680 24216 20686 24268
rect 23201 24259 23259 24265
rect 23201 24256 23213 24259
rect 22388 24228 23213 24256
rect 15979 24160 16528 24188
rect 18877 24191 18935 24197
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 18877 24157 18889 24191
rect 18923 24157 18935 24191
rect 18877 24151 18935 24157
rect 19061 24191 19119 24197
rect 19061 24157 19073 24191
rect 19107 24188 19119 24191
rect 19613 24191 19671 24197
rect 19107 24160 19472 24188
rect 19107 24157 19119 24160
rect 19061 24151 19119 24157
rect 7644 24123 7702 24129
rect 7644 24089 7656 24123
rect 7690 24120 7702 24123
rect 7742 24120 7748 24132
rect 7690 24092 7748 24120
rect 7690 24089 7702 24092
rect 7644 24083 7702 24089
rect 7742 24080 7748 24092
rect 7800 24080 7806 24132
rect 12710 24120 12716 24132
rect 12406 24092 12716 24120
rect 12253 24055 12311 24061
rect 12253 24021 12265 24055
rect 12299 24052 12311 24055
rect 12406 24052 12434 24092
rect 12710 24080 12716 24092
rect 12768 24120 12774 24132
rect 15948 24120 15976 24151
rect 19444 24129 19472 24160
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 12768 24092 15976 24120
rect 19429 24123 19487 24129
rect 12768 24080 12774 24092
rect 19429 24089 19441 24123
rect 19475 24089 19487 24123
rect 19628 24120 19656 24151
rect 19794 24148 19800 24200
rect 19852 24188 19858 24200
rect 19981 24191 20039 24197
rect 19981 24188 19993 24191
rect 19852 24160 19993 24188
rect 19852 24148 19858 24160
rect 19981 24157 19993 24160
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20070 24148 20076 24200
rect 20128 24148 20134 24200
rect 20165 24191 20223 24197
rect 20165 24157 20177 24191
rect 20211 24157 20223 24191
rect 20165 24151 20223 24157
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24188 20315 24191
rect 20640 24188 20668 24216
rect 22388 24200 22416 24228
rect 23201 24225 23213 24228
rect 23247 24225 23259 24259
rect 23201 24219 23259 24225
rect 20303 24160 20668 24188
rect 20303 24157 20315 24160
rect 20257 24151 20315 24157
rect 19812 24120 19840 24148
rect 19628 24092 19840 24120
rect 19429 24083 19487 24089
rect 19886 24080 19892 24132
rect 19944 24120 19950 24132
rect 20180 24120 20208 24151
rect 19944 24092 20208 24120
rect 19944 24080 19950 24092
rect 12299 24024 12434 24052
rect 12299 24021 12311 24024
rect 12253 24015 12311 24021
rect 19794 24012 19800 24064
rect 19852 24052 19858 24064
rect 20272 24052 20300 24151
rect 22370 24148 22376 24200
rect 22428 24148 22434 24200
rect 23014 24148 23020 24200
rect 23072 24148 23078 24200
rect 23106 24148 23112 24200
rect 23164 24148 23170 24200
rect 23290 24148 23296 24200
rect 23348 24148 23354 24200
rect 23385 24191 23443 24197
rect 23385 24157 23397 24191
rect 23431 24157 23443 24191
rect 23385 24151 23443 24157
rect 23032 24120 23060 24148
rect 23400 24120 23428 24151
rect 26142 24148 26148 24200
rect 26200 24148 26206 24200
rect 22066 24092 23428 24120
rect 22066 24052 22094 24092
rect 19852 24024 22094 24052
rect 19852 24012 19858 24024
rect 22462 24012 22468 24064
rect 22520 24052 22526 24064
rect 22925 24055 22983 24061
rect 22925 24052 22937 24055
rect 22520 24024 22937 24052
rect 22520 24012 22526 24024
rect 22925 24021 22937 24024
rect 22971 24021 22983 24055
rect 22925 24015 22983 24021
rect 1104 23962 26656 23984
rect 1104 23910 7298 23962
rect 7350 23910 7362 23962
rect 7414 23910 7426 23962
rect 7478 23910 7490 23962
rect 7542 23910 7554 23962
rect 7606 23910 13646 23962
rect 13698 23910 13710 23962
rect 13762 23910 13774 23962
rect 13826 23910 13838 23962
rect 13890 23910 13902 23962
rect 13954 23910 19994 23962
rect 20046 23910 20058 23962
rect 20110 23910 20122 23962
rect 20174 23910 20186 23962
rect 20238 23910 20250 23962
rect 20302 23910 26342 23962
rect 26394 23910 26406 23962
rect 26458 23910 26470 23962
rect 26522 23910 26534 23962
rect 26586 23910 26598 23962
rect 26650 23910 26656 23962
rect 1104 23888 26656 23910
rect 7742 23808 7748 23860
rect 7800 23808 7806 23860
rect 9493 23851 9551 23857
rect 9493 23817 9505 23851
rect 9539 23817 9551 23851
rect 9493 23811 9551 23817
rect 9677 23851 9735 23857
rect 9677 23817 9689 23851
rect 9723 23848 9735 23851
rect 9766 23848 9772 23860
rect 9723 23820 9772 23848
rect 9723 23817 9735 23820
rect 9677 23811 9735 23817
rect 9508 23780 9536 23811
rect 9766 23808 9772 23820
rect 9824 23808 9830 23860
rect 10042 23808 10048 23860
rect 10100 23808 10106 23860
rect 22097 23851 22155 23857
rect 22097 23817 22109 23851
rect 22143 23848 22155 23851
rect 22143 23820 22784 23848
rect 22143 23817 22155 23820
rect 22097 23811 22155 23817
rect 7944 23752 9536 23780
rect 7944 23721 7972 23752
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 8021 23715 8079 23721
rect 8021 23681 8033 23715
rect 8067 23712 8079 23715
rect 8110 23712 8116 23724
rect 8067 23684 8116 23712
rect 8067 23681 8079 23684
rect 8021 23675 8079 23681
rect 8110 23672 8116 23684
rect 8168 23672 8174 23724
rect 8288 23715 8346 23721
rect 8288 23681 8300 23715
rect 8334 23712 8346 23715
rect 10060 23712 10088 23808
rect 22462 23780 22468 23792
rect 22204 23752 22468 23780
rect 10137 23715 10195 23721
rect 10137 23712 10149 23715
rect 8334 23684 9260 23712
rect 10060 23684 10149 23712
rect 8334 23681 8346 23684
rect 8288 23675 8346 23681
rect 9232 23644 9260 23684
rect 10137 23681 10149 23684
rect 10183 23681 10195 23715
rect 10137 23675 10195 23681
rect 10318 23672 10324 23724
rect 10376 23672 10382 23724
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23712 14519 23715
rect 16022 23712 16028 23724
rect 14507 23684 16028 23712
rect 14507 23681 14519 23684
rect 14461 23675 14519 23681
rect 16022 23672 16028 23684
rect 16080 23672 16086 23724
rect 22204 23721 22232 23752
rect 22462 23740 22468 23752
rect 22520 23740 22526 23792
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 22189 23715 22247 23721
rect 22189 23681 22201 23715
rect 22235 23681 22247 23715
rect 22189 23675 22247 23681
rect 10229 23647 10287 23653
rect 10229 23644 10241 23647
rect 9232 23616 10241 23644
rect 10229 23613 10241 23616
rect 10275 23613 10287 23647
rect 10336 23644 10364 23672
rect 10336 23616 12434 23644
rect 10229 23607 10287 23613
rect 9950 23576 9956 23588
rect 9692 23548 9956 23576
rect 9398 23468 9404 23520
rect 9456 23468 9462 23520
rect 9692 23517 9720 23548
rect 9950 23536 9956 23548
rect 10008 23536 10014 23588
rect 10045 23579 10103 23585
rect 10045 23545 10057 23579
rect 10091 23576 10103 23579
rect 10134 23576 10140 23588
rect 10091 23548 10140 23576
rect 10091 23545 10103 23548
rect 10045 23539 10103 23545
rect 10134 23536 10140 23548
rect 10192 23536 10198 23588
rect 12406 23576 12434 23616
rect 14550 23604 14556 23656
rect 14608 23644 14614 23656
rect 14829 23647 14887 23653
rect 14829 23644 14841 23647
rect 14608 23616 14841 23644
rect 14608 23604 14614 23616
rect 14829 23613 14841 23616
rect 14875 23613 14887 23647
rect 14829 23607 14887 23613
rect 15378 23604 15384 23656
rect 15436 23604 15442 23656
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23644 19763 23647
rect 20346 23644 20352 23656
rect 19751 23616 20352 23644
rect 19751 23613 19763 23616
rect 19705 23607 19763 23613
rect 20346 23604 20352 23616
rect 20404 23604 20410 23656
rect 22020 23644 22048 23675
rect 22278 23672 22284 23724
rect 22336 23672 22342 23724
rect 22370 23672 22376 23724
rect 22428 23672 22434 23724
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23712 22615 23715
rect 22756 23712 22784 23820
rect 23290 23808 23296 23860
rect 23348 23848 23354 23860
rect 23566 23848 23572 23860
rect 23348 23820 23572 23848
rect 23348 23808 23354 23820
rect 23566 23808 23572 23820
rect 23624 23848 23630 23860
rect 24121 23851 24179 23857
rect 24121 23848 24133 23851
rect 23624 23820 24133 23848
rect 23624 23808 23630 23820
rect 24121 23817 24133 23820
rect 24167 23848 24179 23851
rect 24167 23820 24808 23848
rect 24167 23817 24179 23820
rect 24121 23811 24179 23817
rect 24780 23724 24808 23820
rect 22997 23715 23055 23721
rect 22997 23712 23009 23715
rect 22603 23684 22692 23712
rect 22756 23684 23009 23712
rect 22603 23681 22615 23684
rect 22557 23675 22615 23681
rect 22020 23616 22094 23644
rect 15470 23576 15476 23588
rect 12406 23548 15476 23576
rect 15470 23536 15476 23548
rect 15528 23536 15534 23588
rect 22066 23576 22094 23616
rect 22557 23579 22615 23585
rect 22557 23576 22569 23579
rect 22066 23548 22569 23576
rect 22557 23545 22569 23548
rect 22603 23545 22615 23579
rect 22557 23539 22615 23545
rect 9677 23511 9735 23517
rect 9677 23477 9689 23511
rect 9723 23477 9735 23511
rect 9677 23471 9735 23477
rect 14642 23468 14648 23520
rect 14700 23468 14706 23520
rect 15102 23468 15108 23520
rect 15160 23508 15166 23520
rect 18138 23508 18144 23520
rect 15160 23480 18144 23508
rect 15160 23468 15166 23480
rect 18138 23468 18144 23480
rect 18196 23468 18202 23520
rect 19058 23468 19064 23520
rect 19116 23468 19122 23520
rect 22664 23508 22692 23684
rect 22997 23681 23009 23684
rect 23043 23681 23055 23715
rect 22997 23675 23055 23681
rect 24762 23672 24768 23724
rect 24820 23672 24826 23724
rect 22738 23604 22744 23656
rect 22796 23604 22802 23656
rect 23860 23548 24256 23576
rect 23860 23508 23888 23548
rect 24228 23517 24256 23548
rect 22664 23480 23888 23508
rect 24213 23511 24271 23517
rect 24213 23477 24225 23511
rect 24259 23477 24271 23511
rect 24213 23471 24271 23477
rect 1104 23418 26496 23440
rect 1104 23366 4124 23418
rect 4176 23366 4188 23418
rect 4240 23366 4252 23418
rect 4304 23366 4316 23418
rect 4368 23366 4380 23418
rect 4432 23366 10472 23418
rect 10524 23366 10536 23418
rect 10588 23366 10600 23418
rect 10652 23366 10664 23418
rect 10716 23366 10728 23418
rect 10780 23366 16820 23418
rect 16872 23366 16884 23418
rect 16936 23366 16948 23418
rect 17000 23366 17012 23418
rect 17064 23366 17076 23418
rect 17128 23366 23168 23418
rect 23220 23366 23232 23418
rect 23284 23366 23296 23418
rect 23348 23366 23360 23418
rect 23412 23366 23424 23418
rect 23476 23366 26496 23418
rect 1104 23344 26496 23366
rect 10137 23307 10195 23313
rect 10137 23273 10149 23307
rect 10183 23273 10195 23307
rect 10137 23267 10195 23273
rect 10321 23307 10379 23313
rect 10321 23273 10333 23307
rect 10367 23304 10379 23307
rect 11333 23307 11391 23313
rect 11333 23304 11345 23307
rect 10367 23276 11345 23304
rect 10367 23273 10379 23276
rect 10321 23267 10379 23273
rect 11333 23273 11345 23276
rect 11379 23273 11391 23307
rect 13633 23307 13691 23313
rect 13633 23304 13645 23307
rect 11333 23267 11391 23273
rect 11532 23276 13645 23304
rect 10042 23236 10048 23248
rect 9324 23208 10048 23236
rect 9324 23177 9352 23208
rect 10042 23196 10048 23208
rect 10100 23196 10106 23248
rect 10152 23236 10180 23267
rect 10152 23208 10732 23236
rect 9309 23171 9367 23177
rect 9309 23137 9321 23171
rect 9355 23137 9367 23171
rect 9309 23131 9367 23137
rect 9398 23128 9404 23180
rect 9456 23168 9462 23180
rect 10152 23168 10180 23208
rect 9456 23140 10180 23168
rect 9456 23128 9462 23140
rect 10226 23128 10232 23180
rect 10284 23168 10290 23180
rect 10413 23171 10471 23177
rect 10413 23168 10425 23171
rect 10284 23140 10425 23168
rect 10284 23128 10290 23140
rect 10413 23137 10425 23140
rect 10459 23137 10471 23171
rect 10413 23131 10471 23137
rect 9217 23103 9275 23109
rect 9217 23069 9229 23103
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23100 9551 23103
rect 9582 23100 9588 23112
rect 9539 23072 9588 23100
rect 9539 23069 9551 23072
rect 9493 23063 9551 23069
rect 9232 23032 9260 23063
rect 9582 23060 9588 23072
rect 9640 23100 9646 23112
rect 10704 23109 10732 23208
rect 11146 23196 11152 23248
rect 11204 23196 11210 23248
rect 10965 23171 11023 23177
rect 10965 23137 10977 23171
rect 11011 23168 11023 23171
rect 11532 23168 11560 23276
rect 13633 23273 13645 23276
rect 13679 23273 13691 23307
rect 13633 23267 13691 23273
rect 14274 23264 14280 23316
rect 14332 23304 14338 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 14332 23276 14473 23304
rect 14332 23264 14338 23276
rect 14461 23273 14473 23276
rect 14507 23304 14519 23307
rect 15102 23304 15108 23316
rect 14507 23276 15108 23304
rect 14507 23273 14519 23276
rect 14461 23267 14519 23273
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 16945 23307 17003 23313
rect 16945 23273 16957 23307
rect 16991 23304 17003 23307
rect 20809 23307 20867 23313
rect 16991 23276 17448 23304
rect 16991 23273 17003 23276
rect 16945 23267 17003 23273
rect 13078 23196 13084 23248
rect 13136 23236 13142 23248
rect 13725 23239 13783 23245
rect 13725 23236 13737 23239
rect 13136 23208 13737 23236
rect 13136 23196 13142 23208
rect 13725 23205 13737 23208
rect 13771 23205 13783 23239
rect 13725 23199 13783 23205
rect 13817 23171 13875 23177
rect 11011 23140 11560 23168
rect 11808 23140 12480 23168
rect 11011 23137 11023 23140
rect 10965 23131 11023 23137
rect 11164 23112 11192 23140
rect 11808 23112 11836 23140
rect 9769 23103 9827 23109
rect 9769 23100 9781 23103
rect 9640 23072 9781 23100
rect 9640 23060 9646 23072
rect 9769 23069 9781 23072
rect 9815 23100 9827 23103
rect 10689 23103 10747 23109
rect 9815 23072 10272 23100
rect 9815 23069 9827 23072
rect 9769 23063 9827 23069
rect 9950 23032 9956 23044
rect 9232 23004 9956 23032
rect 9950 22992 9956 23004
rect 10008 23032 10014 23044
rect 10137 23035 10195 23041
rect 10137 23032 10149 23035
rect 10008 23004 10149 23032
rect 10008 22992 10014 23004
rect 10137 23001 10149 23004
rect 10183 23001 10195 23035
rect 10244 23032 10272 23072
rect 10689 23069 10701 23103
rect 10735 23069 10747 23103
rect 10689 23063 10747 23069
rect 11146 23060 11152 23112
rect 11204 23060 11210 23112
rect 11698 23060 11704 23112
rect 11756 23060 11762 23112
rect 11790 23060 11796 23112
rect 11848 23060 11854 23112
rect 12158 23060 12164 23112
rect 12216 23060 12222 23112
rect 12452 23109 12480 23140
rect 13817 23137 13829 23171
rect 13863 23168 13875 23171
rect 14292 23168 14320 23264
rect 13863 23140 14320 23168
rect 13863 23137 13875 23140
rect 13817 23131 13875 23137
rect 12437 23103 12495 23109
rect 12437 23069 12449 23103
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 12621 23103 12679 23109
rect 12621 23069 12633 23103
rect 12667 23100 12679 23103
rect 12805 23103 12863 23109
rect 12805 23100 12817 23103
rect 12667 23072 12817 23100
rect 12667 23069 12679 23072
rect 12621 23063 12679 23069
rect 12805 23069 12817 23072
rect 12851 23069 12863 23103
rect 12805 23063 12863 23069
rect 13357 23103 13415 23109
rect 13357 23069 13369 23103
rect 13403 23069 13415 23103
rect 13357 23063 13415 23069
rect 10781 23035 10839 23041
rect 10781 23032 10793 23035
rect 10244 23004 10793 23032
rect 10137 22995 10195 23001
rect 10781 23001 10793 23004
rect 10827 23001 10839 23035
rect 10781 22995 10839 23001
rect 11333 23035 11391 23041
rect 11333 23001 11345 23035
rect 11379 23032 11391 23035
rect 12986 23032 12992 23044
rect 11379 23004 12992 23032
rect 11379 23001 11391 23004
rect 11333 22995 11391 23001
rect 9674 22924 9680 22976
rect 9732 22924 9738 22976
rect 10152 22964 10180 22995
rect 12986 22992 12992 23004
rect 13044 23032 13050 23044
rect 13372 23032 13400 23063
rect 13538 23060 13544 23112
rect 13596 23060 13602 23112
rect 14182 23060 14188 23112
rect 14240 23100 14246 23112
rect 14829 23103 14887 23109
rect 14829 23100 14841 23103
rect 14240 23072 14841 23100
rect 14240 23060 14246 23072
rect 14829 23069 14841 23072
rect 14875 23069 14887 23103
rect 14829 23063 14887 23069
rect 13044 23004 13400 23032
rect 14844 23032 14872 23063
rect 14918 23060 14924 23112
rect 14976 23060 14982 23112
rect 15562 23060 15568 23112
rect 15620 23060 15626 23112
rect 15930 23060 15936 23112
rect 15988 23060 15994 23112
rect 17420 23109 17448 23276
rect 20809 23273 20821 23307
rect 20855 23304 20867 23307
rect 20898 23304 20904 23316
rect 20855 23276 20904 23304
rect 20855 23273 20867 23276
rect 20809 23267 20867 23273
rect 20898 23264 20904 23276
rect 20956 23264 20962 23316
rect 23290 23304 23296 23316
rect 22664 23276 23296 23304
rect 22664 23248 22692 23276
rect 23290 23264 23296 23276
rect 23348 23304 23354 23316
rect 23348 23276 24256 23304
rect 23348 23264 23354 23276
rect 17957 23239 18015 23245
rect 17957 23205 17969 23239
rect 18003 23236 18015 23239
rect 18233 23239 18291 23245
rect 18233 23236 18245 23239
rect 18003 23208 18245 23236
rect 18003 23205 18015 23208
rect 17957 23199 18015 23205
rect 18233 23205 18245 23208
rect 18279 23205 18291 23239
rect 19518 23236 19524 23248
rect 18233 23199 18291 23205
rect 18340 23208 19524 23236
rect 18340 23168 18368 23208
rect 19518 23196 19524 23208
rect 19576 23236 19582 23248
rect 21910 23236 21916 23248
rect 19576 23208 21916 23236
rect 19576 23196 19582 23208
rect 21910 23196 21916 23208
rect 21968 23196 21974 23248
rect 22278 23196 22284 23248
rect 22336 23236 22342 23248
rect 22646 23236 22652 23248
rect 22336 23208 22652 23236
rect 22336 23196 22342 23208
rect 22646 23196 22652 23208
rect 22704 23196 22710 23248
rect 17788 23140 18092 23168
rect 17788 23109 17816 23140
rect 18064 23112 18092 23140
rect 18156 23140 18368 23168
rect 18601 23171 18659 23177
rect 18156 23112 18184 23140
rect 18601 23137 18613 23171
rect 18647 23168 18659 23171
rect 19797 23171 19855 23177
rect 19797 23168 19809 23171
rect 18647 23140 19809 23168
rect 18647 23137 18659 23140
rect 18601 23131 18659 23137
rect 19797 23137 19809 23140
rect 19843 23137 19855 23171
rect 19797 23131 19855 23137
rect 19886 23128 19892 23180
rect 19944 23168 19950 23180
rect 20257 23171 20315 23177
rect 20257 23168 20269 23171
rect 19944 23140 20269 23168
rect 19944 23128 19950 23140
rect 20257 23137 20269 23140
rect 20303 23168 20315 23171
rect 20993 23171 21051 23177
rect 20993 23168 21005 23171
rect 20303 23140 21005 23168
rect 20303 23137 20315 23140
rect 20257 23131 20315 23137
rect 20993 23137 21005 23140
rect 21039 23168 21051 23171
rect 24026 23168 24032 23180
rect 21039 23140 22508 23168
rect 21039 23137 21051 23140
rect 20993 23131 21051 23137
rect 17405 23103 17463 23109
rect 17405 23069 17417 23103
rect 17451 23100 17463 23103
rect 17773 23103 17831 23109
rect 17773 23100 17785 23103
rect 17451 23072 17785 23100
rect 17451 23069 17463 23072
rect 17405 23063 17463 23069
rect 17773 23069 17785 23072
rect 17819 23069 17831 23103
rect 17773 23063 17831 23069
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 16482 23032 16488 23044
rect 14844 23004 16488 23032
rect 13044 22992 13050 23004
rect 16482 22992 16488 23004
rect 16540 23032 16546 23044
rect 17129 23035 17187 23041
rect 17129 23032 17141 23035
rect 16540 23004 17141 23032
rect 16540 22992 16546 23004
rect 17129 23001 17141 23004
rect 17175 23001 17187 23035
rect 17129 22995 17187 23001
rect 17678 22992 17684 23044
rect 17736 23032 17742 23044
rect 17972 23032 18000 23063
rect 18046 23060 18052 23112
rect 18104 23060 18110 23112
rect 18138 23060 18144 23112
rect 18196 23060 18202 23112
rect 18230 23060 18236 23112
rect 18288 23100 18294 23112
rect 18325 23103 18383 23109
rect 18325 23100 18337 23103
rect 18288 23072 18337 23100
rect 18288 23060 18294 23072
rect 18325 23069 18337 23072
rect 18371 23069 18383 23103
rect 18325 23063 18383 23069
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23100 18475 23103
rect 19058 23100 19064 23112
rect 18463 23072 19064 23100
rect 18463 23069 18475 23072
rect 18417 23063 18475 23069
rect 19058 23060 19064 23072
rect 19116 23060 19122 23112
rect 20346 23060 20352 23112
rect 20404 23100 20410 23112
rect 20806 23100 20812 23112
rect 20404 23072 20812 23100
rect 20404 23060 20410 23072
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 21634 23060 21640 23112
rect 21692 23060 21698 23112
rect 21730 23103 21788 23109
rect 21730 23069 21742 23103
rect 21776 23069 21788 23103
rect 21730 23063 21788 23069
rect 17736 23004 18000 23032
rect 21545 23035 21603 23041
rect 17736 22992 17742 23004
rect 21545 23001 21557 23035
rect 21591 23032 21603 23035
rect 21744 23032 21772 23063
rect 22094 23060 22100 23112
rect 22152 23109 22158 23112
rect 22152 23100 22160 23109
rect 22152 23072 22197 23100
rect 22152 23063 22160 23072
rect 22152 23060 22158 23063
rect 22278 23060 22284 23112
rect 22336 23100 22342 23112
rect 22373 23103 22431 23109
rect 22373 23100 22385 23103
rect 22336 23072 22385 23100
rect 22336 23060 22342 23072
rect 22373 23069 22385 23072
rect 22419 23069 22431 23103
rect 22373 23063 22431 23069
rect 21591 23004 21772 23032
rect 21591 23001 21603 23004
rect 21545 22995 21603 23001
rect 21910 22992 21916 23044
rect 21968 22992 21974 23044
rect 22005 23035 22063 23041
rect 22005 23001 22017 23035
rect 22051 23032 22063 23035
rect 22186 23032 22192 23044
rect 22051 23004 22192 23032
rect 22051 23001 22063 23004
rect 22005 22995 22063 23001
rect 22186 22992 22192 23004
rect 22244 22992 22250 23044
rect 22480 23032 22508 23140
rect 23676 23140 24032 23168
rect 22554 23060 22560 23112
rect 22612 23060 22618 23112
rect 22649 23103 22707 23109
rect 22649 23069 22661 23103
rect 22695 23100 22707 23103
rect 22738 23100 22744 23112
rect 22695 23072 22744 23100
rect 22695 23069 22707 23072
rect 22649 23063 22707 23069
rect 22738 23060 22744 23072
rect 22796 23100 22802 23112
rect 23676 23100 23704 23140
rect 24026 23128 24032 23140
rect 24084 23128 24090 23180
rect 22796 23072 23704 23100
rect 24228 23100 24256 23276
rect 24762 23128 24768 23180
rect 24820 23128 24826 23180
rect 24581 23103 24639 23109
rect 24581 23100 24593 23103
rect 24228 23072 24593 23100
rect 22796 23060 22802 23072
rect 24581 23069 24593 23072
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 24670 23060 24676 23112
rect 24728 23060 24734 23112
rect 24857 23103 24915 23109
rect 24857 23069 24869 23103
rect 24903 23069 24915 23103
rect 24857 23063 24915 23069
rect 22922 23041 22928 23044
rect 22480 23004 22876 23032
rect 22848 22976 22876 23004
rect 22916 22995 22928 23041
rect 22922 22992 22928 22995
rect 22980 22992 22986 23044
rect 24872 23032 24900 23063
rect 25314 23060 25320 23112
rect 25372 23060 25378 23112
rect 24946 23032 24952 23044
rect 24044 23004 24952 23032
rect 10597 22967 10655 22973
rect 10597 22964 10609 22967
rect 10152 22936 10609 22964
rect 10597 22933 10609 22936
rect 10643 22933 10655 22967
rect 10597 22927 10655 22933
rect 11974 22924 11980 22976
rect 12032 22924 12038 22976
rect 15010 22924 15016 22976
rect 15068 22924 15074 22976
rect 16206 22924 16212 22976
rect 16264 22964 16270 22976
rect 16577 22967 16635 22973
rect 16577 22964 16589 22967
rect 16264 22936 16589 22964
rect 16264 22924 16270 22936
rect 16577 22933 16589 22936
rect 16623 22933 16635 22967
rect 16577 22927 16635 22933
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 16761 22967 16819 22973
rect 16761 22964 16773 22967
rect 16724 22936 16773 22964
rect 16724 22924 16730 22936
rect 16761 22933 16773 22936
rect 16807 22933 16819 22967
rect 16761 22927 16819 22933
rect 16929 22967 16987 22973
rect 16929 22933 16941 22967
rect 16975 22964 16987 22967
rect 17402 22964 17408 22976
rect 16975 22936 17408 22964
rect 16975 22933 16987 22936
rect 16929 22927 16987 22933
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 17497 22967 17555 22973
rect 17497 22933 17509 22967
rect 17543 22964 17555 22967
rect 17954 22964 17960 22976
rect 17543 22936 17960 22964
rect 17543 22933 17555 22936
rect 17497 22927 17555 22933
rect 17954 22924 17960 22936
rect 18012 22924 18018 22976
rect 19242 22924 19248 22976
rect 19300 22924 19306 22976
rect 20438 22924 20444 22976
rect 20496 22924 20502 22976
rect 22278 22924 22284 22976
rect 22336 22924 22342 22976
rect 22462 22924 22468 22976
rect 22520 22924 22526 22976
rect 22830 22924 22836 22976
rect 22888 22924 22894 22976
rect 23658 22924 23664 22976
rect 23716 22964 23722 22976
rect 24044 22973 24072 23004
rect 24946 22992 24952 23004
rect 25004 22992 25010 23044
rect 24029 22967 24087 22973
rect 24029 22964 24041 22967
rect 23716 22936 24041 22964
rect 23716 22924 23722 22936
rect 24029 22933 24041 22936
rect 24075 22933 24087 22967
rect 24029 22927 24087 22933
rect 24118 22924 24124 22976
rect 24176 22964 24182 22976
rect 24397 22967 24455 22973
rect 24397 22964 24409 22967
rect 24176 22936 24409 22964
rect 24176 22924 24182 22936
rect 24397 22933 24409 22936
rect 24443 22933 24455 22967
rect 24397 22927 24455 22933
rect 25130 22924 25136 22976
rect 25188 22924 25194 22976
rect 1104 22874 26656 22896
rect 1104 22822 7298 22874
rect 7350 22822 7362 22874
rect 7414 22822 7426 22874
rect 7478 22822 7490 22874
rect 7542 22822 7554 22874
rect 7606 22822 13646 22874
rect 13698 22822 13710 22874
rect 13762 22822 13774 22874
rect 13826 22822 13838 22874
rect 13890 22822 13902 22874
rect 13954 22822 19994 22874
rect 20046 22822 20058 22874
rect 20110 22822 20122 22874
rect 20174 22822 20186 22874
rect 20238 22822 20250 22874
rect 20302 22822 26342 22874
rect 26394 22822 26406 22874
rect 26458 22822 26470 22874
rect 26522 22822 26534 22874
rect 26586 22822 26598 22874
rect 26650 22822 26656 22874
rect 1104 22800 26656 22822
rect 9674 22720 9680 22772
rect 9732 22720 9738 22772
rect 9950 22720 9956 22772
rect 10008 22720 10014 22772
rect 11146 22720 11152 22772
rect 11204 22720 11210 22772
rect 11333 22763 11391 22769
rect 11333 22729 11345 22763
rect 11379 22760 11391 22763
rect 11790 22760 11796 22772
rect 11379 22732 11796 22760
rect 11379 22729 11391 22732
rect 11333 22723 11391 22729
rect 11790 22720 11796 22732
rect 11848 22720 11854 22772
rect 11974 22720 11980 22772
rect 12032 22720 12038 22772
rect 12158 22720 12164 22772
rect 12216 22760 12222 22772
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 12216 22732 13093 22760
rect 12216 22720 12222 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 13081 22723 13139 22729
rect 13354 22720 13360 22772
rect 13412 22760 13418 22772
rect 15105 22763 15163 22769
rect 13412 22732 13676 22760
rect 13412 22720 13418 22732
rect 9692 22692 9720 22720
rect 10689 22695 10747 22701
rect 10689 22692 10701 22695
rect 9692 22664 10701 22692
rect 10689 22661 10701 22664
rect 10735 22661 10747 22695
rect 10689 22655 10747 22661
rect 8110 22584 8116 22636
rect 8168 22624 8174 22636
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 8168 22596 8585 22624
rect 8168 22584 8174 22596
rect 8573 22593 8585 22596
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 8840 22627 8898 22633
rect 8840 22593 8852 22627
rect 8886 22624 8898 22627
rect 9306 22624 9312 22636
rect 8886 22596 9312 22624
rect 8886 22593 8898 22596
rect 8840 22587 8898 22593
rect 9306 22584 9312 22596
rect 9364 22584 9370 22636
rect 9950 22584 9956 22636
rect 10008 22624 10014 22636
rect 11164 22633 11192 22720
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 10008 22596 10241 22624
rect 10008 22584 10014 22596
rect 10229 22593 10241 22596
rect 10275 22593 10287 22627
rect 10229 22587 10287 22593
rect 10413 22627 10471 22633
rect 10413 22593 10425 22627
rect 10459 22624 10471 22627
rect 11149 22627 11207 22633
rect 11149 22624 11161 22627
rect 10459 22596 11161 22624
rect 10459 22593 10471 22596
rect 10413 22587 10471 22593
rect 11149 22593 11161 22596
rect 11195 22593 11207 22627
rect 11149 22587 11207 22593
rect 11238 22584 11244 22636
rect 11296 22624 11302 22636
rect 11609 22627 11667 22633
rect 11609 22624 11621 22627
rect 11296 22596 11621 22624
rect 11296 22584 11302 22596
rect 11609 22593 11621 22596
rect 11655 22593 11667 22627
rect 11609 22587 11667 22593
rect 11698 22584 11704 22636
rect 11756 22584 11762 22636
rect 11808 22624 11836 22720
rect 11876 22695 11934 22701
rect 11876 22661 11888 22695
rect 11922 22692 11934 22695
rect 11992 22692 12020 22720
rect 11922 22664 12020 22692
rect 11922 22661 11934 22664
rect 11876 22655 11934 22661
rect 12526 22652 12532 22704
rect 12584 22692 12590 22704
rect 13446 22692 13452 22704
rect 12584 22664 13452 22692
rect 12584 22652 12590 22664
rect 13446 22652 13452 22664
rect 13504 22692 13510 22704
rect 13504 22664 13584 22692
rect 13504 22652 13510 22664
rect 12158 22624 12164 22636
rect 11808 22596 12164 22624
rect 12158 22584 12164 22596
rect 12216 22624 12222 22636
rect 13556 22633 13584 22664
rect 13648 22633 13676 22732
rect 15105 22729 15117 22763
rect 15151 22729 15163 22763
rect 15105 22723 15163 22729
rect 15197 22763 15255 22769
rect 15197 22729 15209 22763
rect 15243 22760 15255 22763
rect 15562 22760 15568 22772
rect 15243 22732 15568 22760
rect 15243 22729 15255 22732
rect 15197 22723 15255 22729
rect 15120 22692 15148 22723
rect 15562 22720 15568 22732
rect 15620 22720 15626 22772
rect 15841 22763 15899 22769
rect 15841 22729 15853 22763
rect 15887 22760 15899 22763
rect 16022 22760 16028 22772
rect 15887 22732 16028 22760
rect 15887 22729 15899 22732
rect 15841 22723 15899 22729
rect 16022 22720 16028 22732
rect 16080 22720 16086 22772
rect 16485 22763 16543 22769
rect 16485 22729 16497 22763
rect 16531 22729 16543 22763
rect 16485 22723 16543 22729
rect 15378 22692 15384 22704
rect 15120 22664 15384 22692
rect 15378 22652 15384 22664
rect 15436 22652 15442 22704
rect 16500 22692 16528 22723
rect 20438 22720 20444 22772
rect 20496 22760 20502 22772
rect 21085 22763 21143 22769
rect 21085 22760 21097 22763
rect 20496 22732 21097 22760
rect 20496 22720 20502 22732
rect 21085 22729 21097 22732
rect 21131 22760 21143 22763
rect 21131 22732 22232 22760
rect 21131 22729 21143 22732
rect 21085 22723 21143 22729
rect 17006 22695 17064 22701
rect 17006 22692 17018 22695
rect 16500 22664 17018 22692
rect 17006 22661 17018 22664
rect 17052 22661 17064 22695
rect 18322 22692 18328 22704
rect 17006 22655 17064 22661
rect 18248 22664 18328 22692
rect 13998 22633 14004 22636
rect 13265 22627 13323 22633
rect 13265 22624 13277 22627
rect 12216 22596 13277 22624
rect 12216 22584 12222 22596
rect 13265 22593 13277 22596
rect 13311 22593 13323 22627
rect 13265 22587 13323 22593
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22593 13599 22627
rect 13541 22587 13599 22593
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 13992 22587 14004 22633
rect 10965 22559 11023 22565
rect 10965 22525 10977 22559
rect 11011 22556 11023 22559
rect 11716 22556 11744 22584
rect 11011 22528 11744 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 12986 22516 12992 22568
rect 13044 22556 13050 22568
rect 13372 22556 13400 22587
rect 13998 22584 14004 22587
rect 14056 22584 14062 22636
rect 15470 22584 15476 22636
rect 15528 22584 15534 22636
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22624 15991 22627
rect 16206 22624 16212 22636
rect 15979 22596 16212 22624
rect 15979 22593 15991 22596
rect 15933 22587 15991 22593
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22624 16359 22627
rect 16666 22624 16672 22636
rect 16347 22596 16672 22624
rect 16347 22593 16359 22596
rect 16301 22587 16359 22593
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 18248 22633 18276 22664
rect 18322 22652 18328 22664
rect 18380 22692 18386 22704
rect 22002 22692 22008 22704
rect 18380 22664 21312 22692
rect 18380 22652 18386 22664
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22593 18291 22627
rect 18233 22587 18291 22593
rect 18500 22627 18558 22633
rect 18500 22593 18512 22627
rect 18546 22624 18558 22627
rect 19242 22624 19248 22636
rect 18546 22596 19248 22624
rect 18546 22593 18558 22596
rect 18500 22587 18558 22593
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 19720 22633 19748 22664
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22593 19763 22627
rect 19705 22587 19763 22593
rect 19794 22584 19800 22636
rect 19852 22624 19858 22636
rect 19961 22627 20019 22633
rect 19961 22624 19973 22627
rect 19852 22596 19973 22624
rect 19852 22584 19858 22596
rect 19961 22593 19973 22596
rect 20007 22593 20019 22627
rect 19961 22587 20019 22593
rect 13044 22528 13400 22556
rect 13044 22516 13050 22528
rect 13722 22516 13728 22568
rect 13780 22516 13786 22568
rect 15488 22556 15516 22584
rect 21284 22568 21312 22664
rect 21468 22664 22008 22692
rect 21468 22633 21496 22664
rect 22002 22652 22008 22664
rect 22060 22652 22066 22704
rect 21361 22627 21419 22633
rect 21361 22593 21373 22627
rect 21407 22593 21419 22627
rect 21361 22587 21419 22593
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 22204 22624 22232 22732
rect 22278 22720 22284 22772
rect 22336 22720 22342 22772
rect 22462 22720 22468 22772
rect 22520 22720 22526 22772
rect 22554 22720 22560 22772
rect 22612 22760 22618 22772
rect 23293 22763 23351 22769
rect 23293 22760 23305 22763
rect 22612 22732 23305 22760
rect 22612 22720 22618 22732
rect 23293 22729 23305 22732
rect 23339 22729 23351 22763
rect 23293 22723 23351 22729
rect 23566 22720 23572 22772
rect 23624 22720 23630 22772
rect 23658 22720 23664 22772
rect 23716 22720 23722 22772
rect 24210 22760 24216 22772
rect 23860 22732 24216 22760
rect 22296 22692 22324 22720
rect 22480 22692 22508 22720
rect 23860 22701 23888 22732
rect 24210 22720 24216 22732
rect 24268 22720 24274 22772
rect 24305 22763 24363 22769
rect 24305 22729 24317 22763
rect 24351 22760 24363 22763
rect 24351 22732 24440 22760
rect 24351 22729 24363 22732
rect 24305 22723 24363 22729
rect 24412 22704 24440 22732
rect 24486 22720 24492 22772
rect 24544 22760 24550 22772
rect 25774 22760 25780 22772
rect 24544 22732 25780 22760
rect 24544 22720 24550 22732
rect 25774 22720 25780 22732
rect 25832 22760 25838 22772
rect 25961 22763 26019 22769
rect 25961 22760 25973 22763
rect 25832 22732 25973 22760
rect 25832 22720 25838 22732
rect 25961 22729 25973 22732
rect 26007 22729 26019 22763
rect 25961 22723 26019 22729
rect 23043 22695 23101 22701
rect 23043 22692 23055 22695
rect 22296 22664 22416 22692
rect 22480 22664 23055 22692
rect 22278 22624 22284 22636
rect 22204 22596 22284 22624
rect 21453 22587 21511 22593
rect 16574 22556 16580 22568
rect 15488 22528 16580 22556
rect 16574 22516 16580 22528
rect 16632 22516 16638 22568
rect 16758 22516 16764 22568
rect 16816 22516 16822 22568
rect 21266 22516 21272 22568
rect 21324 22516 21330 22568
rect 21376 22556 21404 22587
rect 22278 22584 22284 22596
rect 22336 22584 22342 22636
rect 22388 22630 22416 22664
rect 23043 22661 23055 22664
rect 23089 22661 23101 22695
rect 23043 22655 23101 22661
rect 23845 22695 23903 22701
rect 23845 22661 23857 22695
rect 23891 22661 23903 22695
rect 23845 22655 23903 22661
rect 24026 22652 24032 22704
rect 24084 22692 24090 22704
rect 24084 22664 24348 22692
rect 24084 22652 24090 22664
rect 22465 22630 22523 22633
rect 22388 22627 22523 22630
rect 22388 22602 22477 22627
rect 22465 22593 22477 22602
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 22741 22627 22799 22633
rect 22741 22593 22753 22627
rect 22787 22593 22799 22627
rect 22741 22587 22799 22593
rect 22557 22559 22615 22565
rect 22557 22556 22569 22559
rect 21376 22528 22569 22556
rect 22557 22525 22569 22528
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 22646 22516 22652 22568
rect 22704 22556 22710 22568
rect 22756 22556 22784 22587
rect 22830 22584 22836 22636
rect 22888 22584 22894 22636
rect 22925 22627 22983 22633
rect 22925 22593 22937 22627
rect 22971 22593 22983 22627
rect 23477 22627 23535 22633
rect 23477 22624 23489 22627
rect 22925 22587 22983 22593
rect 23012 22596 23489 22624
rect 22940 22556 22968 22587
rect 22704 22528 22784 22556
rect 22848 22528 22968 22556
rect 22704 22516 22710 22528
rect 10042 22380 10048 22432
rect 10100 22380 10106 22432
rect 10597 22423 10655 22429
rect 10597 22389 10609 22423
rect 10643 22420 10655 22423
rect 12526 22420 12532 22432
rect 10643 22392 12532 22420
rect 10643 22389 10655 22392
rect 10597 22383 10655 22389
rect 12526 22380 12532 22392
rect 12584 22380 12590 22432
rect 13004 22429 13032 22516
rect 15565 22491 15623 22497
rect 15565 22457 15577 22491
rect 15611 22488 15623 22491
rect 18230 22488 18236 22500
rect 15611 22460 16804 22488
rect 15611 22457 15623 22460
rect 15565 22451 15623 22457
rect 12989 22423 13047 22429
rect 12989 22389 13001 22423
rect 13035 22389 13047 22423
rect 12989 22383 13047 22389
rect 15657 22423 15715 22429
rect 15657 22389 15669 22423
rect 15703 22420 15715 22423
rect 16114 22420 16120 22432
rect 15703 22392 16120 22420
rect 15703 22389 15715 22392
rect 15657 22383 15715 22389
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 16776 22420 16804 22460
rect 17972 22460 18236 22488
rect 17972 22420 18000 22460
rect 18230 22448 18236 22460
rect 18288 22448 18294 22500
rect 20806 22448 20812 22500
rect 20864 22448 20870 22500
rect 20990 22448 20996 22500
rect 21048 22488 21054 22500
rect 21048 22460 21312 22488
rect 21048 22448 21054 22460
rect 16776 22392 18000 22420
rect 18046 22380 18052 22432
rect 18104 22420 18110 22432
rect 18141 22423 18199 22429
rect 18141 22420 18153 22423
rect 18104 22392 18153 22420
rect 18104 22380 18110 22392
rect 18141 22389 18153 22392
rect 18187 22389 18199 22423
rect 18141 22383 18199 22389
rect 19613 22423 19671 22429
rect 19613 22389 19625 22423
rect 19659 22420 19671 22423
rect 20824 22420 20852 22448
rect 19659 22392 20852 22420
rect 19659 22389 19671 22392
rect 19613 22383 19671 22389
rect 21174 22380 21180 22432
rect 21232 22380 21238 22432
rect 21284 22420 21312 22460
rect 21450 22448 21456 22500
rect 21508 22488 21514 22500
rect 22848 22488 22876 22528
rect 21508 22460 22876 22488
rect 21508 22448 21514 22460
rect 21821 22423 21879 22429
rect 21821 22420 21833 22423
rect 21284 22392 21833 22420
rect 21821 22389 21833 22392
rect 21867 22389 21879 22423
rect 21821 22383 21879 22389
rect 22186 22380 22192 22432
rect 22244 22420 22250 22432
rect 23012 22420 23040 22596
rect 23477 22593 23489 22596
rect 23523 22624 23535 22627
rect 23750 22624 23756 22636
rect 23523 22596 23756 22624
rect 23523 22593 23535 22596
rect 23477 22587 23535 22593
rect 23750 22584 23756 22596
rect 23808 22584 23814 22636
rect 24121 22627 24179 22633
rect 24121 22593 24133 22627
rect 24167 22593 24179 22627
rect 24121 22587 24179 22593
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 23106 22516 23112 22568
rect 23164 22556 23170 22568
rect 23201 22559 23259 22565
rect 23201 22556 23213 22559
rect 23164 22528 23213 22556
rect 23164 22516 23170 22528
rect 23201 22525 23213 22528
rect 23247 22525 23259 22559
rect 23201 22519 23259 22525
rect 23216 22488 23244 22519
rect 23290 22516 23296 22568
rect 23348 22556 23354 22568
rect 24136 22556 24164 22587
rect 23348 22528 24164 22556
rect 23348 22516 23354 22528
rect 24228 22488 24256 22587
rect 24320 22556 24348 22664
rect 24394 22652 24400 22704
rect 24452 22652 24458 22704
rect 24946 22692 24952 22704
rect 24668 22664 24952 22692
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22624 24547 22627
rect 24668 22624 24696 22664
rect 24946 22652 24952 22664
rect 25004 22652 25010 22704
rect 24854 22633 24860 22636
rect 24535 22596 24696 22624
rect 24837 22627 24860 22633
rect 24535 22593 24547 22596
rect 24489 22587 24547 22593
rect 24837 22593 24849 22627
rect 24837 22587 24860 22593
rect 24854 22584 24860 22587
rect 24912 22584 24918 22636
rect 24581 22559 24639 22565
rect 24581 22556 24593 22559
rect 24320 22528 24593 22556
rect 24581 22525 24593 22528
rect 24627 22525 24639 22559
rect 24581 22519 24639 22525
rect 24486 22488 24492 22500
rect 23216 22460 24492 22488
rect 24486 22448 24492 22460
rect 24544 22448 24550 22500
rect 22244 22392 23040 22420
rect 23937 22423 23995 22429
rect 22244 22380 22250 22392
rect 23937 22389 23949 22423
rect 23983 22420 23995 22423
rect 24762 22420 24768 22432
rect 23983 22392 24768 22420
rect 23983 22389 23995 22392
rect 23937 22383 23995 22389
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 1104 22330 26496 22352
rect 1104 22278 4124 22330
rect 4176 22278 4188 22330
rect 4240 22278 4252 22330
rect 4304 22278 4316 22330
rect 4368 22278 4380 22330
rect 4432 22278 10472 22330
rect 10524 22278 10536 22330
rect 10588 22278 10600 22330
rect 10652 22278 10664 22330
rect 10716 22278 10728 22330
rect 10780 22278 16820 22330
rect 16872 22278 16884 22330
rect 16936 22278 16948 22330
rect 17000 22278 17012 22330
rect 17064 22278 17076 22330
rect 17128 22278 23168 22330
rect 23220 22278 23232 22330
rect 23284 22278 23296 22330
rect 23348 22278 23360 22330
rect 23412 22278 23424 22330
rect 23476 22278 26496 22330
rect 1104 22256 26496 22278
rect 9306 22176 9312 22228
rect 9364 22176 9370 22228
rect 13538 22176 13544 22228
rect 13596 22216 13602 22228
rect 13725 22219 13783 22225
rect 13725 22216 13737 22219
rect 13596 22188 13737 22216
rect 13596 22176 13602 22188
rect 13725 22185 13737 22188
rect 13771 22185 13783 22219
rect 13725 22179 13783 22185
rect 13998 22176 14004 22228
rect 14056 22216 14062 22228
rect 14093 22219 14151 22225
rect 14093 22216 14105 22219
rect 14056 22188 14105 22216
rect 14056 22176 14062 22188
rect 14093 22185 14105 22188
rect 14139 22185 14151 22219
rect 14093 22179 14151 22185
rect 16114 22176 16120 22228
rect 16172 22176 16178 22228
rect 16209 22219 16267 22225
rect 16209 22185 16221 22219
rect 16255 22185 16267 22219
rect 16209 22179 16267 22185
rect 16393 22219 16451 22225
rect 16393 22185 16405 22219
rect 16439 22216 16451 22219
rect 16482 22216 16488 22228
rect 16439 22188 16488 22216
rect 16439 22185 16451 22188
rect 16393 22179 16451 22185
rect 16224 22092 16252 22179
rect 16482 22176 16488 22188
rect 16540 22176 16546 22228
rect 18138 22176 18144 22228
rect 18196 22176 18202 22228
rect 19794 22176 19800 22228
rect 19852 22176 19858 22228
rect 19886 22176 19892 22228
rect 19944 22176 19950 22228
rect 22738 22216 22744 22228
rect 22296 22188 22744 22216
rect 18156 22148 18184 22176
rect 17972 22120 18184 22148
rect 18233 22151 18291 22157
rect 12989 22083 13047 22089
rect 12989 22049 13001 22083
rect 13035 22080 13047 22083
rect 13722 22080 13728 22092
rect 13035 22052 13728 22080
rect 13035 22049 13047 22052
rect 12989 22043 13047 22049
rect 13722 22040 13728 22052
rect 13780 22080 13786 22092
rect 14734 22080 14740 22092
rect 13780 22052 14740 22080
rect 13780 22040 13786 22052
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 16206 22040 16212 22092
rect 16264 22040 16270 22092
rect 9401 22015 9459 22021
rect 9401 21981 9413 22015
rect 9447 22012 9459 22015
rect 10042 22012 10048 22024
rect 9447 21984 10048 22012
rect 9447 21981 9459 21984
rect 9401 21975 9459 21981
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 13081 22015 13139 22021
rect 13081 21981 13093 22015
rect 13127 21981 13139 22015
rect 13081 21975 13139 21981
rect 12342 21904 12348 21956
rect 12400 21944 12406 21956
rect 12722 21947 12780 21953
rect 12722 21944 12734 21947
rect 12400 21916 12734 21944
rect 12400 21904 12406 21916
rect 12722 21913 12734 21916
rect 12768 21913 12780 21947
rect 12722 21907 12780 21913
rect 11609 21879 11667 21885
rect 11609 21845 11621 21879
rect 11655 21876 11667 21879
rect 11698 21876 11704 21888
rect 11655 21848 11704 21876
rect 11655 21845 11667 21848
rect 11609 21839 11667 21845
rect 11698 21836 11704 21848
rect 11756 21876 11762 21888
rect 13096 21876 13124 21975
rect 13630 21972 13636 22024
rect 13688 21972 13694 22024
rect 14274 21972 14280 22024
rect 14332 21972 14338 22024
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 13648 21944 13676 21972
rect 14476 21944 14504 21975
rect 14550 21972 14556 22024
rect 14608 21972 14614 22024
rect 14752 22012 14780 22040
rect 16666 22012 16672 22024
rect 14752 21984 16672 22012
rect 16666 21972 16672 21984
rect 16724 22012 16730 22024
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16724 21984 16865 22012
rect 16724 21972 16730 21984
rect 16853 21981 16865 21984
rect 16899 21981 16911 22015
rect 16853 21975 16911 21981
rect 13648 21916 14504 21944
rect 14642 21904 14648 21956
rect 14700 21944 14706 21956
rect 14982 21947 15040 21953
rect 14982 21944 14994 21947
rect 14700 21916 14994 21944
rect 14700 21904 14706 21916
rect 14982 21913 14994 21916
rect 15028 21913 15040 21947
rect 14982 21907 15040 21913
rect 15378 21904 15384 21956
rect 15436 21904 15442 21956
rect 16390 21953 16396 21956
rect 16377 21947 16396 21953
rect 16377 21913 16389 21947
rect 16377 21907 16396 21913
rect 16390 21904 16396 21907
rect 16448 21904 16454 21956
rect 16577 21947 16635 21953
rect 16577 21913 16589 21947
rect 16623 21913 16635 21947
rect 16577 21907 16635 21913
rect 17120 21947 17178 21953
rect 17120 21913 17132 21947
rect 17166 21944 17178 21947
rect 17972 21944 18000 22120
rect 18233 22117 18245 22151
rect 18279 22148 18291 22151
rect 22296 22148 22324 22188
rect 22738 22176 22744 22188
rect 22796 22176 22802 22228
rect 22922 22176 22928 22228
rect 22980 22176 22986 22228
rect 24397 22219 24455 22225
rect 24397 22185 24409 22219
rect 24443 22216 24455 22219
rect 24854 22216 24860 22228
rect 24443 22188 24860 22216
rect 24443 22185 24455 22188
rect 24397 22179 24455 22185
rect 24854 22176 24860 22188
rect 24912 22176 24918 22228
rect 18279 22120 18368 22148
rect 18279 22117 18291 22120
rect 18233 22111 18291 22117
rect 18138 22040 18144 22092
rect 18196 22080 18202 22092
rect 18340 22089 18368 22120
rect 22204 22120 22324 22148
rect 22649 22151 22707 22157
rect 18325 22083 18383 22089
rect 18325 22080 18337 22083
rect 18196 22052 18337 22080
rect 18196 22040 18202 22052
rect 18325 22049 18337 22052
rect 18371 22049 18383 22083
rect 18325 22043 18383 22049
rect 21266 22040 21272 22092
rect 21324 22080 21330 22092
rect 22097 22083 22155 22089
rect 22097 22080 22109 22083
rect 21324 22052 22109 22080
rect 21324 22040 21330 22052
rect 22097 22049 22109 22052
rect 22143 22080 22155 22083
rect 22204 22080 22232 22120
rect 22649 22117 22661 22151
rect 22695 22148 22707 22151
rect 22940 22148 22968 22176
rect 22695 22120 22968 22148
rect 22695 22117 22707 22120
rect 22649 22111 22707 22117
rect 22925 22083 22983 22089
rect 22925 22080 22937 22083
rect 22143 22052 22232 22080
rect 22480 22052 22937 22080
rect 22143 22049 22155 22052
rect 22097 22043 22155 22049
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 17166 21916 17356 21944
rect 17166 21913 17178 21916
rect 17120 21907 17178 21913
rect 11756 21848 13124 21876
rect 15396 21876 15424 21904
rect 16592 21876 16620 21907
rect 17328 21888 17356 21916
rect 17788 21916 18000 21944
rect 19628 21944 19656 21975
rect 20990 21972 20996 22024
rect 21048 22021 21054 22024
rect 21048 21975 21060 22021
rect 21048 21972 21054 21975
rect 21634 21972 21640 22024
rect 21692 22012 21698 22024
rect 22480 22012 22508 22052
rect 22925 22049 22937 22052
rect 22971 22049 22983 22083
rect 22925 22043 22983 22049
rect 23017 22083 23075 22089
rect 23017 22049 23029 22083
rect 23063 22080 23075 22083
rect 24118 22080 24124 22092
rect 23063 22052 24124 22080
rect 23063 22049 23075 22052
rect 23017 22043 23075 22049
rect 24118 22040 24124 22052
rect 24176 22040 24182 22092
rect 25130 22080 25136 22092
rect 24228 22052 25136 22080
rect 21692 21984 22508 22012
rect 22833 22015 22891 22021
rect 21692 21972 21698 21984
rect 22833 21981 22845 22015
rect 22879 21981 22891 22015
rect 23845 22015 23903 22021
rect 23845 22012 23857 22015
rect 22833 21975 22891 21981
rect 23768 21984 23857 22012
rect 21174 21944 21180 21956
rect 19628 21916 21180 21944
rect 17788 21888 17816 21916
rect 21174 21904 21180 21916
rect 21232 21904 21238 21956
rect 21358 21904 21364 21956
rect 21416 21904 21422 21956
rect 22848 21944 22876 21975
rect 23658 21944 23664 21956
rect 22848 21916 23664 21944
rect 23658 21904 23664 21916
rect 23716 21904 23722 21956
rect 15396 21848 16620 21876
rect 11756 21836 11762 21848
rect 17310 21836 17316 21888
rect 17368 21836 17374 21888
rect 17770 21836 17776 21888
rect 17828 21836 17834 21888
rect 18966 21836 18972 21888
rect 19024 21836 19030 21888
rect 22922 21836 22928 21888
rect 22980 21876 22986 21888
rect 23768 21876 23796 21984
rect 23845 21981 23857 21984
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 24026 21972 24032 22024
rect 24084 22012 24090 22024
rect 24228 22012 24256 22052
rect 25130 22040 25136 22052
rect 25188 22040 25194 22092
rect 25774 22040 25780 22092
rect 25832 22040 25838 22092
rect 24084 21984 24256 22012
rect 24581 22015 24639 22021
rect 24084 21972 24090 21984
rect 24581 21981 24593 22015
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 23937 21947 23995 21953
rect 23937 21913 23949 21947
rect 23983 21944 23995 21947
rect 24596 21944 24624 21975
rect 24762 21972 24768 22024
rect 24820 21972 24826 22024
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 22012 24915 22015
rect 25225 22015 25283 22021
rect 25225 22012 25237 22015
rect 24903 21984 25237 22012
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 25225 21981 25237 21984
rect 25271 21981 25283 22015
rect 25225 21975 25283 21981
rect 23983 21916 24624 21944
rect 23983 21913 23995 21916
rect 23937 21907 23995 21913
rect 22980 21848 23796 21876
rect 22980 21836 22986 21848
rect 1104 21786 26656 21808
rect 1104 21734 7298 21786
rect 7350 21734 7362 21786
rect 7414 21734 7426 21786
rect 7478 21734 7490 21786
rect 7542 21734 7554 21786
rect 7606 21734 13646 21786
rect 13698 21734 13710 21786
rect 13762 21734 13774 21786
rect 13826 21734 13838 21786
rect 13890 21734 13902 21786
rect 13954 21734 19994 21786
rect 20046 21734 20058 21786
rect 20110 21734 20122 21786
rect 20174 21734 20186 21786
rect 20238 21734 20250 21786
rect 20302 21734 26342 21786
rect 26394 21734 26406 21786
rect 26458 21734 26470 21786
rect 26522 21734 26534 21786
rect 26586 21734 26598 21786
rect 26650 21734 26656 21786
rect 1104 21712 26656 21734
rect 8110 21632 8116 21684
rect 8168 21632 8174 21684
rect 12253 21675 12311 21681
rect 12253 21641 12265 21675
rect 12299 21672 12311 21675
rect 12342 21672 12348 21684
rect 12299 21644 12348 21672
rect 12299 21641 12311 21644
rect 12253 21635 12311 21641
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 14734 21632 14740 21684
rect 14792 21632 14798 21684
rect 15378 21632 15384 21684
rect 15436 21632 15442 21684
rect 15841 21675 15899 21681
rect 15841 21641 15853 21675
rect 15887 21672 15899 21675
rect 15930 21672 15936 21684
rect 15887 21644 15936 21672
rect 15887 21641 15899 21644
rect 15841 21635 15899 21641
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 16022 21632 16028 21684
rect 16080 21632 16086 21684
rect 17310 21632 17316 21684
rect 17368 21632 17374 21684
rect 17402 21632 17408 21684
rect 17460 21672 17466 21684
rect 17589 21675 17647 21681
rect 17589 21672 17601 21675
rect 17460 21644 17601 21672
rect 17460 21632 17466 21644
rect 17589 21641 17601 21644
rect 17635 21641 17647 21675
rect 17589 21635 17647 21641
rect 8128 21604 8156 21632
rect 14752 21604 14780 21632
rect 7668 21576 8156 21604
rect 14476 21576 14780 21604
rect 7668 21545 7696 21576
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 12158 21496 12164 21548
rect 12216 21496 12222 21548
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21536 12403 21539
rect 13078 21536 13084 21548
rect 12391 21508 13084 21536
rect 12391 21505 12403 21508
rect 12345 21499 12403 21505
rect 13078 21496 13084 21508
rect 13136 21496 13142 21548
rect 14476 21545 14504 21576
rect 15010 21564 15016 21616
rect 15068 21564 15074 21616
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21505 14519 21539
rect 14461 21499 14519 21505
rect 14728 21539 14786 21545
rect 14728 21505 14740 21539
rect 14774 21536 14786 21539
rect 15028 21536 15056 21564
rect 14774 21508 15056 21536
rect 15396 21536 15424 21632
rect 16574 21564 16580 21616
rect 16632 21604 16638 21616
rect 17037 21607 17095 21613
rect 17037 21604 17049 21607
rect 16632 21576 17049 21604
rect 16632 21564 16638 21576
rect 17037 21573 17049 21576
rect 17083 21604 17095 21607
rect 17604 21604 17632 21635
rect 17678 21632 17684 21684
rect 17736 21632 17742 21684
rect 17773 21675 17831 21681
rect 17773 21641 17785 21675
rect 17819 21672 17831 21675
rect 18046 21672 18052 21684
rect 17819 21644 18052 21672
rect 17819 21641 17831 21644
rect 17773 21635 17831 21641
rect 17972 21604 18000 21644
rect 18046 21632 18052 21644
rect 18104 21632 18110 21684
rect 18141 21675 18199 21681
rect 18141 21641 18153 21675
rect 18187 21672 18199 21675
rect 18230 21672 18236 21684
rect 18187 21644 18236 21672
rect 18187 21641 18199 21644
rect 18141 21635 18199 21641
rect 18230 21632 18236 21644
rect 18288 21632 18294 21684
rect 18966 21672 18972 21684
rect 18616 21644 18972 21672
rect 18616 21613 18644 21644
rect 18966 21632 18972 21644
rect 19024 21632 19030 21684
rect 21453 21675 21511 21681
rect 21453 21641 21465 21675
rect 21499 21672 21511 21675
rect 21910 21672 21916 21684
rect 21499 21644 21916 21672
rect 21499 21641 21511 21644
rect 21453 21635 21511 21641
rect 21910 21632 21916 21644
rect 21968 21632 21974 21684
rect 22646 21672 22652 21684
rect 22066 21644 22652 21672
rect 18417 21607 18475 21613
rect 18417 21604 18429 21607
rect 17083 21576 17540 21604
rect 17604 21576 17825 21604
rect 17972 21576 18429 21604
rect 17083 21573 17095 21576
rect 17037 21567 17095 21573
rect 16117 21539 16175 21545
rect 16117 21536 16129 21539
rect 15396 21508 16129 21536
rect 14774 21505 14786 21508
rect 14728 21499 14786 21505
rect 16117 21505 16129 21508
rect 16163 21505 16175 21539
rect 16117 21499 16175 21505
rect 16206 21496 16212 21548
rect 16264 21536 16270 21548
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 16264 21508 16681 21536
rect 16264 21496 16270 21508
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 16758 21496 16764 21548
rect 16816 21496 16822 21548
rect 17313 21539 17371 21545
rect 17313 21505 17325 21539
rect 17359 21536 17371 21539
rect 17402 21536 17408 21548
rect 17359 21508 17408 21536
rect 17359 21505 17371 21508
rect 17313 21499 17371 21505
rect 17402 21496 17408 21508
rect 17460 21496 17466 21548
rect 17512 21536 17540 21576
rect 17586 21536 17592 21548
rect 17512 21508 17592 21536
rect 17586 21496 17592 21508
rect 17644 21496 17650 21548
rect 17797 21536 17825 21576
rect 18417 21573 18429 21576
rect 18463 21573 18475 21607
rect 18417 21567 18475 21573
rect 18601 21607 18659 21613
rect 18601 21573 18613 21607
rect 18647 21573 18659 21607
rect 18601 21567 18659 21573
rect 19886 21564 19892 21616
rect 19944 21564 19950 21616
rect 22066 21604 22094 21644
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 23658 21632 23664 21684
rect 23716 21672 23722 21684
rect 24762 21672 24768 21684
rect 23716 21644 24768 21672
rect 23716 21632 23722 21644
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 25314 21632 25320 21684
rect 25372 21672 25378 21684
rect 25501 21675 25559 21681
rect 25501 21672 25513 21675
rect 25372 21644 25513 21672
rect 25372 21632 25378 21644
rect 25501 21641 25513 21644
rect 25547 21641 25559 21675
rect 25501 21635 25559 21641
rect 23017 21607 23075 21613
rect 23017 21604 23029 21607
rect 21560 21576 22094 21604
rect 22480 21576 23029 21604
rect 17862 21536 17868 21548
rect 17797 21508 17868 21536
rect 17862 21496 17868 21508
rect 17920 21496 17926 21548
rect 18046 21496 18052 21548
rect 18104 21496 18110 21548
rect 18230 21496 18236 21548
rect 18288 21496 18294 21548
rect 18322 21496 18328 21548
rect 18380 21496 18386 21548
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20622 21536 20628 21548
rect 20303 21508 20628 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 20806 21496 20812 21548
rect 20864 21536 20870 21548
rect 21361 21539 21419 21545
rect 21361 21536 21373 21539
rect 20864 21508 21373 21536
rect 20864 21496 20870 21508
rect 21361 21505 21373 21508
rect 21407 21536 21419 21539
rect 21450 21536 21456 21548
rect 21407 21508 21456 21536
rect 21407 21505 21419 21508
rect 21361 21499 21419 21505
rect 21450 21496 21456 21508
rect 21508 21496 21514 21548
rect 21560 21545 21588 21576
rect 21545 21539 21603 21545
rect 21545 21505 21557 21539
rect 21591 21505 21603 21539
rect 21545 21499 21603 21505
rect 22002 21496 22008 21548
rect 22060 21496 22066 21548
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22480 21545 22508 21576
rect 23017 21573 23029 21576
rect 23063 21573 23075 21607
rect 24780 21604 24808 21632
rect 24780 21576 25728 21604
rect 23017 21567 23075 21573
rect 22281 21539 22339 21545
rect 22281 21536 22293 21539
rect 22152 21508 22293 21536
rect 22152 21496 22158 21508
rect 22281 21505 22293 21508
rect 22327 21505 22339 21539
rect 22281 21499 22339 21505
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21536 22707 21539
rect 22833 21539 22891 21545
rect 22695 21508 22784 21536
rect 22695 21505 22707 21508
rect 22649 21499 22707 21505
rect 7926 21428 7932 21480
rect 7984 21428 7990 21480
rect 22296 21468 22324 21499
rect 22572 21468 22600 21499
rect 22296 21440 22600 21468
rect 22756 21468 22784 21508
rect 22833 21505 22845 21539
rect 22879 21536 22891 21539
rect 23658 21536 23664 21548
rect 22879 21508 23664 21536
rect 22879 21505 22891 21508
rect 22833 21499 22891 21505
rect 23658 21496 23664 21508
rect 23716 21496 23722 21548
rect 23934 21496 23940 21548
rect 23992 21496 23998 21548
rect 24118 21496 24124 21548
rect 24176 21536 24182 21548
rect 25700 21545 25728 21576
rect 24213 21539 24271 21545
rect 24213 21536 24225 21539
rect 24176 21508 24225 21536
rect 24176 21496 24182 21508
rect 24213 21505 24225 21508
rect 24259 21505 24271 21539
rect 24213 21499 24271 21505
rect 24397 21539 24455 21545
rect 24397 21505 24409 21539
rect 24443 21536 24455 21539
rect 24765 21539 24823 21545
rect 24765 21536 24777 21539
rect 24443 21508 24777 21536
rect 24443 21505 24455 21508
rect 24397 21499 24455 21505
rect 24765 21505 24777 21508
rect 24811 21505 24823 21539
rect 24765 21499 24823 21505
rect 25685 21539 25743 21545
rect 25685 21505 25697 21539
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 25774 21496 25780 21548
rect 25832 21496 25838 21548
rect 23566 21468 23572 21480
rect 22756 21440 23572 21468
rect 22572 21412 22600 21440
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 25314 21428 25320 21480
rect 25372 21428 25378 21480
rect 17218 21360 17224 21412
rect 17276 21360 17282 21412
rect 17957 21403 18015 21409
rect 17957 21369 17969 21403
rect 18003 21400 18015 21403
rect 18046 21400 18052 21412
rect 18003 21372 18052 21400
rect 18003 21369 18015 21372
rect 17957 21363 18015 21369
rect 18046 21360 18052 21372
rect 18104 21360 18110 21412
rect 18598 21360 18604 21412
rect 18656 21360 18662 21412
rect 22554 21360 22560 21412
rect 22612 21400 22618 21412
rect 24026 21400 24032 21412
rect 22612 21372 24032 21400
rect 22612 21360 22618 21372
rect 24026 21360 24032 21372
rect 24084 21360 24090 21412
rect 9401 21335 9459 21341
rect 9401 21301 9413 21335
rect 9447 21332 9459 21335
rect 9582 21332 9588 21344
rect 9447 21304 9588 21332
rect 9447 21301 9459 21304
rect 9401 21295 9459 21301
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 17405 21335 17463 21341
rect 17405 21301 17417 21335
rect 17451 21332 17463 21335
rect 17494 21332 17500 21344
rect 17451 21304 17500 21332
rect 17451 21301 17463 21304
rect 17405 21295 17463 21301
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 21821 21335 21879 21341
rect 21821 21301 21833 21335
rect 21867 21332 21879 21335
rect 22094 21332 22100 21344
rect 21867 21304 22100 21332
rect 21867 21301 21879 21304
rect 21821 21295 21879 21301
rect 22094 21292 22100 21304
rect 22152 21292 22158 21344
rect 22830 21292 22836 21344
rect 22888 21292 22894 21344
rect 23753 21335 23811 21341
rect 23753 21301 23765 21335
rect 23799 21332 23811 21335
rect 24210 21332 24216 21344
rect 23799 21304 24216 21332
rect 23799 21301 23811 21304
rect 23753 21295 23811 21301
rect 24210 21292 24216 21304
rect 24268 21292 24274 21344
rect 1104 21242 26496 21264
rect 1104 21190 4124 21242
rect 4176 21190 4188 21242
rect 4240 21190 4252 21242
rect 4304 21190 4316 21242
rect 4368 21190 4380 21242
rect 4432 21190 10472 21242
rect 10524 21190 10536 21242
rect 10588 21190 10600 21242
rect 10652 21190 10664 21242
rect 10716 21190 10728 21242
rect 10780 21190 16820 21242
rect 16872 21190 16884 21242
rect 16936 21190 16948 21242
rect 17000 21190 17012 21242
rect 17064 21190 17076 21242
rect 17128 21190 23168 21242
rect 23220 21190 23232 21242
rect 23284 21190 23296 21242
rect 23348 21190 23360 21242
rect 23412 21190 23424 21242
rect 23476 21190 26496 21242
rect 1104 21168 26496 21190
rect 16316 21100 17356 21128
rect 8128 21032 9628 21060
rect 8021 20927 8079 20933
rect 8021 20893 8033 20927
rect 8067 20924 8079 20927
rect 8128 20924 8156 21032
rect 8220 20964 8800 20992
rect 8220 20933 8248 20964
rect 8772 20936 8800 20964
rect 9600 20936 9628 21032
rect 11330 20992 11336 21004
rect 10796 20964 11336 20992
rect 8067 20896 8156 20924
rect 8205 20927 8263 20933
rect 8067 20893 8079 20896
rect 8021 20887 8079 20893
rect 8205 20893 8217 20927
rect 8251 20893 8263 20927
rect 8205 20887 8263 20893
rect 8481 20927 8539 20933
rect 8481 20893 8493 20927
rect 8527 20924 8539 20927
rect 8570 20924 8576 20936
rect 8527 20896 8576 20924
rect 8527 20893 8539 20896
rect 8481 20887 8539 20893
rect 8570 20884 8576 20896
rect 8628 20884 8634 20936
rect 8754 20884 8760 20936
rect 8812 20884 8818 20936
rect 9493 20927 9551 20933
rect 9493 20924 9505 20927
rect 9416 20896 9505 20924
rect 8113 20859 8171 20865
rect 8113 20825 8125 20859
rect 8159 20856 8171 20859
rect 8386 20856 8392 20868
rect 8159 20828 8392 20856
rect 8159 20825 8171 20828
rect 8113 20819 8171 20825
rect 8386 20816 8392 20828
rect 8444 20816 8450 20868
rect 9416 20800 9444 20896
rect 9493 20893 9505 20896
rect 9539 20893 9551 20927
rect 9493 20887 9551 20893
rect 9582 20884 9588 20936
rect 9640 20924 9646 20936
rect 10796 20933 10824 20964
rect 11330 20952 11336 20964
rect 11388 20952 11394 21004
rect 14734 20952 14740 21004
rect 14792 20992 14798 21004
rect 15473 20995 15531 21001
rect 15473 20992 15485 20995
rect 14792 20964 15485 20992
rect 14792 20952 14798 20964
rect 15473 20961 15485 20964
rect 15519 20961 15531 20995
rect 15473 20955 15531 20961
rect 16316 20936 16344 21100
rect 16482 21020 16488 21072
rect 16540 21060 16546 21072
rect 16761 21063 16819 21069
rect 16540 21032 16712 21060
rect 16540 21020 16546 21032
rect 10229 20927 10287 20933
rect 10229 20924 10241 20927
rect 9640 20896 10241 20924
rect 9640 20884 9646 20896
rect 10229 20893 10241 20896
rect 10275 20893 10287 20927
rect 10229 20887 10287 20893
rect 10781 20927 10839 20933
rect 10781 20893 10793 20927
rect 10827 20893 10839 20927
rect 10781 20887 10839 20893
rect 11057 20927 11115 20933
rect 11057 20893 11069 20927
rect 11103 20893 11115 20927
rect 11057 20887 11115 20893
rect 11072 20856 11100 20887
rect 16298 20884 16304 20936
rect 16356 20884 16362 20936
rect 16485 20927 16543 20933
rect 16485 20893 16497 20927
rect 16531 20893 16543 20927
rect 16684 20924 16712 21032
rect 16761 21029 16773 21063
rect 16807 21060 16819 21063
rect 17034 21060 17040 21072
rect 16807 21032 17040 21060
rect 16807 21029 16819 21032
rect 16761 21023 16819 21029
rect 17034 21020 17040 21032
rect 17092 21020 17098 21072
rect 17126 21020 17132 21072
rect 17184 21060 17190 21072
rect 17221 21063 17279 21069
rect 17221 21060 17233 21063
rect 17184 21032 17233 21060
rect 17184 21020 17190 21032
rect 17221 21029 17233 21032
rect 17267 21029 17279 21063
rect 17328 21060 17356 21100
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 18230 21128 18236 21140
rect 17920 21100 18236 21128
rect 17920 21088 17926 21100
rect 18230 21088 18236 21100
rect 18288 21128 18294 21140
rect 18325 21131 18383 21137
rect 18325 21128 18337 21131
rect 18288 21100 18337 21128
rect 18288 21088 18294 21100
rect 18325 21097 18337 21100
rect 18371 21097 18383 21131
rect 18325 21091 18383 21097
rect 22002 21088 22008 21140
rect 22060 21128 22066 21140
rect 22373 21131 22431 21137
rect 22373 21128 22385 21131
rect 22060 21100 22385 21128
rect 22060 21088 22066 21100
rect 22373 21097 22385 21100
rect 22419 21097 22431 21131
rect 22373 21091 22431 21097
rect 23198 21088 23204 21140
rect 23256 21128 23262 21140
rect 25314 21128 25320 21140
rect 23256 21100 25320 21128
rect 23256 21088 23262 21100
rect 25314 21088 25320 21100
rect 25372 21128 25378 21140
rect 25777 21131 25835 21137
rect 25777 21128 25789 21131
rect 25372 21100 25789 21128
rect 25372 21088 25378 21100
rect 25777 21097 25789 21100
rect 25823 21097 25835 21131
rect 25777 21091 25835 21097
rect 17328 21032 19334 21060
rect 17221 21023 17279 21029
rect 16761 20927 16819 20933
rect 16761 20924 16773 20927
rect 16684 20896 16773 20924
rect 16485 20887 16543 20893
rect 16761 20893 16773 20896
rect 16807 20893 16819 20927
rect 16761 20887 16819 20893
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20893 16911 20927
rect 16853 20887 16911 20893
rect 11238 20856 11244 20868
rect 11072 20828 11244 20856
rect 11238 20816 11244 20828
rect 11296 20816 11302 20868
rect 11333 20859 11391 20865
rect 11333 20825 11345 20859
rect 11379 20825 11391 20859
rect 12618 20856 12624 20868
rect 12558 20828 12624 20856
rect 11333 20819 11391 20825
rect 7834 20748 7840 20800
rect 7892 20788 7898 20800
rect 8294 20788 8300 20800
rect 7892 20760 8300 20788
rect 7892 20748 7898 20760
rect 8294 20748 8300 20760
rect 8352 20748 8358 20800
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 8846 20788 8852 20800
rect 8720 20760 8852 20788
rect 8720 20748 8726 20760
rect 8846 20748 8852 20760
rect 8904 20748 8910 20800
rect 8938 20748 8944 20800
rect 8996 20748 9002 20800
rect 9398 20748 9404 20800
rect 9456 20748 9462 20800
rect 9674 20748 9680 20800
rect 9732 20748 9738 20800
rect 10965 20791 11023 20797
rect 10965 20757 10977 20791
rect 11011 20788 11023 20791
rect 11348 20788 11376 20819
rect 12618 20816 12624 20828
rect 12676 20816 12682 20868
rect 16500 20856 16528 20887
rect 16868 20856 16896 20887
rect 17034 20884 17040 20936
rect 17092 20924 17098 20936
rect 17773 20927 17831 20933
rect 17773 20924 17785 20927
rect 17092 20896 17785 20924
rect 17092 20884 17098 20896
rect 17773 20893 17785 20896
rect 17819 20893 17831 20927
rect 17773 20887 17831 20893
rect 18138 20884 18144 20936
rect 18196 20924 18202 20936
rect 18233 20927 18291 20933
rect 18233 20924 18245 20927
rect 18196 20896 18245 20924
rect 18196 20884 18202 20896
rect 18233 20893 18245 20896
rect 18279 20893 18291 20927
rect 18233 20887 18291 20893
rect 18598 20884 18604 20936
rect 18656 20884 18662 20936
rect 19306 20924 19334 21032
rect 24397 20995 24455 21001
rect 24397 20992 24409 20995
rect 22664 20964 23428 20992
rect 21358 20924 21364 20936
rect 19306 20896 21364 20924
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 22554 20884 22560 20936
rect 22612 20884 22618 20936
rect 22664 20933 22692 20964
rect 23400 20936 23428 20964
rect 23492 20964 24409 20992
rect 22649 20927 22707 20933
rect 22649 20893 22661 20927
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 22738 20884 22744 20936
rect 22796 20924 22802 20936
rect 22833 20927 22891 20933
rect 22833 20924 22845 20927
rect 22796 20896 22845 20924
rect 22796 20884 22802 20896
rect 22833 20893 22845 20896
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 22922 20884 22928 20936
rect 22980 20884 22986 20936
rect 23017 20927 23075 20933
rect 23017 20893 23029 20927
rect 23063 20924 23075 20927
rect 23198 20924 23204 20936
rect 23063 20896 23204 20924
rect 23063 20893 23075 20896
rect 23017 20887 23075 20893
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 23382 20884 23388 20936
rect 23440 20884 23446 20936
rect 16500 20828 16896 20856
rect 16684 20800 16712 20828
rect 16942 20816 16948 20868
rect 17000 20816 17006 20868
rect 17129 20859 17187 20865
rect 17129 20825 17141 20859
rect 17175 20825 17187 20859
rect 17129 20819 17187 20825
rect 11011 20760 11376 20788
rect 11011 20757 11023 20760
rect 10965 20751 11023 20757
rect 12802 20748 12808 20800
rect 12860 20748 12866 20800
rect 16574 20748 16580 20800
rect 16632 20748 16638 20800
rect 16666 20748 16672 20800
rect 16724 20748 16730 20800
rect 17034 20797 17040 20800
rect 17030 20751 17040 20797
rect 17034 20748 17040 20751
rect 17092 20748 17098 20800
rect 17147 20788 17175 20819
rect 22186 20816 22192 20868
rect 22244 20856 22250 20868
rect 23492 20856 23520 20964
rect 24397 20961 24409 20964
rect 24443 20961 24455 20995
rect 24397 20955 24455 20961
rect 23566 20884 23572 20936
rect 23624 20924 23630 20936
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 23624 20896 23765 20924
rect 23624 20884 23630 20896
rect 23753 20893 23765 20896
rect 23799 20893 23811 20927
rect 23753 20887 23811 20893
rect 24210 20884 24216 20936
rect 24268 20924 24274 20936
rect 24653 20927 24711 20933
rect 24653 20924 24665 20927
rect 24268 20896 24665 20924
rect 24268 20884 24274 20896
rect 24653 20893 24665 20896
rect 24699 20893 24711 20927
rect 24653 20887 24711 20893
rect 22244 20828 23520 20856
rect 22244 20816 22250 20828
rect 18230 20788 18236 20800
rect 17147 20760 18236 20788
rect 18230 20748 18236 20760
rect 18288 20748 18294 20800
rect 18322 20748 18328 20800
rect 18380 20748 18386 20800
rect 18414 20748 18420 20800
rect 18472 20748 18478 20800
rect 22738 20748 22744 20800
rect 22796 20788 22802 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 22796 20760 23305 20788
rect 22796 20748 22802 20760
rect 23293 20757 23305 20760
rect 23339 20788 23351 20791
rect 23750 20788 23756 20800
rect 23339 20760 23756 20788
rect 23339 20757 23351 20760
rect 23293 20751 23351 20757
rect 23750 20748 23756 20760
rect 23808 20748 23814 20800
rect 1104 20698 26656 20720
rect 1104 20646 7298 20698
rect 7350 20646 7362 20698
rect 7414 20646 7426 20698
rect 7478 20646 7490 20698
rect 7542 20646 7554 20698
rect 7606 20646 13646 20698
rect 13698 20646 13710 20698
rect 13762 20646 13774 20698
rect 13826 20646 13838 20698
rect 13890 20646 13902 20698
rect 13954 20646 19994 20698
rect 20046 20646 20058 20698
rect 20110 20646 20122 20698
rect 20174 20646 20186 20698
rect 20238 20646 20250 20698
rect 20302 20646 26342 20698
rect 26394 20646 26406 20698
rect 26458 20646 26470 20698
rect 26522 20646 26534 20698
rect 26586 20646 26598 20698
rect 26650 20646 26656 20698
rect 1104 20624 26656 20646
rect 8662 20544 8668 20596
rect 8720 20544 8726 20596
rect 11330 20544 11336 20596
rect 11388 20584 11394 20596
rect 11517 20587 11575 20593
rect 11517 20584 11529 20587
rect 11388 20556 11529 20584
rect 11388 20544 11394 20556
rect 11517 20553 11529 20556
rect 11563 20553 11575 20587
rect 11974 20584 11980 20596
rect 11517 20547 11575 20553
rect 11624 20556 11980 20584
rect 8680 20516 8708 20544
rect 11624 20528 11652 20556
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 15102 20584 15108 20596
rect 12545 20556 15108 20584
rect 7392 20488 8708 20516
rect 7392 20457 7420 20488
rect 9030 20476 9036 20528
rect 9088 20476 9094 20528
rect 10689 20519 10747 20525
rect 10689 20485 10701 20519
rect 10735 20516 10747 20519
rect 11238 20516 11244 20528
rect 10735 20488 11244 20516
rect 10735 20485 10747 20488
rect 10689 20479 10747 20485
rect 11238 20476 11244 20488
rect 11296 20476 11302 20528
rect 11606 20476 11612 20528
rect 11664 20476 11670 20528
rect 12545 20516 12573 20556
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 16592 20556 17724 20584
rect 16592 20528 16620 20556
rect 12802 20516 12808 20528
rect 11808 20488 12573 20516
rect 12636 20488 12808 20516
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 7558 20408 7564 20460
rect 7616 20408 7622 20460
rect 7653 20451 7711 20457
rect 7653 20417 7665 20451
rect 7699 20417 7711 20451
rect 7653 20411 7711 20417
rect 7745 20451 7803 20457
rect 7745 20417 7757 20451
rect 7791 20448 7803 20451
rect 7834 20448 7840 20460
rect 7791 20420 7840 20448
rect 7791 20417 7803 20420
rect 7745 20411 7803 20417
rect 7668 20244 7696 20411
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 8018 20408 8024 20460
rect 8076 20408 8082 20460
rect 9858 20408 9864 20460
rect 9916 20448 9922 20460
rect 11808 20448 11836 20488
rect 9916 20420 11836 20448
rect 9916 20408 9922 20420
rect 11882 20408 11888 20460
rect 11940 20408 11946 20460
rect 8297 20383 8355 20389
rect 8297 20380 8309 20383
rect 7944 20352 8309 20380
rect 7944 20321 7972 20352
rect 8297 20349 8309 20352
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 9030 20340 9036 20392
rect 9088 20380 9094 20392
rect 10042 20380 10048 20392
rect 9088 20352 10048 20380
rect 9088 20340 9094 20352
rect 10042 20340 10048 20352
rect 10100 20340 10106 20392
rect 12161 20383 12219 20389
rect 12161 20349 12173 20383
rect 12207 20380 12219 20383
rect 12636 20380 12664 20488
rect 12802 20476 12808 20488
rect 12860 20516 12866 20528
rect 12860 20488 14044 20516
rect 12860 20476 12866 20488
rect 13170 20408 13176 20460
rect 13228 20448 13234 20460
rect 14016 20457 14044 20488
rect 16574 20476 16580 20528
rect 16632 20476 16638 20528
rect 16669 20519 16727 20525
rect 16669 20485 16681 20519
rect 16715 20516 16727 20519
rect 16758 20516 16764 20528
rect 16715 20488 16764 20516
rect 16715 20485 16727 20488
rect 16669 20479 16727 20485
rect 16758 20476 16764 20488
rect 16816 20476 16822 20528
rect 16960 20488 17448 20516
rect 13817 20451 13875 20457
rect 13817 20448 13829 20451
rect 13228 20420 13829 20448
rect 13228 20408 13234 20420
rect 13817 20417 13829 20420
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20448 14059 20451
rect 14090 20448 14096 20460
rect 14047 20420 14096 20448
rect 14047 20417 14059 20420
rect 14001 20411 14059 20417
rect 14090 20408 14096 20420
rect 14148 20408 14154 20460
rect 14550 20408 14556 20460
rect 14608 20448 14614 20460
rect 15105 20451 15163 20457
rect 15105 20448 15117 20451
rect 14608 20420 15117 20448
rect 14608 20408 14614 20420
rect 15105 20417 15117 20420
rect 15151 20417 15163 20451
rect 15105 20411 15163 20417
rect 15286 20408 15292 20460
rect 15344 20408 15350 20460
rect 16960 20457 16988 20488
rect 17420 20460 17448 20488
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20448 15531 20451
rect 15565 20451 15623 20457
rect 15565 20448 15577 20451
rect 15519 20420 15577 20448
rect 15519 20417 15531 20420
rect 15473 20411 15531 20417
rect 15565 20417 15577 20420
rect 15611 20417 15623 20451
rect 15565 20411 15623 20417
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 17126 20408 17132 20460
rect 17184 20408 17190 20460
rect 17402 20408 17408 20460
rect 17460 20408 17466 20460
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20417 17647 20451
rect 17696 20448 17724 20556
rect 18506 20544 18512 20596
rect 18564 20544 18570 20596
rect 20993 20587 21051 20593
rect 20993 20553 21005 20587
rect 21039 20584 21051 20587
rect 22738 20584 22744 20596
rect 21039 20556 22744 20584
rect 21039 20553 21051 20556
rect 20993 20547 21051 20553
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 23658 20544 23664 20596
rect 23716 20544 23722 20596
rect 23934 20544 23940 20596
rect 23992 20544 23998 20596
rect 24946 20593 24952 20596
rect 24923 20587 24952 20593
rect 24923 20584 24935 20587
rect 24136 20556 24935 20584
rect 22094 20525 22100 20528
rect 22066 20519 22100 20525
rect 22066 20485 22078 20519
rect 22066 20479 22100 20485
rect 22094 20476 22100 20479
rect 22152 20476 22158 20528
rect 23216 20488 23428 20516
rect 23216 20460 23244 20488
rect 17865 20451 17923 20457
rect 17865 20448 17877 20451
rect 17696 20420 17877 20448
rect 17589 20411 17647 20417
rect 17865 20417 17877 20420
rect 17911 20448 17923 20451
rect 18322 20448 18328 20460
rect 17911 20420 18328 20448
rect 17911 20417 17923 20420
rect 17865 20411 17923 20417
rect 12207 20352 12664 20380
rect 12207 20349 12219 20352
rect 12161 20343 12219 20349
rect 12802 20340 12808 20392
rect 12860 20380 12866 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12860 20352 13093 20380
rect 12860 20340 12866 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 16853 20383 16911 20389
rect 16853 20349 16865 20383
rect 16899 20380 16911 20383
rect 17144 20380 17172 20408
rect 16899 20352 17172 20380
rect 17313 20383 17371 20389
rect 16899 20349 16911 20352
rect 16853 20343 16911 20349
rect 17313 20349 17325 20383
rect 17359 20349 17371 20383
rect 17604 20380 17632 20411
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 18598 20408 18604 20460
rect 18656 20448 18662 20460
rect 19153 20451 19211 20457
rect 19153 20448 19165 20451
rect 18656 20420 19165 20448
rect 18656 20408 18662 20420
rect 19153 20417 19165 20420
rect 19199 20417 19211 20451
rect 19153 20411 19211 20417
rect 19334 20408 19340 20460
rect 19392 20408 19398 20460
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 20588 20420 20637 20448
rect 20588 20408 20594 20420
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20448 20867 20451
rect 20898 20448 20904 20460
rect 20855 20420 20904 20448
rect 20855 20417 20867 20420
rect 20809 20411 20867 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 21085 20451 21143 20457
rect 21085 20417 21097 20451
rect 21131 20448 21143 20451
rect 22554 20448 22560 20460
rect 21131 20420 22560 20448
rect 21131 20417 21143 20420
rect 21085 20411 21143 20417
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 23198 20408 23204 20460
rect 23256 20408 23262 20460
rect 23400 20457 23428 20488
rect 23474 20476 23480 20528
rect 23532 20516 23538 20528
rect 23569 20519 23627 20525
rect 23569 20516 23581 20519
rect 23532 20488 23581 20516
rect 23532 20476 23538 20488
rect 23569 20485 23581 20488
rect 23615 20485 23627 20519
rect 23676 20516 23704 20544
rect 24029 20519 24087 20525
rect 24029 20516 24041 20519
rect 23676 20488 24041 20516
rect 23569 20479 23627 20485
rect 24029 20485 24041 20488
rect 24075 20485 24087 20519
rect 24029 20479 24087 20485
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20417 23351 20451
rect 23293 20411 23351 20417
rect 23386 20451 23444 20457
rect 23386 20417 23398 20451
rect 23432 20417 23444 20451
rect 23386 20411 23444 20417
rect 17770 20380 17776 20392
rect 17604 20352 17776 20380
rect 17313 20343 17371 20349
rect 7929 20315 7987 20321
rect 7929 20281 7941 20315
rect 7975 20281 7987 20315
rect 7929 20275 7987 20281
rect 13446 20272 13452 20324
rect 13504 20312 13510 20324
rect 13633 20315 13691 20321
rect 13633 20312 13645 20315
rect 13504 20284 13645 20312
rect 13504 20272 13510 20284
rect 13633 20281 13645 20284
rect 13679 20281 13691 20315
rect 17328 20312 17356 20343
rect 17770 20340 17776 20352
rect 17828 20380 17834 20392
rect 19352 20380 19380 20408
rect 17828 20352 19380 20380
rect 21821 20383 21879 20389
rect 17828 20340 17834 20352
rect 21821 20349 21833 20383
rect 21867 20349 21879 20383
rect 21821 20343 21879 20349
rect 18601 20315 18659 20321
rect 18601 20312 18613 20315
rect 17328 20284 18613 20312
rect 13633 20275 13691 20281
rect 18601 20281 18613 20284
rect 18647 20281 18659 20315
rect 21634 20312 21640 20324
rect 18601 20275 18659 20281
rect 20364 20284 21640 20312
rect 8938 20244 8944 20256
rect 7668 20216 8944 20244
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 9769 20247 9827 20253
rect 9769 20244 9781 20247
rect 9456 20216 9781 20244
rect 9456 20204 9462 20216
rect 9769 20213 9781 20216
rect 9815 20213 9827 20247
rect 9769 20207 9827 20213
rect 13538 20204 13544 20256
rect 13596 20204 13602 20256
rect 15749 20247 15807 20253
rect 15749 20213 15761 20247
rect 15795 20244 15807 20247
rect 15930 20244 15936 20256
rect 15795 20216 15936 20244
rect 15795 20213 15807 20216
rect 15749 20207 15807 20213
rect 15930 20204 15936 20216
rect 15988 20204 15994 20256
rect 16945 20247 17003 20253
rect 16945 20213 16957 20247
rect 16991 20244 17003 20247
rect 17310 20244 17316 20256
rect 16991 20216 17316 20244
rect 16991 20213 17003 20216
rect 16945 20207 17003 20213
rect 17310 20204 17316 20216
rect 17368 20204 17374 20256
rect 17678 20204 17684 20256
rect 17736 20244 17742 20256
rect 17773 20247 17831 20253
rect 17773 20244 17785 20247
rect 17736 20216 17785 20244
rect 17736 20204 17742 20216
rect 17773 20213 17785 20216
rect 17819 20213 17831 20247
rect 17773 20207 17831 20213
rect 20254 20204 20260 20256
rect 20312 20244 20318 20256
rect 20364 20253 20392 20284
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 20349 20247 20407 20253
rect 20349 20244 20361 20247
rect 20312 20216 20361 20244
rect 20312 20204 20318 20216
rect 20349 20213 20361 20216
rect 20395 20213 20407 20247
rect 20349 20207 20407 20213
rect 20806 20204 20812 20256
rect 20864 20204 20870 20256
rect 21836 20244 21864 20343
rect 22922 20340 22928 20392
rect 22980 20380 22986 20392
rect 23308 20380 23336 20411
rect 23658 20408 23664 20460
rect 23716 20408 23722 20460
rect 23799 20451 23857 20457
rect 23799 20417 23811 20451
rect 23845 20448 23857 20451
rect 24136 20448 24164 20556
rect 24923 20553 24935 20556
rect 24923 20547 24952 20553
rect 24946 20544 24952 20547
rect 25004 20544 25010 20596
rect 25133 20519 25191 20525
rect 23845 20420 24164 20448
rect 24596 20488 24854 20516
rect 23845 20417 23857 20420
rect 23799 20411 23857 20417
rect 22980 20352 23336 20380
rect 22980 20340 22986 20352
rect 23566 20340 23572 20392
rect 23624 20380 23630 20392
rect 24596 20389 24624 20488
rect 24826 20448 24854 20488
rect 25133 20485 25145 20519
rect 25179 20485 25191 20519
rect 25133 20479 25191 20485
rect 25148 20448 25176 20479
rect 24826 20420 25176 20448
rect 24581 20383 24639 20389
rect 24581 20380 24593 20383
rect 23624 20352 24593 20380
rect 23624 20340 23630 20352
rect 24581 20349 24593 20352
rect 24627 20349 24639 20383
rect 24581 20343 24639 20349
rect 23201 20315 23259 20321
rect 23201 20281 23213 20315
rect 23247 20312 23259 20315
rect 23382 20312 23388 20324
rect 23247 20284 23388 20312
rect 23247 20281 23259 20284
rect 23201 20275 23259 20281
rect 23382 20272 23388 20284
rect 23440 20312 23446 20324
rect 23440 20284 24992 20312
rect 23440 20272 23446 20284
rect 22186 20244 22192 20256
rect 21836 20216 22192 20244
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 23474 20204 23480 20256
rect 23532 20244 23538 20256
rect 23658 20244 23664 20256
rect 23532 20216 23664 20244
rect 23532 20204 23538 20216
rect 23658 20204 23664 20216
rect 23716 20244 23722 20256
rect 24118 20244 24124 20256
rect 23716 20216 24124 20244
rect 23716 20204 23722 20216
rect 24118 20204 24124 20216
rect 24176 20244 24182 20256
rect 24964 20253 24992 20284
rect 24765 20247 24823 20253
rect 24765 20244 24777 20247
rect 24176 20216 24777 20244
rect 24176 20204 24182 20216
rect 24765 20213 24777 20216
rect 24811 20213 24823 20247
rect 24765 20207 24823 20213
rect 24949 20247 25007 20253
rect 24949 20213 24961 20247
rect 24995 20213 25007 20247
rect 24949 20207 25007 20213
rect 1104 20154 26496 20176
rect 1104 20102 4124 20154
rect 4176 20102 4188 20154
rect 4240 20102 4252 20154
rect 4304 20102 4316 20154
rect 4368 20102 4380 20154
rect 4432 20102 10472 20154
rect 10524 20102 10536 20154
rect 10588 20102 10600 20154
rect 10652 20102 10664 20154
rect 10716 20102 10728 20154
rect 10780 20102 16820 20154
rect 16872 20102 16884 20154
rect 16936 20102 16948 20154
rect 17000 20102 17012 20154
rect 17064 20102 17076 20154
rect 17128 20102 23168 20154
rect 23220 20102 23232 20154
rect 23284 20102 23296 20154
rect 23348 20102 23360 20154
rect 23412 20102 23424 20154
rect 23476 20102 26496 20154
rect 1104 20080 26496 20102
rect 7558 20000 7564 20052
rect 7616 20000 7622 20052
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 8021 20043 8079 20049
rect 8021 20040 8033 20043
rect 7984 20012 8033 20040
rect 7984 20000 7990 20012
rect 8021 20009 8033 20012
rect 8067 20009 8079 20043
rect 8021 20003 8079 20009
rect 8754 20000 8760 20052
rect 8812 20040 8818 20052
rect 9033 20043 9091 20049
rect 9033 20040 9045 20043
rect 8812 20012 9045 20040
rect 8812 20000 8818 20012
rect 9033 20009 9045 20012
rect 9079 20009 9091 20043
rect 9033 20003 9091 20009
rect 9214 20000 9220 20052
rect 9272 20040 9278 20052
rect 9585 20043 9643 20049
rect 9585 20040 9597 20043
rect 9272 20012 9597 20040
rect 9272 20000 9278 20012
rect 9585 20009 9597 20012
rect 9631 20009 9643 20043
rect 9585 20003 9643 20009
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 12618 20040 12624 20052
rect 10100 20012 12624 20040
rect 10100 20000 10106 20012
rect 12618 20000 12624 20012
rect 12676 20000 12682 20052
rect 15105 20043 15163 20049
rect 15105 20009 15117 20043
rect 15151 20040 15163 20043
rect 15286 20040 15292 20052
rect 15151 20012 15292 20040
rect 15151 20009 15163 20012
rect 15105 20003 15163 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 17129 20043 17187 20049
rect 17129 20040 17141 20043
rect 16632 20012 17141 20040
rect 16632 20000 16638 20012
rect 17129 20009 17141 20012
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 17402 20000 17408 20052
rect 17460 20000 17466 20052
rect 18598 20000 18604 20052
rect 18656 20040 18662 20052
rect 18785 20043 18843 20049
rect 18785 20040 18797 20043
rect 18656 20012 18797 20040
rect 18656 20000 18662 20012
rect 18785 20009 18797 20012
rect 18831 20009 18843 20043
rect 18785 20003 18843 20009
rect 20806 20000 20812 20052
rect 20864 20000 20870 20052
rect 20898 20000 20904 20052
rect 20956 20040 20962 20052
rect 21085 20043 21143 20049
rect 21085 20040 21097 20043
rect 20956 20012 21097 20040
rect 20956 20000 20962 20012
rect 21085 20009 21097 20012
rect 21131 20009 21143 20043
rect 21085 20003 21143 20009
rect 23566 20000 23572 20052
rect 23624 20000 23630 20052
rect 7576 19904 7604 20000
rect 9048 19944 9444 19972
rect 7576 19876 8156 19904
rect 7469 19839 7527 19845
rect 7469 19805 7481 19839
rect 7515 19805 7527 19839
rect 7469 19799 7527 19805
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 7650 19836 7656 19848
rect 7607 19808 7656 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 7484 19768 7512 19799
rect 7650 19796 7656 19808
rect 7708 19796 7714 19848
rect 8018 19768 8024 19780
rect 7484 19740 8024 19768
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7285 19703 7343 19709
rect 7285 19700 7297 19703
rect 7064 19672 7297 19700
rect 7064 19660 7070 19672
rect 7285 19669 7297 19672
rect 7331 19669 7343 19703
rect 7285 19663 7343 19669
rect 7926 19660 7932 19712
rect 7984 19660 7990 19712
rect 8128 19700 8156 19876
rect 8294 19864 8300 19916
rect 8352 19864 8358 19916
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 8312 19836 8340 19864
rect 8251 19808 8340 19836
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 8386 19796 8392 19848
rect 8444 19796 8450 19848
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 8846 19836 8852 19848
rect 8619 19808 8852 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 8846 19796 8852 19808
rect 8904 19796 8910 19848
rect 8938 19796 8944 19848
rect 8996 19796 9002 19848
rect 9048 19836 9076 19944
rect 9416 19904 9444 19944
rect 12434 19932 12440 19984
rect 12492 19972 12498 19984
rect 16945 19975 17003 19981
rect 12492 19944 12664 19972
rect 12492 19932 12498 19944
rect 10502 19904 10508 19916
rect 9416 19876 10508 19904
rect 9416 19848 9444 19876
rect 10502 19864 10508 19876
rect 10560 19864 10566 19916
rect 12636 19904 12664 19944
rect 16945 19941 16957 19975
rect 16991 19972 17003 19975
rect 17420 19972 17448 20000
rect 16991 19944 17448 19972
rect 16991 19941 17003 19944
rect 16945 19935 17003 19941
rect 14458 19904 14464 19916
rect 12636 19876 14464 19904
rect 14458 19864 14464 19876
rect 14516 19904 14522 19916
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 14516 19876 14841 19904
rect 14516 19864 14522 19876
rect 14829 19873 14841 19876
rect 14875 19873 14887 19907
rect 15657 19907 15715 19913
rect 15657 19904 15669 19907
rect 14829 19867 14887 19873
rect 14936 19876 15669 19904
rect 9116 19839 9174 19845
rect 9116 19836 9128 19839
rect 9048 19808 9128 19836
rect 9116 19805 9128 19808
rect 9162 19805 9174 19839
rect 9116 19799 9174 19805
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19830 9275 19839
rect 9306 19830 9312 19848
rect 9263 19805 9312 19830
rect 9217 19802 9312 19805
rect 9217 19799 9275 19802
rect 9306 19796 9312 19802
rect 9364 19796 9370 19848
rect 9398 19796 9404 19848
rect 9456 19796 9462 19848
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 9674 19796 9680 19848
rect 9732 19796 9738 19848
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19805 11115 19839
rect 11057 19799 11115 19805
rect 8297 19771 8355 19777
rect 8297 19737 8309 19771
rect 8343 19768 8355 19771
rect 9692 19768 9720 19796
rect 8343 19740 9720 19768
rect 11072 19768 11100 19799
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 12860 19808 13553 19836
rect 12860 19796 12866 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 14936 19836 14964 19876
rect 15657 19873 15669 19876
rect 15703 19873 15715 19907
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 15657 19867 15715 19873
rect 18984 19876 19625 19904
rect 18984 19848 19012 19876
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 19613 19867 19671 19873
rect 14700 19808 14964 19836
rect 14700 19796 14706 19808
rect 15102 19796 15108 19848
rect 15160 19836 15166 19848
rect 15841 19839 15899 19845
rect 15841 19836 15853 19839
rect 15160 19808 15853 19836
rect 15160 19796 15166 19808
rect 15841 19805 15853 19808
rect 15887 19836 15899 19839
rect 16298 19836 16304 19848
rect 15887 19808 16304 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 17678 19845 17684 19848
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 16592 19808 17417 19836
rect 16592 19780 16620 19808
rect 17405 19805 17417 19808
rect 17451 19805 17463 19839
rect 17672 19836 17684 19845
rect 17639 19808 17684 19836
rect 17405 19799 17463 19805
rect 17672 19799 17684 19808
rect 17678 19796 17684 19799
rect 17736 19796 17742 19848
rect 18966 19796 18972 19848
rect 19024 19796 19030 19848
rect 19337 19839 19395 19845
rect 19337 19805 19349 19839
rect 19383 19805 19395 19839
rect 19337 19799 19395 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19836 19579 19839
rect 20824 19836 20852 20000
rect 20993 19975 21051 19981
rect 20993 19941 21005 19975
rect 21039 19972 21051 19975
rect 21039 19944 21680 19972
rect 21039 19941 21051 19944
rect 20993 19935 21051 19941
rect 21652 19913 21680 19944
rect 21637 19907 21695 19913
rect 21637 19873 21649 19907
rect 21683 19873 21695 19907
rect 21637 19867 21695 19873
rect 22186 19864 22192 19916
rect 22244 19864 22250 19916
rect 19567 19808 20852 19836
rect 19567 19805 19579 19808
rect 19521 19799 19579 19805
rect 11238 19768 11244 19780
rect 11072 19740 11244 19768
rect 8343 19737 8355 19740
rect 8297 19731 8355 19737
rect 11238 19728 11244 19740
rect 11296 19728 11302 19780
rect 11333 19771 11391 19777
rect 11333 19737 11345 19771
rect 11379 19768 11391 19771
rect 11606 19768 11612 19780
rect 11379 19740 11612 19768
rect 11379 19737 11391 19740
rect 11333 19731 11391 19737
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 12618 19768 12624 19780
rect 12558 19740 12624 19768
rect 12618 19728 12624 19740
rect 12676 19728 12682 19780
rect 16574 19728 16580 19780
rect 16632 19728 16638 19780
rect 17313 19771 17371 19777
rect 17313 19737 17325 19771
rect 17359 19768 17371 19771
rect 18414 19768 18420 19780
rect 17359 19740 18420 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 18414 19728 18420 19740
rect 18472 19728 18478 19780
rect 9309 19703 9367 19709
rect 9309 19700 9321 19703
rect 8128 19672 9321 19700
rect 9309 19669 9321 19672
rect 9355 19669 9367 19703
rect 9309 19663 9367 19669
rect 12802 19660 12808 19712
rect 12860 19660 12866 19712
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 12989 19703 13047 19709
rect 12989 19700 13001 19703
rect 12952 19672 13001 19700
rect 12952 19660 12958 19672
rect 12989 19669 13001 19672
rect 13035 19669 13047 19703
rect 12989 19663 13047 19669
rect 13998 19660 14004 19712
rect 14056 19700 14062 19712
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 14056 19672 14289 19700
rect 14056 19660 14062 19672
rect 14277 19669 14289 19672
rect 14323 19669 14335 19703
rect 14277 19663 14335 19669
rect 14737 19703 14795 19709
rect 14737 19669 14749 19703
rect 14783 19700 14795 19703
rect 15194 19700 15200 19712
rect 14783 19672 15200 19700
rect 14783 19669 14795 19672
rect 14737 19663 14795 19669
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 16666 19660 16672 19712
rect 16724 19700 16730 19712
rect 17113 19703 17171 19709
rect 17113 19700 17125 19703
rect 16724 19672 17125 19700
rect 16724 19660 16730 19672
rect 17113 19669 17125 19672
rect 17159 19700 17171 19703
rect 17494 19700 17500 19712
rect 17159 19672 17500 19700
rect 17159 19669 17171 19672
rect 17113 19663 17171 19669
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 17586 19660 17592 19712
rect 17644 19700 17650 19712
rect 19352 19700 19380 19799
rect 19429 19771 19487 19777
rect 19429 19737 19441 19771
rect 19475 19768 19487 19771
rect 19858 19771 19916 19777
rect 19858 19768 19870 19771
rect 19475 19740 19870 19768
rect 19475 19737 19487 19740
rect 19429 19731 19487 19737
rect 19858 19737 19870 19740
rect 19904 19737 19916 19771
rect 19858 19731 19916 19737
rect 22456 19771 22514 19777
rect 22456 19737 22468 19771
rect 22502 19768 22514 19771
rect 22738 19768 22744 19780
rect 22502 19740 22744 19768
rect 22502 19737 22514 19740
rect 22456 19731 22514 19737
rect 22738 19728 22744 19740
rect 22796 19728 22802 19780
rect 20254 19700 20260 19712
rect 17644 19672 20260 19700
rect 17644 19660 17650 19672
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 1104 19610 26656 19632
rect 1104 19558 7298 19610
rect 7350 19558 7362 19610
rect 7414 19558 7426 19610
rect 7478 19558 7490 19610
rect 7542 19558 7554 19610
rect 7606 19558 13646 19610
rect 13698 19558 13710 19610
rect 13762 19558 13774 19610
rect 13826 19558 13838 19610
rect 13890 19558 13902 19610
rect 13954 19558 19994 19610
rect 20046 19558 20058 19610
rect 20110 19558 20122 19610
rect 20174 19558 20186 19610
rect 20238 19558 20250 19610
rect 20302 19558 26342 19610
rect 26394 19558 26406 19610
rect 26458 19558 26470 19610
rect 26522 19558 26534 19610
rect 26586 19558 26598 19610
rect 26650 19558 26656 19610
rect 1104 19536 26656 19558
rect 7377 19499 7435 19505
rect 7377 19465 7389 19499
rect 7423 19496 7435 19499
rect 7650 19496 7656 19508
rect 7423 19468 7656 19496
rect 7423 19465 7435 19468
rect 7377 19459 7435 19465
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 7926 19456 7932 19508
rect 7984 19496 7990 19508
rect 8113 19499 8171 19505
rect 8113 19496 8125 19499
rect 7984 19468 8125 19496
rect 7984 19456 7990 19468
rect 8113 19465 8125 19468
rect 8159 19465 8171 19499
rect 8113 19459 8171 19465
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 8938 19456 8944 19508
rect 8996 19496 9002 19508
rect 9033 19499 9091 19505
rect 9033 19496 9045 19499
rect 8996 19468 9045 19496
rect 8996 19456 9002 19468
rect 9033 19465 9045 19468
rect 9079 19496 9091 19499
rect 9122 19496 9128 19508
rect 9079 19468 9128 19496
rect 9079 19465 9091 19468
rect 9033 19459 9091 19465
rect 9122 19456 9128 19468
rect 9180 19496 9186 19508
rect 9490 19496 9496 19508
rect 9180 19468 9496 19496
rect 9180 19456 9186 19468
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 9677 19499 9735 19505
rect 9677 19465 9689 19499
rect 9723 19465 9735 19499
rect 9950 19496 9956 19508
rect 9677 19459 9735 19465
rect 9784 19468 9956 19496
rect 8772 19428 8800 19456
rect 8496 19400 8800 19428
rect 9217 19431 9275 19437
rect 1762 19320 1768 19372
rect 1820 19320 1826 19372
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19360 6423 19363
rect 7098 19360 7104 19372
rect 6411 19332 7104 19360
rect 6411 19329 6423 19332
rect 6365 19323 6423 19329
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 8496 19369 8524 19400
rect 9217 19397 9229 19431
rect 9263 19428 9275 19431
rect 9398 19428 9404 19440
rect 9263 19400 9404 19428
rect 9263 19397 9275 19400
rect 9217 19391 9275 19397
rect 9398 19388 9404 19400
rect 9456 19388 9462 19440
rect 9692 19428 9720 19459
rect 9508 19400 9720 19428
rect 9508 19372 9536 19400
rect 8297 19363 8355 19369
rect 8297 19329 8309 19363
rect 8343 19329 8355 19363
rect 8297 19323 8355 19329
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19329 8539 19363
rect 8481 19323 8539 19329
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19360 8815 19363
rect 9030 19360 9036 19372
rect 8803 19332 9036 19360
rect 8803 19329 8815 19332
rect 8757 19323 8815 19329
rect 8021 19295 8079 19301
rect 8021 19261 8033 19295
rect 8067 19292 8079 19295
rect 8312 19292 8340 19323
rect 9030 19320 9036 19332
rect 9088 19320 9094 19372
rect 9125 19363 9183 19369
rect 9125 19329 9137 19363
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 8386 19292 8392 19304
rect 8067 19264 8392 19292
rect 8067 19261 8079 19264
rect 8021 19255 8079 19261
rect 8386 19252 8392 19264
rect 8444 19292 8450 19304
rect 9140 19292 9168 19323
rect 9490 19320 9496 19372
rect 9548 19320 9554 19372
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9784 19360 9812 19468
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 12526 19496 12532 19508
rect 12347 19468 12532 19496
rect 11517 19431 11575 19437
rect 9876 19400 11468 19428
rect 9876 19369 9904 19400
rect 11440 19372 11468 19400
rect 11517 19397 11529 19431
rect 11563 19428 11575 19431
rect 11606 19428 11612 19440
rect 11563 19400 11612 19428
rect 11563 19397 11575 19400
rect 11517 19391 11575 19397
rect 11606 19388 11612 19400
rect 11664 19388 11670 19440
rect 11882 19388 11888 19440
rect 11940 19428 11946 19440
rect 12347 19428 12375 19468
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 12621 19499 12679 19505
rect 12621 19465 12633 19499
rect 12667 19496 12679 19499
rect 13170 19496 13176 19508
rect 12667 19468 13176 19496
rect 12667 19465 12679 19468
rect 12621 19459 12679 19465
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 14384 19468 16252 19496
rect 11940 19400 12375 19428
rect 11940 19388 11946 19400
rect 9723 19332 9812 19360
rect 9861 19363 9919 19369
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 9861 19329 9873 19363
rect 9907 19329 9919 19363
rect 9861 19323 9919 19329
rect 9953 19363 10011 19369
rect 9953 19329 9965 19363
rect 9999 19329 10011 19363
rect 9953 19323 10011 19329
rect 10229 19363 10287 19369
rect 10229 19329 10241 19363
rect 10275 19360 10287 19363
rect 10318 19360 10324 19372
rect 10275 19332 10324 19360
rect 10275 19329 10287 19332
rect 10229 19323 10287 19329
rect 9968 19292 9996 19323
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 10502 19320 10508 19372
rect 10560 19320 10566 19372
rect 10597 19363 10655 19369
rect 10597 19329 10609 19363
rect 10643 19360 10655 19363
rect 11054 19360 11060 19372
rect 10643 19332 11060 19360
rect 10643 19329 10655 19332
rect 10597 19323 10655 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 11146 19320 11152 19372
rect 11204 19320 11210 19372
rect 11330 19320 11336 19372
rect 11388 19320 11394 19372
rect 11422 19320 11428 19372
rect 11480 19360 11486 19372
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11480 19332 11713 19360
rect 11480 19320 11486 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19329 11851 19363
rect 11793 19323 11851 19329
rect 10137 19295 10195 19301
rect 8444 19264 9536 19292
rect 9968 19264 10088 19292
rect 8444 19252 8450 19264
rect 9030 19184 9036 19236
rect 9088 19224 9094 19236
rect 9401 19227 9459 19233
rect 9401 19224 9413 19227
rect 9088 19196 9413 19224
rect 9088 19184 9094 19196
rect 9401 19193 9413 19196
rect 9447 19193 9459 19227
rect 9508 19224 9536 19264
rect 10060 19224 10088 19264
rect 10137 19261 10149 19295
rect 10183 19292 10195 19295
rect 10870 19292 10876 19304
rect 10183 19264 10876 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 10965 19295 11023 19301
rect 10965 19261 10977 19295
rect 11011 19292 11023 19295
rect 11808 19292 11836 19323
rect 11974 19320 11980 19372
rect 12032 19369 12038 19372
rect 12032 19363 12061 19369
rect 12049 19329 12061 19363
rect 12032 19323 12061 19329
rect 12032 19320 12038 19323
rect 12250 19320 12256 19372
rect 12308 19320 12314 19372
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12434 19360 12440 19372
rect 12400 19332 12440 19360
rect 12400 19320 12406 19332
rect 12434 19320 12440 19332
rect 12492 19360 12498 19372
rect 12492 19332 12537 19360
rect 12492 19320 12498 19332
rect 12618 19320 12624 19372
rect 12676 19360 12682 19372
rect 14384 19369 14412 19468
rect 14369 19363 14427 19369
rect 12676 19332 13018 19360
rect 12676 19320 12682 19332
rect 14369 19329 14381 19363
rect 14415 19329 14427 19363
rect 14918 19360 14924 19372
rect 14858 19332 14924 19360
rect 14369 19323 14427 19329
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 11011 19264 11836 19292
rect 11011 19261 11023 19264
rect 10965 19255 11023 19261
rect 11882 19252 11888 19304
rect 11940 19292 11946 19304
rect 11992 19292 12020 19320
rect 11940 19264 12020 19292
rect 12161 19295 12219 19301
rect 11940 19252 11946 19264
rect 12161 19261 12173 19295
rect 12207 19292 12219 19295
rect 12894 19292 12900 19304
rect 12207 19264 12900 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 13354 19252 13360 19304
rect 13412 19292 13418 19304
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13412 19264 14105 19292
rect 13412 19252 13418 19264
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 15470 19252 15476 19304
rect 15528 19292 15534 19304
rect 16224 19301 16252 19468
rect 16482 19456 16488 19508
rect 16540 19496 16546 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 16540 19468 18337 19496
rect 16540 19456 16546 19468
rect 18325 19465 18337 19468
rect 18371 19465 18383 19499
rect 18325 19459 18383 19465
rect 18506 19456 18512 19508
rect 18564 19456 18570 19508
rect 18984 19468 21220 19496
rect 17120 19431 17178 19437
rect 17120 19397 17132 19431
rect 17166 19428 17178 19431
rect 17218 19428 17224 19440
rect 17166 19400 17224 19428
rect 17166 19397 17178 19400
rect 17120 19391 17178 19397
rect 17218 19388 17224 19400
rect 17276 19388 17282 19440
rect 18322 19360 18328 19372
rect 18248 19332 18328 19360
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15528 19264 15945 19292
rect 15528 19252 15534 19264
rect 15933 19261 15945 19264
rect 15979 19261 15991 19295
rect 15933 19255 15991 19261
rect 16209 19295 16267 19301
rect 16209 19261 16221 19295
rect 16255 19292 16267 19295
rect 16574 19292 16580 19304
rect 16255 19264 16580 19292
rect 16255 19261 16267 19264
rect 16209 19255 16267 19261
rect 16574 19252 16580 19264
rect 16632 19292 16638 19304
rect 16853 19295 16911 19301
rect 16853 19292 16865 19295
rect 16632 19264 16865 19292
rect 16632 19252 16638 19264
rect 16853 19261 16865 19264
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 10226 19224 10232 19236
rect 9508 19196 10232 19224
rect 9401 19187 9459 19193
rect 934 19116 940 19168
rect 992 19156 998 19168
rect 1489 19159 1547 19165
rect 1489 19156 1501 19159
rect 992 19128 1501 19156
rect 992 19116 998 19128
rect 1489 19125 1501 19128
rect 1535 19125 1547 19159
rect 1489 19119 1547 19125
rect 6546 19116 6552 19168
rect 6604 19116 6610 19168
rect 8478 19116 8484 19168
rect 8536 19116 8542 19168
rect 8570 19116 8576 19168
rect 8628 19156 8634 19168
rect 8849 19159 8907 19165
rect 8849 19156 8861 19159
rect 8628 19128 8861 19156
rect 8628 19116 8634 19128
rect 8849 19125 8861 19128
rect 8895 19125 8907 19159
rect 9416 19156 9444 19187
rect 10226 19184 10232 19196
rect 10284 19184 10290 19236
rect 10410 19184 10416 19236
rect 10468 19184 10474 19236
rect 11330 19184 11336 19236
rect 11388 19224 11394 19236
rect 12342 19224 12348 19236
rect 11388 19196 12348 19224
rect 11388 19184 11394 19196
rect 12342 19184 12348 19196
rect 12400 19184 12406 19236
rect 18248 19233 18276 19332
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18414 19320 18420 19372
rect 18472 19320 18478 19372
rect 18524 19360 18552 19456
rect 18984 19440 19012 19468
rect 18966 19388 18972 19440
rect 19024 19388 19030 19440
rect 20898 19388 20904 19440
rect 20956 19428 20962 19440
rect 20993 19431 21051 19437
rect 20993 19428 21005 19431
rect 20956 19400 21005 19428
rect 20956 19388 20962 19400
rect 20993 19397 21005 19400
rect 21039 19397 21051 19431
rect 21192 19428 21220 19468
rect 21634 19456 21640 19508
rect 21692 19496 21698 19508
rect 21692 19468 22508 19496
rect 21692 19456 21698 19468
rect 22480 19437 22508 19468
rect 22738 19456 22744 19508
rect 22796 19456 22802 19508
rect 22465 19431 22523 19437
rect 21192 19400 21312 19428
rect 20993 19391 21051 19397
rect 21284 19369 21312 19400
rect 22465 19397 22477 19431
rect 22511 19397 22523 19431
rect 22465 19391 22523 19397
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 18524 19332 19073 19360
rect 19061 19329 19073 19332
rect 19107 19329 19119 19363
rect 21269 19363 21327 19369
rect 19061 19323 19119 19329
rect 18432 19292 18460 19320
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 18432 19264 18889 19292
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19904 19292 19932 19346
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 22186 19360 22192 19372
rect 21315 19332 22192 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22741 19363 22799 19369
rect 22741 19329 22753 19363
rect 22787 19360 22799 19363
rect 23658 19360 23664 19372
rect 22787 19332 23664 19360
rect 22787 19329 22799 19332
rect 22741 19323 22799 19329
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 19392 19264 19932 19292
rect 22649 19295 22707 19301
rect 19392 19252 19398 19264
rect 22649 19261 22661 19295
rect 22695 19292 22707 19295
rect 22830 19292 22836 19304
rect 22695 19264 22836 19292
rect 22695 19261 22707 19264
rect 22649 19255 22707 19261
rect 22830 19252 22836 19264
rect 22888 19252 22894 19304
rect 18233 19227 18291 19233
rect 18233 19193 18245 19227
rect 18279 19193 18291 19227
rect 18233 19187 18291 19193
rect 18322 19184 18328 19236
rect 18380 19224 18386 19236
rect 19521 19227 19579 19233
rect 18380 19196 19288 19224
rect 18380 19184 18386 19196
rect 9582 19156 9588 19168
rect 9416 19128 9588 19156
rect 8849 19119 8907 19125
rect 9582 19116 9588 19128
rect 9640 19156 9646 19168
rect 10137 19159 10195 19165
rect 10137 19156 10149 19159
rect 9640 19128 10149 19156
rect 9640 19116 9646 19128
rect 10137 19125 10149 19128
rect 10183 19156 10195 19159
rect 12066 19156 12072 19168
rect 10183 19128 12072 19156
rect 10183 19125 10195 19128
rect 10137 19119 10195 19125
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 12253 19159 12311 19165
rect 12253 19156 12265 19159
rect 12216 19128 12265 19156
rect 12216 19116 12222 19128
rect 12253 19125 12265 19128
rect 12299 19125 12311 19159
rect 12253 19119 12311 19125
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 14090 19156 14096 19168
rect 13688 19128 14096 19156
rect 13688 19116 13694 19128
rect 14090 19116 14096 19128
rect 14148 19116 14154 19168
rect 14461 19159 14519 19165
rect 14461 19125 14473 19159
rect 14507 19156 14519 19159
rect 15194 19156 15200 19168
rect 14507 19128 15200 19156
rect 14507 19125 14519 19128
rect 14461 19119 14519 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 17494 19116 17500 19168
rect 17552 19156 17558 19168
rect 19260 19165 19288 19196
rect 19521 19193 19533 19227
rect 19567 19224 19579 19227
rect 19794 19224 19800 19236
rect 19567 19196 19800 19224
rect 19567 19193 19579 19196
rect 19521 19187 19579 19193
rect 19794 19184 19800 19196
rect 19852 19184 19858 19236
rect 19153 19159 19211 19165
rect 19153 19156 19165 19159
rect 17552 19128 19165 19156
rect 17552 19116 17558 19128
rect 19153 19125 19165 19128
rect 19199 19125 19211 19159
rect 19153 19119 19211 19125
rect 19245 19159 19303 19165
rect 19245 19125 19257 19159
rect 19291 19125 19303 19159
rect 19245 19119 19303 19125
rect 1104 19066 26496 19088
rect 1104 19014 4124 19066
rect 4176 19014 4188 19066
rect 4240 19014 4252 19066
rect 4304 19014 4316 19066
rect 4368 19014 4380 19066
rect 4432 19014 10472 19066
rect 10524 19014 10536 19066
rect 10588 19014 10600 19066
rect 10652 19014 10664 19066
rect 10716 19014 10728 19066
rect 10780 19014 16820 19066
rect 16872 19014 16884 19066
rect 16936 19014 16948 19066
rect 17000 19014 17012 19066
rect 17064 19014 17076 19066
rect 17128 19014 23168 19066
rect 23220 19014 23232 19066
rect 23284 19014 23296 19066
rect 23348 19014 23360 19066
rect 23412 19014 23424 19066
rect 23476 19014 26496 19066
rect 1104 18992 26496 19014
rect 7098 18912 7104 18964
rect 7156 18952 7162 18964
rect 7929 18955 7987 18961
rect 7929 18952 7941 18955
rect 7156 18924 7941 18952
rect 7156 18912 7162 18924
rect 7929 18921 7941 18924
rect 7975 18921 7987 18955
rect 7929 18915 7987 18921
rect 8386 18912 8392 18964
rect 8444 18912 8450 18964
rect 9490 18952 9496 18964
rect 9324 18924 9496 18952
rect 7837 18887 7895 18893
rect 7837 18853 7849 18887
rect 7883 18884 7895 18887
rect 8404 18884 8432 18912
rect 7883 18856 8432 18884
rect 7883 18853 7895 18856
rect 7837 18847 7895 18853
rect 6089 18819 6147 18825
rect 6089 18785 6101 18819
rect 6135 18816 6147 18819
rect 6362 18816 6368 18828
rect 6135 18788 6368 18816
rect 6135 18785 6147 18788
rect 6089 18779 6147 18785
rect 6362 18776 6368 18788
rect 6420 18776 6426 18828
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 8352 18788 8401 18816
rect 8352 18776 8358 18788
rect 8389 18785 8401 18788
rect 8435 18785 8447 18819
rect 8389 18779 8447 18785
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18785 8539 18819
rect 8481 18779 8539 18785
rect 8496 18748 8524 18779
rect 8128 18720 8524 18748
rect 6365 18683 6423 18689
rect 6365 18649 6377 18683
rect 6411 18649 6423 18683
rect 6365 18643 6423 18649
rect 6380 18612 6408 18643
rect 6914 18640 6920 18692
rect 6972 18640 6978 18692
rect 8128 18624 8156 18720
rect 8662 18708 8668 18760
rect 8720 18708 8726 18760
rect 9214 18708 9220 18760
rect 9272 18708 9278 18760
rect 9324 18757 9352 18924
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 12434 18952 12440 18964
rect 11204 18924 12296 18952
rect 11204 18912 11210 18924
rect 11698 18884 11704 18896
rect 9416 18856 11704 18884
rect 9416 18760 9444 18856
rect 11698 18844 11704 18856
rect 11756 18844 11762 18896
rect 11882 18844 11888 18896
rect 11940 18844 11946 18896
rect 12268 18884 12296 18924
rect 12360 18924 12440 18952
rect 12360 18884 12388 18924
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12529 18955 12587 18961
rect 12529 18921 12541 18955
rect 12575 18952 12587 18955
rect 13354 18952 13360 18964
rect 12575 18924 13360 18952
rect 12575 18921 12587 18924
rect 12529 18915 12587 18921
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 13538 18912 13544 18964
rect 13596 18912 13602 18964
rect 14461 18955 14519 18961
rect 14461 18921 14473 18955
rect 14507 18952 14519 18955
rect 14642 18952 14648 18964
rect 14507 18924 14648 18952
rect 14507 18921 14519 18924
rect 14461 18915 14519 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 18414 18912 18420 18964
rect 18472 18912 18478 18964
rect 12268 18856 12388 18884
rect 12452 18884 12480 18912
rect 12710 18884 12716 18896
rect 12452 18856 12716 18884
rect 12710 18844 12716 18856
rect 12768 18844 12774 18896
rect 11900 18816 11928 18844
rect 11900 18788 12388 18816
rect 12360 18760 12388 18788
rect 12618 18776 12624 18828
rect 12676 18816 12682 18828
rect 13449 18819 13507 18825
rect 13449 18816 13461 18819
rect 12676 18788 13461 18816
rect 12676 18776 12682 18788
rect 13449 18785 13461 18788
rect 13495 18785 13507 18819
rect 13556 18816 13584 18912
rect 14274 18884 14280 18896
rect 14108 18856 14280 18884
rect 14108 18825 14136 18856
rect 14274 18844 14280 18856
rect 14332 18844 14338 18896
rect 19334 18844 19340 18896
rect 19392 18884 19398 18896
rect 20349 18887 20407 18893
rect 20349 18884 20361 18887
rect 19392 18856 20361 18884
rect 19392 18844 19398 18856
rect 20349 18853 20361 18856
rect 20395 18853 20407 18887
rect 20349 18847 20407 18853
rect 13725 18819 13783 18825
rect 13725 18816 13737 18819
rect 13556 18788 13737 18816
rect 13449 18779 13507 18785
rect 13725 18785 13737 18788
rect 13771 18785 13783 18819
rect 13725 18779 13783 18785
rect 14093 18819 14151 18825
rect 14093 18785 14105 18819
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 14292 18788 14688 18816
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9677 18751 9735 18757
rect 9677 18717 9689 18751
rect 9723 18748 9735 18751
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9723 18720 9781 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 10410 18708 10416 18760
rect 10468 18708 10474 18760
rect 11146 18708 11152 18760
rect 11204 18748 11210 18760
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 11204 18720 11989 18748
rect 11204 18708 11210 18720
rect 11977 18717 11989 18720
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 8202 18640 8208 18692
rect 8260 18680 8266 18692
rect 8680 18680 8708 18708
rect 9519 18683 9577 18689
rect 9519 18680 9531 18683
rect 8260 18652 9531 18680
rect 8260 18640 8266 18652
rect 9519 18649 9531 18652
rect 9565 18649 9577 18683
rect 9519 18643 9577 18649
rect 9858 18640 9864 18692
rect 9916 18680 9922 18692
rect 10505 18683 10563 18689
rect 10505 18680 10517 18683
rect 9916 18652 10517 18680
rect 9916 18640 9922 18652
rect 10505 18649 10517 18652
rect 10551 18649 10563 18683
rect 10505 18643 10563 18649
rect 11238 18640 11244 18692
rect 11296 18640 11302 18692
rect 7006 18612 7012 18624
rect 6380 18584 7012 18612
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 8110 18572 8116 18624
rect 8168 18572 8174 18624
rect 8294 18572 8300 18624
rect 8352 18572 8358 18624
rect 9030 18572 9036 18624
rect 9088 18572 9094 18624
rect 11992 18612 12020 18711
rect 12342 18708 12348 18760
rect 12400 18708 12406 18760
rect 13170 18708 13176 18760
rect 13228 18708 13234 18760
rect 13538 18708 13544 18760
rect 13596 18708 13602 18760
rect 14292 18757 14320 18788
rect 14660 18760 14688 18788
rect 15930 18776 15936 18828
rect 15988 18776 15994 18828
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18717 14335 18751
rect 14277 18711 14335 18717
rect 12158 18640 12164 18692
rect 12216 18640 12222 18692
rect 12253 18683 12311 18689
rect 12253 18649 12265 18683
rect 12299 18680 12311 18683
rect 12621 18683 12679 18689
rect 12621 18680 12633 18683
rect 12299 18652 12633 18680
rect 12299 18649 12311 18652
rect 12253 18643 12311 18649
rect 12621 18649 12633 18652
rect 12667 18649 12679 18683
rect 12621 18643 12679 18649
rect 13078 18640 13084 18692
rect 13136 18680 13142 18692
rect 13648 18680 13676 18711
rect 14366 18708 14372 18760
rect 14424 18708 14430 18760
rect 14642 18708 14648 18760
rect 14700 18708 14706 18760
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18748 16267 18751
rect 16574 18748 16580 18760
rect 16255 18720 16580 18748
rect 16255 18717 16267 18720
rect 16209 18711 16267 18717
rect 16574 18708 16580 18720
rect 16632 18748 16638 18760
rect 17310 18757 17316 18760
rect 17037 18751 17095 18757
rect 17037 18748 17049 18751
rect 16632 18720 17049 18748
rect 16632 18708 16638 18720
rect 17037 18717 17049 18720
rect 17083 18717 17095 18751
rect 17304 18748 17316 18757
rect 17271 18720 17316 18748
rect 17037 18711 17095 18717
rect 17304 18711 17316 18720
rect 17310 18708 17316 18711
rect 17368 18708 17374 18760
rect 20165 18751 20223 18757
rect 20165 18717 20177 18751
rect 20211 18748 20223 18751
rect 20346 18748 20352 18760
rect 20211 18720 20352 18748
rect 20211 18717 20223 18720
rect 20165 18711 20223 18717
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18748 20499 18751
rect 20714 18748 20720 18760
rect 20487 18720 20720 18748
rect 20487 18717 20499 18720
rect 20441 18711 20499 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 22830 18708 22836 18760
rect 22888 18708 22894 18760
rect 14182 18680 14188 18692
rect 13136 18652 13676 18680
rect 13924 18652 14188 18680
rect 13136 18640 13142 18652
rect 13446 18612 13452 18624
rect 11992 18584 13452 18612
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 13924 18621 13952 18652
rect 14182 18640 14188 18652
rect 14240 18640 14246 18692
rect 15654 18680 15660 18692
rect 15502 18652 15660 18680
rect 13909 18615 13967 18621
rect 13909 18581 13921 18615
rect 13955 18581 13967 18615
rect 13909 18575 13967 18581
rect 14090 18572 14096 18624
rect 14148 18572 14154 18624
rect 14918 18572 14924 18624
rect 14976 18612 14982 18624
rect 15580 18612 15608 18652
rect 15654 18640 15660 18652
rect 15712 18680 15718 18692
rect 17494 18680 17500 18692
rect 15712 18652 17500 18680
rect 15712 18640 15718 18652
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 14976 18584 15608 18612
rect 14976 18572 14982 18584
rect 19702 18572 19708 18624
rect 19760 18612 19766 18624
rect 19981 18615 20039 18621
rect 19981 18612 19993 18615
rect 19760 18584 19993 18612
rect 19760 18572 19766 18584
rect 19981 18581 19993 18584
rect 20027 18581 20039 18615
rect 19981 18575 20039 18581
rect 23017 18615 23075 18621
rect 23017 18581 23029 18615
rect 23063 18612 23075 18615
rect 23290 18612 23296 18624
rect 23063 18584 23296 18612
rect 23063 18581 23075 18584
rect 23017 18575 23075 18581
rect 23290 18572 23296 18584
rect 23348 18572 23354 18624
rect 1104 18522 26656 18544
rect 1104 18470 7298 18522
rect 7350 18470 7362 18522
rect 7414 18470 7426 18522
rect 7478 18470 7490 18522
rect 7542 18470 7554 18522
rect 7606 18470 13646 18522
rect 13698 18470 13710 18522
rect 13762 18470 13774 18522
rect 13826 18470 13838 18522
rect 13890 18470 13902 18522
rect 13954 18470 19994 18522
rect 20046 18470 20058 18522
rect 20110 18470 20122 18522
rect 20174 18470 20186 18522
rect 20238 18470 20250 18522
rect 20302 18470 26342 18522
rect 26394 18470 26406 18522
rect 26458 18470 26470 18522
rect 26522 18470 26534 18522
rect 26586 18470 26598 18522
rect 26650 18470 26656 18522
rect 1104 18448 26656 18470
rect 1762 18368 1768 18420
rect 1820 18408 1826 18420
rect 2133 18411 2191 18417
rect 2133 18408 2145 18411
rect 1820 18380 2145 18408
rect 1820 18368 1826 18380
rect 2133 18377 2145 18380
rect 2179 18377 2191 18411
rect 2133 18371 2191 18377
rect 8110 18368 8116 18420
rect 8168 18368 8174 18420
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 8294 18408 8300 18420
rect 8251 18380 8300 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 11238 18408 11244 18420
rect 8680 18380 11244 18408
rect 6546 18300 6552 18352
rect 6604 18340 6610 18352
rect 6641 18343 6699 18349
rect 6641 18340 6653 18343
rect 6604 18312 6653 18340
rect 6604 18300 6610 18312
rect 6641 18309 6653 18312
rect 6687 18309 6699 18343
rect 6641 18303 6699 18309
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 7926 18272 7932 18284
rect 2363 18244 2774 18272
rect 7774 18244 7932 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 2746 18068 2774 18244
rect 7926 18232 7932 18244
rect 7984 18232 7990 18284
rect 6362 18164 6368 18216
rect 6420 18164 6426 18216
rect 7098 18068 7104 18080
rect 2746 18040 7104 18068
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 8128 18068 8156 18368
rect 8570 18300 8576 18352
rect 8628 18300 8634 18352
rect 8389 18275 8447 18281
rect 8389 18241 8401 18275
rect 8435 18272 8447 18275
rect 8588 18272 8616 18300
rect 8680 18281 8708 18380
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 11422 18368 11428 18420
rect 11480 18408 11486 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 11480 18380 12173 18408
rect 11480 18368 11486 18380
rect 12161 18377 12173 18380
rect 12207 18377 12219 18411
rect 12161 18371 12219 18377
rect 14090 18368 14096 18420
rect 14148 18368 14154 18420
rect 14366 18368 14372 18420
rect 14424 18368 14430 18420
rect 15105 18411 15163 18417
rect 15105 18377 15117 18411
rect 15151 18408 15163 18411
rect 15470 18408 15476 18420
rect 15151 18380 15476 18408
rect 15151 18377 15163 18380
rect 15105 18371 15163 18377
rect 15470 18368 15476 18380
rect 15528 18368 15534 18420
rect 19702 18368 19708 18420
rect 19760 18368 19766 18420
rect 22066 18380 23520 18408
rect 8941 18343 8999 18349
rect 8941 18309 8953 18343
rect 8987 18340 8999 18343
rect 9030 18340 9036 18352
rect 8987 18312 9036 18340
rect 8987 18309 8999 18312
rect 8941 18303 8999 18309
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 12434 18340 12440 18352
rect 10244 18312 11284 18340
rect 8435 18244 8616 18272
rect 8665 18275 8723 18281
rect 8435 18241 8447 18244
rect 8389 18235 8447 18241
rect 8665 18241 8677 18275
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 9950 18232 9956 18284
rect 10008 18232 10014 18284
rect 10042 18232 10048 18284
rect 10100 18232 10106 18284
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 8938 18204 8944 18216
rect 8619 18176 8944 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 8938 18164 8944 18176
rect 8996 18204 9002 18216
rect 9398 18204 9404 18216
rect 8996 18176 9404 18204
rect 8996 18164 9002 18176
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9968 18204 9996 18232
rect 10244 18204 10272 18312
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 10376 18244 10517 18272
rect 10376 18232 10382 18244
rect 10505 18241 10517 18244
rect 10551 18241 10563 18275
rect 10505 18235 10563 18241
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 10686 18272 10692 18284
rect 10643 18244 10692 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 10612 18204 10640 18235
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 10781 18275 10839 18281
rect 10781 18241 10793 18275
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 10881 18275 10939 18281
rect 10881 18241 10893 18275
rect 10927 18272 10939 18275
rect 10980 18272 11008 18312
rect 10927 18244 11008 18272
rect 10927 18241 10939 18244
rect 10881 18235 10939 18241
rect 9968 18176 10272 18204
rect 10336 18176 10640 18204
rect 10796 18204 10824 18235
rect 11054 18232 11060 18284
rect 11112 18232 11118 18284
rect 11256 18281 11284 18312
rect 12176 18312 12440 18340
rect 11241 18275 11299 18281
rect 11241 18241 11253 18275
rect 11287 18241 11299 18275
rect 11241 18235 11299 18241
rect 11330 18232 11336 18284
rect 11388 18232 11394 18284
rect 12066 18232 12072 18284
rect 12124 18232 12130 18284
rect 12176 18281 12204 18312
rect 12434 18300 12440 18312
rect 12492 18340 12498 18352
rect 12492 18312 13216 18340
rect 12492 18300 12498 18312
rect 12161 18275 12219 18281
rect 12161 18241 12173 18275
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 10962 18204 10968 18216
rect 10796 18176 10968 18204
rect 10336 18068 10364 18176
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 11072 18204 11100 18232
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 11072 18176 11805 18204
rect 11793 18173 11805 18176
rect 11839 18173 11851 18207
rect 11793 18167 11851 18173
rect 10410 18096 10416 18148
rect 10468 18136 10474 18148
rect 11330 18136 11336 18148
rect 10468 18108 11336 18136
rect 10468 18096 10474 18108
rect 11330 18096 11336 18108
rect 11388 18096 11394 18148
rect 11808 18136 11836 18167
rect 12066 18136 12072 18148
rect 11808 18108 12072 18136
rect 12066 18096 12072 18108
rect 12124 18096 12130 18148
rect 8128 18040 10364 18068
rect 11054 18028 11060 18080
rect 11112 18028 11118 18080
rect 11514 18028 11520 18080
rect 11572 18028 11578 18080
rect 11977 18071 12035 18077
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12176 18068 12204 18235
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 12345 18275 12403 18281
rect 12345 18272 12357 18275
rect 12308 18244 12357 18272
rect 12308 18232 12314 18244
rect 12345 18241 12357 18244
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 13078 18232 13084 18284
rect 13136 18232 13142 18284
rect 13096 18204 13124 18232
rect 13188 18213 13216 18312
rect 13372 18312 14044 18340
rect 13372 18281 13400 18312
rect 14016 18284 14044 18312
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18241 13415 18275
rect 13357 18235 13415 18241
rect 13446 18232 13452 18284
rect 13504 18232 13510 18284
rect 13538 18232 13544 18284
rect 13596 18272 13602 18284
rect 13817 18275 13875 18281
rect 13817 18272 13829 18275
rect 13596 18244 13829 18272
rect 13596 18232 13602 18244
rect 13817 18241 13829 18244
rect 13863 18241 13875 18275
rect 13817 18235 13875 18241
rect 13998 18232 14004 18284
rect 14056 18232 14062 18284
rect 14108 18272 14136 18368
rect 14384 18340 14412 18368
rect 15289 18343 15347 18349
rect 15289 18340 15301 18343
rect 14384 18312 15301 18340
rect 15289 18309 15301 18312
rect 15335 18309 15347 18343
rect 15289 18303 15347 18309
rect 19429 18343 19487 18349
rect 19429 18309 19441 18343
rect 19475 18340 19487 18343
rect 19720 18340 19748 18368
rect 22066 18340 22094 18380
rect 19475 18312 19748 18340
rect 22020 18312 22094 18340
rect 22204 18312 23152 18340
rect 19475 18309 19487 18312
rect 19429 18303 19487 18309
rect 14461 18275 14519 18281
rect 14461 18272 14473 18275
rect 14108 18244 14473 18272
rect 14461 18241 14473 18244
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 15194 18232 15200 18284
rect 15252 18232 15258 18284
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 19024 18244 19165 18272
rect 19024 18232 19030 18244
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 20530 18232 20536 18284
rect 20588 18232 20594 18284
rect 12406 18176 13124 18204
rect 13173 18207 13231 18213
rect 12250 18096 12256 18148
rect 12308 18136 12314 18148
rect 12406 18136 12434 18176
rect 13173 18173 13185 18207
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18204 13323 18207
rect 13464 18204 13492 18232
rect 22020 18216 22048 18312
rect 22204 18284 22232 18312
rect 22186 18232 22192 18284
rect 22244 18232 22250 18284
rect 22738 18232 22744 18284
rect 22796 18232 22802 18284
rect 23124 18281 23152 18312
rect 23290 18300 23296 18352
rect 23348 18340 23354 18352
rect 23385 18343 23443 18349
rect 23385 18340 23397 18343
rect 23348 18312 23397 18340
rect 23348 18300 23354 18312
rect 23385 18309 23397 18312
rect 23431 18309 23443 18343
rect 23492 18340 23520 18380
rect 23492 18312 23874 18340
rect 23385 18303 23443 18309
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 13311 18176 13492 18204
rect 13633 18207 13691 18213
rect 13311 18173 13323 18176
rect 13265 18167 13323 18173
rect 13633 18173 13645 18207
rect 13679 18173 13691 18207
rect 13633 18167 13691 18173
rect 13648 18136 13676 18167
rect 22002 18164 22008 18216
rect 22060 18164 22066 18216
rect 22922 18164 22928 18216
rect 22980 18204 22986 18216
rect 23017 18207 23075 18213
rect 23017 18204 23029 18207
rect 22980 18176 23029 18204
rect 22980 18164 22986 18176
rect 23017 18173 23029 18176
rect 23063 18173 23075 18207
rect 23124 18204 23152 18235
rect 23382 18204 23388 18216
rect 23124 18176 23388 18204
rect 23017 18167 23075 18173
rect 23382 18164 23388 18176
rect 23440 18164 23446 18216
rect 25130 18164 25136 18216
rect 25188 18164 25194 18216
rect 12308 18108 12434 18136
rect 13188 18108 13676 18136
rect 12308 18096 12314 18108
rect 13188 18080 13216 18108
rect 12023 18040 12204 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 13170 18028 13176 18080
rect 13228 18028 13234 18080
rect 13538 18028 13544 18080
rect 13596 18028 13602 18080
rect 14001 18071 14059 18077
rect 14001 18037 14013 18071
rect 14047 18068 14059 18071
rect 14458 18068 14464 18080
rect 14047 18040 14464 18068
rect 14047 18037 14059 18040
rect 14001 18031 14059 18037
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 20898 18028 20904 18080
rect 20956 18028 20962 18080
rect 22554 18028 22560 18080
rect 22612 18028 22618 18080
rect 22925 18071 22983 18077
rect 22925 18037 22937 18071
rect 22971 18068 22983 18071
rect 24118 18068 24124 18080
rect 22971 18040 24124 18068
rect 22971 18037 22983 18040
rect 22925 18031 22983 18037
rect 24118 18028 24124 18040
rect 24176 18028 24182 18080
rect 1104 17978 26496 18000
rect 1104 17926 4124 17978
rect 4176 17926 4188 17978
rect 4240 17926 4252 17978
rect 4304 17926 4316 17978
rect 4368 17926 4380 17978
rect 4432 17926 10472 17978
rect 10524 17926 10536 17978
rect 10588 17926 10600 17978
rect 10652 17926 10664 17978
rect 10716 17926 10728 17978
rect 10780 17926 16820 17978
rect 16872 17926 16884 17978
rect 16936 17926 16948 17978
rect 17000 17926 17012 17978
rect 17064 17926 17076 17978
rect 17128 17926 23168 17978
rect 23220 17926 23232 17978
rect 23284 17926 23296 17978
rect 23348 17926 23360 17978
rect 23412 17926 23424 17978
rect 23476 17926 26496 17978
rect 1104 17904 26496 17926
rect 8113 17867 8171 17873
rect 8113 17833 8125 17867
rect 8159 17864 8171 17867
rect 8202 17864 8208 17876
rect 8159 17836 8208 17864
rect 8159 17833 8171 17836
rect 8113 17827 8171 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 8386 17824 8392 17876
rect 8444 17824 8450 17876
rect 8570 17824 8576 17876
rect 8628 17824 8634 17876
rect 9122 17824 9128 17876
rect 9180 17824 9186 17876
rect 11974 17864 11980 17876
rect 9876 17836 11980 17864
rect 5721 17731 5779 17737
rect 5721 17697 5733 17731
rect 5767 17728 5779 17731
rect 5994 17728 6000 17740
rect 5767 17700 6000 17728
rect 5767 17697 5779 17700
rect 5721 17691 5779 17697
rect 5994 17688 6000 17700
rect 6052 17688 6058 17740
rect 8588 17728 8616 17824
rect 9876 17796 9904 17836
rect 11974 17824 11980 17836
rect 12032 17864 12038 17876
rect 12032 17836 12204 17864
rect 12032 17824 12038 17836
rect 8404 17700 8616 17728
rect 8864 17768 9904 17796
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 8404 17669 8432 17700
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 5868 17632 6469 17660
rect 5868 17620 5874 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17629 8447 17663
rect 8389 17623 8447 17629
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 8573 17663 8631 17669
rect 8573 17660 8585 17663
rect 8536 17632 8585 17660
rect 8536 17620 8542 17632
rect 8573 17629 8585 17632
rect 8619 17660 8631 17663
rect 8864 17660 8892 17768
rect 9950 17728 9956 17740
rect 8956 17700 9956 17728
rect 8956 17669 8984 17700
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10413 17731 10471 17737
rect 10413 17697 10425 17731
rect 10459 17728 10471 17731
rect 11054 17728 11060 17740
rect 10459 17700 11060 17728
rect 10459 17697 10471 17700
rect 10413 17691 10471 17697
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 11164 17700 11560 17728
rect 8619 17632 8892 17660
rect 8941 17663 8999 17669
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 8941 17629 8953 17663
rect 8987 17629 8999 17663
rect 8941 17623 8999 17629
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 9766 17660 9772 17672
rect 9232 17632 9772 17660
rect 5445 17595 5503 17601
rect 5445 17561 5457 17595
rect 5491 17592 5503 17595
rect 5905 17595 5963 17601
rect 5905 17592 5917 17595
rect 5491 17564 5917 17592
rect 5491 17561 5503 17564
rect 5445 17555 5503 17561
rect 5905 17561 5917 17564
rect 5951 17561 5963 17595
rect 5905 17555 5963 17561
rect 4614 17484 4620 17536
rect 4672 17524 4678 17536
rect 5077 17527 5135 17533
rect 5077 17524 5089 17527
rect 4672 17496 5089 17524
rect 4672 17484 4678 17496
rect 5077 17493 5089 17496
rect 5123 17493 5135 17527
rect 5077 17487 5135 17493
rect 5537 17527 5595 17533
rect 5537 17493 5549 17527
rect 5583 17524 5595 17527
rect 6638 17524 6644 17536
rect 5583 17496 6644 17524
rect 5583 17493 5595 17496
rect 5537 17487 5595 17493
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 9232 17524 9260 17632
rect 9766 17620 9772 17632
rect 9824 17660 9830 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 9824 17632 10149 17660
rect 9824 17620 9830 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17660 11023 17663
rect 11164 17660 11192 17700
rect 11532 17672 11560 17700
rect 12176 17672 12204 17836
rect 12342 17824 12348 17876
rect 12400 17824 12406 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22189 17867 22247 17873
rect 22189 17864 22201 17867
rect 22152 17836 22201 17864
rect 22152 17824 22158 17836
rect 22189 17833 22201 17836
rect 22235 17833 22247 17867
rect 22189 17827 22247 17833
rect 22830 17824 22836 17876
rect 22888 17864 22894 17876
rect 23201 17867 23259 17873
rect 23201 17864 23213 17867
rect 22888 17836 23213 17864
rect 22888 17824 22894 17836
rect 23201 17833 23213 17836
rect 23247 17833 23259 17867
rect 24854 17864 24860 17876
rect 23201 17827 23259 17833
rect 23308 17836 24860 17864
rect 12526 17756 12532 17808
rect 12584 17756 12590 17808
rect 21082 17728 21088 17740
rect 20732 17700 21088 17728
rect 11011 17632 11192 17660
rect 11241 17663 11299 17669
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 10796 17592 10824 17623
rect 11146 17592 11152 17604
rect 9646 17564 10732 17592
rect 10796 17564 11152 17592
rect 7984 17496 9260 17524
rect 7984 17484 7990 17496
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 9646 17524 9674 17564
rect 9364 17496 9674 17524
rect 9953 17527 10011 17533
rect 9364 17484 9370 17496
rect 9953 17493 9965 17527
rect 9999 17524 10011 17527
rect 10042 17524 10048 17536
rect 9999 17496 10048 17524
rect 9999 17493 10011 17496
rect 9953 17487 10011 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 10704 17524 10732 17564
rect 11146 17552 11152 17564
rect 11204 17552 11210 17604
rect 11256 17592 11284 17623
rect 11330 17620 11336 17672
rect 11388 17620 11394 17672
rect 11514 17620 11520 17672
rect 11572 17620 11578 17672
rect 12066 17620 12072 17672
rect 12124 17620 12130 17672
rect 12158 17620 12164 17672
rect 12216 17620 12222 17672
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 15654 17660 15660 17672
rect 14608 17632 15660 17660
rect 14608 17620 14614 17632
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 18141 17663 18199 17669
rect 18141 17629 18153 17663
rect 18187 17660 18199 17663
rect 18233 17663 18291 17669
rect 18233 17660 18245 17663
rect 18187 17632 18245 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 18233 17629 18245 17632
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 18598 17660 18604 17672
rect 18463 17632 18604 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17660 18751 17663
rect 18782 17660 18788 17672
rect 18739 17632 18788 17660
rect 18739 17629 18751 17632
rect 18693 17623 18751 17629
rect 18782 17620 18788 17632
rect 18840 17620 18846 17672
rect 18874 17620 18880 17672
rect 18932 17660 18938 17672
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 18932 17632 19809 17660
rect 18932 17620 18938 17632
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 20530 17620 20536 17672
rect 20588 17660 20594 17672
rect 20732 17660 20760 17700
rect 21082 17688 21088 17700
rect 21140 17688 21146 17740
rect 22097 17731 22155 17737
rect 22097 17697 22109 17731
rect 22143 17728 22155 17731
rect 22186 17728 22192 17740
rect 22143 17700 22192 17728
rect 22143 17697 22155 17700
rect 22097 17691 22155 17697
rect 22186 17688 22192 17700
rect 22244 17688 22250 17740
rect 23308 17728 23336 17836
rect 24854 17824 24860 17836
rect 24912 17864 24918 17876
rect 24912 17836 25820 17864
rect 24912 17824 24918 17836
rect 23566 17756 23572 17808
rect 23624 17796 23630 17808
rect 23624 17768 24440 17796
rect 23624 17756 23630 17768
rect 22296 17700 23336 17728
rect 23845 17731 23903 17737
rect 20588 17646 20760 17660
rect 20588 17632 20746 17646
rect 20588 17620 20594 17632
rect 11606 17592 11612 17604
rect 11256 17564 11612 17592
rect 11606 17552 11612 17564
rect 11664 17552 11670 17604
rect 12710 17552 12716 17604
rect 12768 17552 12774 17604
rect 20073 17595 20131 17601
rect 20073 17561 20085 17595
rect 20119 17561 20131 17595
rect 20073 17555 20131 17561
rect 21821 17595 21879 17601
rect 21821 17561 21833 17595
rect 21867 17592 21879 17595
rect 22094 17592 22100 17604
rect 21867 17564 22100 17592
rect 21867 17561 21879 17564
rect 21821 17555 21879 17561
rect 11422 17524 11428 17536
rect 10704 17496 11428 17524
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 11793 17527 11851 17533
rect 11793 17493 11805 17527
rect 11839 17524 11851 17527
rect 12250 17524 12256 17536
rect 11839 17496 12256 17524
rect 11839 17493 11851 17496
rect 11793 17487 11851 17493
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 14826 17484 14832 17536
rect 14884 17484 14890 17536
rect 17218 17484 17224 17536
rect 17276 17524 17282 17536
rect 17497 17527 17555 17533
rect 17497 17524 17509 17527
rect 17276 17496 17509 17524
rect 17276 17484 17282 17496
rect 17497 17493 17509 17496
rect 17543 17493 17555 17527
rect 17497 17487 17555 17493
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 18601 17527 18659 17533
rect 18601 17524 18613 17527
rect 18472 17496 18613 17524
rect 18472 17484 18478 17496
rect 18601 17493 18613 17496
rect 18647 17493 18659 17527
rect 18601 17487 18659 17493
rect 19058 17484 19064 17536
rect 19116 17524 19122 17536
rect 19245 17527 19303 17533
rect 19245 17524 19257 17527
rect 19116 17496 19257 17524
rect 19116 17484 19122 17496
rect 19245 17493 19257 17496
rect 19291 17493 19303 17527
rect 20088 17524 20116 17555
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 22296 17592 22324 17700
rect 23845 17697 23857 17731
rect 23891 17697 23903 17731
rect 23845 17691 23903 17697
rect 22370 17620 22376 17672
rect 22428 17660 22434 17672
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 22428 17632 22753 17660
rect 22428 17620 22434 17632
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 22922 17620 22928 17672
rect 22980 17620 22986 17672
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17660 23167 17663
rect 23860 17660 23888 17691
rect 24118 17688 24124 17740
rect 24176 17688 24182 17740
rect 24412 17737 24440 17768
rect 24397 17731 24455 17737
rect 24397 17697 24409 17731
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 23155 17632 23888 17660
rect 24136 17660 24164 17688
rect 24213 17663 24271 17669
rect 24213 17660 24225 17663
rect 24136 17632 24225 17660
rect 23155 17629 23167 17632
rect 23109 17623 23167 17629
rect 22204 17564 22324 17592
rect 20990 17524 20996 17536
rect 20088 17496 20996 17524
rect 19245 17487 19303 17493
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 22204 17524 22232 17564
rect 22830 17552 22836 17604
rect 22888 17592 22894 17604
rect 23124 17592 23152 17623
rect 23860 17592 23888 17632
rect 24213 17629 24225 17632
rect 24259 17629 24271 17663
rect 25792 17646 25820 17836
rect 24213 17623 24271 17629
rect 24673 17595 24731 17601
rect 22888 17564 23152 17592
rect 23584 17564 23796 17592
rect 23860 17564 24256 17592
rect 22888 17552 22894 17564
rect 21140 17496 22232 17524
rect 21140 17484 21146 17496
rect 22278 17484 22284 17536
rect 22336 17524 22342 17536
rect 22925 17527 22983 17533
rect 22925 17524 22937 17527
rect 22336 17496 22937 17524
rect 22336 17484 22342 17496
rect 22925 17493 22937 17496
rect 22971 17524 22983 17527
rect 23014 17524 23020 17536
rect 22971 17496 23020 17524
rect 22971 17493 22983 17496
rect 22925 17487 22983 17493
rect 23014 17484 23020 17496
rect 23072 17484 23078 17536
rect 23584 17533 23612 17564
rect 23768 17536 23796 17564
rect 23569 17527 23627 17533
rect 23569 17493 23581 17527
rect 23615 17493 23627 17527
rect 23569 17487 23627 17493
rect 23658 17484 23664 17536
rect 23716 17484 23722 17536
rect 23750 17484 23756 17536
rect 23808 17484 23814 17536
rect 24026 17484 24032 17536
rect 24084 17524 24090 17536
rect 24121 17527 24179 17533
rect 24121 17524 24133 17527
rect 24084 17496 24133 17524
rect 24084 17484 24090 17496
rect 24121 17493 24133 17496
rect 24167 17493 24179 17527
rect 24228 17524 24256 17564
rect 24673 17561 24685 17595
rect 24719 17592 24731 17595
rect 24946 17592 24952 17604
rect 24719 17564 24952 17592
rect 24719 17561 24731 17564
rect 24673 17555 24731 17561
rect 24946 17552 24952 17564
rect 25004 17552 25010 17604
rect 25038 17524 25044 17536
rect 24228 17496 25044 17524
rect 24121 17487 24179 17493
rect 25038 17484 25044 17496
rect 25096 17484 25102 17536
rect 26142 17484 26148 17536
rect 26200 17484 26206 17536
rect 1104 17434 26656 17456
rect 1104 17382 7298 17434
rect 7350 17382 7362 17434
rect 7414 17382 7426 17434
rect 7478 17382 7490 17434
rect 7542 17382 7554 17434
rect 7606 17382 13646 17434
rect 13698 17382 13710 17434
rect 13762 17382 13774 17434
rect 13826 17382 13838 17434
rect 13890 17382 13902 17434
rect 13954 17382 19994 17434
rect 20046 17382 20058 17434
rect 20110 17382 20122 17434
rect 20174 17382 20186 17434
rect 20238 17382 20250 17434
rect 20302 17382 26342 17434
rect 26394 17382 26406 17434
rect 26458 17382 26470 17434
rect 26522 17382 26534 17434
rect 26586 17382 26598 17434
rect 26650 17382 26656 17434
rect 1104 17360 26656 17382
rect 11606 17280 11612 17332
rect 11664 17280 11670 17332
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12710 17320 12716 17332
rect 12483 17292 12716 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 13725 17323 13783 17329
rect 13725 17289 13737 17323
rect 13771 17320 13783 17323
rect 14550 17320 14556 17332
rect 13771 17292 14556 17320
rect 13771 17289 13783 17292
rect 13725 17283 13783 17289
rect 14550 17280 14556 17292
rect 14608 17280 14614 17332
rect 17218 17280 17224 17332
rect 17276 17280 17282 17332
rect 18414 17280 18420 17332
rect 18472 17280 18478 17332
rect 18874 17280 18880 17332
rect 18932 17280 18938 17332
rect 19058 17280 19064 17332
rect 19116 17320 19122 17332
rect 19116 17292 19380 17320
rect 19116 17280 19122 17292
rect 14274 17252 14280 17264
rect 12176 17224 13032 17252
rect 3970 17184 3976 17196
rect 3818 17156 3976 17184
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17184 6239 17187
rect 6270 17184 6276 17196
rect 6227 17156 6276 17184
rect 6227 17153 6239 17156
rect 6181 17147 6239 17153
rect 6270 17144 6276 17156
rect 6328 17184 6334 17196
rect 9858 17184 9864 17196
rect 6328 17156 9864 17184
rect 6328 17144 6334 17156
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 12176 17193 12204 17224
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 2406 17076 2412 17128
rect 2464 17076 2470 17128
rect 2685 17119 2743 17125
rect 2685 17085 2697 17119
rect 2731 17116 2743 17119
rect 3234 17116 3240 17128
rect 2731 17088 3240 17116
rect 2731 17085 2743 17088
rect 2685 17079 2743 17085
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17116 4215 17119
rect 4890 17116 4896 17128
rect 4203 17088 4896 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17116 5503 17119
rect 5534 17116 5540 17128
rect 5491 17088 5540 17116
rect 5491 17085 5503 17088
rect 5445 17079 5503 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 6454 17076 6460 17128
rect 6512 17076 6518 17128
rect 10226 17076 10232 17128
rect 10284 17116 10290 17128
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 10284 17088 10609 17116
rect 10284 17076 10290 17088
rect 10597 17085 10609 17088
rect 10643 17116 10655 17119
rect 10962 17116 10968 17128
rect 10643 17088 10968 17116
rect 10643 17085 10655 17088
rect 10597 17079 10655 17085
rect 10962 17076 10968 17088
rect 11020 17116 11026 17128
rect 11532 17116 11560 17147
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 12544 17193 12572 17224
rect 13004 17196 13032 17224
rect 13924 17224 14136 17252
rect 12529 17187 12587 17193
rect 12529 17153 12541 17187
rect 12575 17184 12587 17187
rect 12713 17187 12771 17193
rect 12575 17156 12609 17184
rect 12575 17153 12587 17156
rect 12529 17147 12587 17153
rect 12713 17153 12725 17187
rect 12759 17184 12771 17187
rect 12894 17184 12900 17196
rect 12759 17156 12900 17184
rect 12759 17153 12771 17156
rect 12713 17147 12771 17153
rect 11020 17088 11560 17116
rect 12268 17116 12296 17144
rect 12728 17116 12756 17147
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 12986 17144 12992 17196
rect 13044 17144 13050 17196
rect 13924 17193 13952 17224
rect 13909 17187 13967 17193
rect 13909 17153 13921 17187
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 14016 17116 14044 17147
rect 12268 17088 14044 17116
rect 14108 17116 14136 17224
rect 14200 17224 14280 17252
rect 14200 17193 14228 17224
rect 14274 17212 14280 17224
rect 14332 17252 14338 17264
rect 16301 17255 16359 17261
rect 16301 17252 16313 17255
rect 14332 17224 16313 17252
rect 14332 17212 14338 17224
rect 16301 17221 16313 17224
rect 16347 17221 16359 17255
rect 16301 17215 16359 17221
rect 16945 17255 17003 17261
rect 16945 17221 16957 17255
rect 16991 17252 17003 17255
rect 17236 17252 17264 17280
rect 16991 17224 17264 17252
rect 19245 17255 19303 17261
rect 16991 17221 17003 17224
rect 16945 17215 17003 17221
rect 19245 17221 19257 17255
rect 19291 17252 19303 17255
rect 19352 17252 19380 17292
rect 20714 17280 20720 17332
rect 20772 17280 20778 17332
rect 21913 17323 21971 17329
rect 21913 17289 21925 17323
rect 21959 17320 21971 17323
rect 22278 17320 22284 17332
rect 21959 17292 22284 17320
rect 21959 17289 21971 17292
rect 21913 17283 21971 17289
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 22741 17323 22799 17329
rect 22741 17289 22753 17323
rect 22787 17320 22799 17323
rect 22830 17320 22836 17332
rect 22787 17292 22836 17320
rect 22787 17289 22799 17292
rect 22741 17283 22799 17289
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 24210 17280 24216 17332
rect 24268 17320 24274 17332
rect 25038 17320 25044 17332
rect 24268 17292 25044 17320
rect 24268 17280 24274 17292
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 20530 17252 20536 17264
rect 19291 17224 19380 17252
rect 20470 17224 20536 17252
rect 19291 17221 19303 17224
rect 19245 17215 19303 17221
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 22462 17218 22468 17264
rect 22388 17212 22468 17218
rect 22520 17212 22526 17264
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 15194 17144 15200 17196
rect 15252 17144 15258 17196
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17184 16175 17187
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 16163 17156 16221 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 18601 17187 18659 17193
rect 16209 17147 16267 17153
rect 14108 17088 14688 17116
rect 11020 17076 11026 17088
rect 12158 17008 12164 17060
rect 12216 17048 12222 17060
rect 12621 17051 12679 17057
rect 12621 17048 12633 17051
rect 12216 17020 12633 17048
rect 12216 17008 12222 17020
rect 12621 17017 12633 17020
rect 12667 17017 12679 17051
rect 12621 17011 12679 17017
rect 14001 17051 14059 17057
rect 14001 17017 14013 17051
rect 14047 17048 14059 17051
rect 14550 17048 14556 17060
rect 14047 17020 14556 17048
rect 14047 17017 14059 17020
rect 14001 17011 14059 17017
rect 14550 17008 14556 17020
rect 14608 17008 14614 17060
rect 4249 16983 4307 16989
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 4522 16980 4528 16992
rect 4295 16952 4528 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 4522 16940 4528 16952
rect 4580 16940 4586 16992
rect 7101 16983 7159 16989
rect 7101 16949 7113 16983
rect 7147 16980 7159 16983
rect 7558 16980 7564 16992
rect 7147 16952 7564 16980
rect 7147 16949 7159 16952
rect 7101 16943 7159 16949
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 11241 16983 11299 16989
rect 11241 16949 11253 16983
rect 11287 16980 11299 16983
rect 11422 16980 11428 16992
rect 11287 16952 11428 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 14366 16940 14372 16992
rect 14424 16940 14430 16992
rect 14660 16980 14688 17088
rect 15010 17076 15016 17128
rect 15068 17076 15074 17128
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 15473 17119 15531 17125
rect 15473 17116 15485 17119
rect 15344 17088 15485 17116
rect 15344 17076 15350 17088
rect 15473 17085 15485 17088
rect 15519 17085 15531 17119
rect 15473 17079 15531 17085
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 16669 17119 16727 17125
rect 16669 17116 16681 17119
rect 16632 17088 16681 17116
rect 16632 17076 16638 17088
rect 16669 17085 16681 17088
rect 16715 17085 16727 17119
rect 18064 17116 18092 17170
rect 18601 17153 18613 17187
rect 18647 17184 18659 17187
rect 18690 17184 18696 17196
rect 18647 17156 18696 17184
rect 18647 17153 18659 17156
rect 18601 17147 18659 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 20898 17144 20904 17196
rect 20956 17184 20962 17196
rect 21361 17187 21419 17193
rect 21361 17184 21373 17187
rect 20956 17156 21373 17184
rect 20956 17144 20962 17156
rect 21361 17153 21373 17156
rect 21407 17153 21419 17187
rect 21361 17147 21419 17153
rect 22094 17144 22100 17196
rect 22152 17144 22158 17196
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 16669 17079 16727 17085
rect 16776 17088 18092 17116
rect 14826 17008 14832 17060
rect 14884 17048 14890 17060
rect 16776 17048 16804 17088
rect 18874 17076 18880 17128
rect 18932 17076 18938 17128
rect 18966 17076 18972 17128
rect 19024 17076 19030 17128
rect 19242 17076 19248 17128
rect 19300 17116 19306 17128
rect 20622 17116 20628 17128
rect 19300 17088 20628 17116
rect 19300 17076 19306 17088
rect 20622 17076 20628 17088
rect 20680 17116 20686 17128
rect 21174 17116 21180 17128
rect 20680 17088 21180 17116
rect 20680 17076 20686 17088
rect 21174 17076 21180 17088
rect 21232 17116 21238 17128
rect 22002 17116 22008 17128
rect 21232 17088 22008 17116
rect 21232 17076 21238 17088
rect 22002 17076 22008 17088
rect 22060 17076 22066 17128
rect 14884 17020 16804 17048
rect 22204 17048 22232 17147
rect 22278 17144 22284 17196
rect 22336 17144 22342 17196
rect 22388 17190 22508 17212
rect 22388 17187 22457 17190
rect 22388 17156 22411 17187
rect 22399 17153 22411 17156
rect 22445 17153 22457 17187
rect 22399 17147 22457 17153
rect 22646 17144 22652 17196
rect 22704 17144 22710 17196
rect 23290 17144 23296 17196
rect 23348 17144 23354 17196
rect 24854 17184 24860 17196
rect 24702 17156 24860 17184
rect 24854 17144 24860 17156
rect 24912 17144 24918 17196
rect 25314 17144 25320 17196
rect 25372 17184 25378 17196
rect 25409 17187 25467 17193
rect 25409 17184 25421 17187
rect 25372 17156 25421 17184
rect 25372 17144 25378 17156
rect 25409 17153 25421 17156
rect 25455 17184 25467 17187
rect 26142 17184 26148 17196
rect 25455 17156 26148 17184
rect 25455 17153 25467 17156
rect 25409 17147 25467 17153
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 22557 17119 22615 17125
rect 22557 17085 22569 17119
rect 22603 17116 22615 17119
rect 22738 17116 22744 17128
rect 22603 17088 22744 17116
rect 22603 17085 22615 17088
rect 22557 17079 22615 17085
rect 22738 17076 22744 17088
rect 22796 17116 22802 17128
rect 22922 17116 22928 17128
rect 22796 17088 22928 17116
rect 22796 17076 22802 17088
rect 22922 17076 22928 17088
rect 22980 17076 22986 17128
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17085 23167 17119
rect 23109 17079 23167 17085
rect 22646 17048 22652 17060
rect 22204 17020 22652 17048
rect 14884 17008 14890 17020
rect 22646 17008 22652 17020
rect 22704 17008 22710 17060
rect 23124 17048 23152 17079
rect 23566 17076 23572 17128
rect 23624 17076 23630 17128
rect 22848 17020 23152 17048
rect 15289 16983 15347 16989
rect 15289 16980 15301 16983
rect 14660 16952 15301 16980
rect 15289 16949 15301 16952
rect 15335 16980 15347 16983
rect 15746 16980 15752 16992
rect 15335 16952 15752 16980
rect 15335 16949 15347 16952
rect 15289 16943 15347 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 18690 16940 18696 16992
rect 18748 16940 18754 16992
rect 18874 16940 18880 16992
rect 18932 16980 18938 16992
rect 19334 16980 19340 16992
rect 18932 16952 19340 16980
rect 18932 16940 18938 16952
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 20806 16940 20812 16992
rect 20864 16940 20870 16992
rect 22370 16940 22376 16992
rect 22428 16980 22434 16992
rect 22848 16980 22876 17020
rect 22428 16952 22876 16980
rect 22428 16940 22434 16952
rect 22922 16940 22928 16992
rect 22980 16940 22986 16992
rect 23124 16980 23152 17020
rect 24210 16980 24216 16992
rect 23124 16952 24216 16980
rect 24210 16940 24216 16952
rect 24268 16940 24274 16992
rect 25958 16940 25964 16992
rect 26016 16940 26022 16992
rect 1104 16890 26496 16912
rect 1104 16838 4124 16890
rect 4176 16838 4188 16890
rect 4240 16838 4252 16890
rect 4304 16838 4316 16890
rect 4368 16838 4380 16890
rect 4432 16838 10472 16890
rect 10524 16838 10536 16890
rect 10588 16838 10600 16890
rect 10652 16838 10664 16890
rect 10716 16838 10728 16890
rect 10780 16838 16820 16890
rect 16872 16838 16884 16890
rect 16936 16838 16948 16890
rect 17000 16838 17012 16890
rect 17064 16838 17076 16890
rect 17128 16838 23168 16890
rect 23220 16838 23232 16890
rect 23284 16838 23296 16890
rect 23348 16838 23360 16890
rect 23412 16838 23424 16890
rect 23476 16838 26496 16890
rect 1104 16816 26496 16838
rect 2406 16736 2412 16788
rect 2464 16776 2470 16788
rect 2464 16748 2774 16776
rect 2464 16736 2470 16748
rect 2746 16640 2774 16748
rect 3234 16736 3240 16788
rect 3292 16736 3298 16788
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 8033 16779 8091 16785
rect 8033 16776 8045 16779
rect 7616 16748 8045 16776
rect 7616 16736 7622 16748
rect 8033 16745 8045 16748
rect 8079 16745 8091 16779
rect 8033 16739 8091 16745
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 11480 16748 12296 16776
rect 11480 16736 11486 16748
rect 12066 16668 12072 16720
rect 12124 16708 12130 16720
rect 12161 16711 12219 16717
rect 12161 16708 12173 16711
rect 12124 16680 12173 16708
rect 12124 16668 12130 16680
rect 12161 16677 12173 16680
rect 12207 16677 12219 16711
rect 12161 16671 12219 16677
rect 4709 16643 4767 16649
rect 4709 16640 4721 16643
rect 2746 16612 4721 16640
rect 4709 16609 4721 16612
rect 4755 16640 4767 16643
rect 6362 16640 6368 16652
rect 4755 16612 6368 16640
rect 4755 16609 4767 16612
rect 4709 16603 4767 16609
rect 6362 16600 6368 16612
rect 6420 16640 6426 16652
rect 7006 16640 7012 16652
rect 6420 16612 7012 16640
rect 6420 16600 6426 16612
rect 7006 16600 7012 16612
rect 7064 16640 7070 16652
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 7064 16612 8309 16640
rect 7064 16600 7070 16612
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 9585 16643 9643 16649
rect 9585 16609 9597 16643
rect 9631 16640 9643 16643
rect 10318 16640 10324 16652
rect 9631 16612 10324 16640
rect 9631 16609 9643 16612
rect 9585 16603 9643 16609
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16640 10471 16643
rect 11238 16640 11244 16652
rect 10459 16612 11244 16640
rect 10459 16609 10471 16612
rect 10413 16603 10471 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 12268 16649 12296 16748
rect 14366 16736 14372 16788
rect 14424 16736 14430 16788
rect 14550 16736 14556 16788
rect 14608 16736 14614 16788
rect 16472 16779 16530 16785
rect 16472 16745 16484 16779
rect 16518 16776 16530 16779
rect 18877 16779 18935 16785
rect 18877 16776 18889 16779
rect 16518 16748 18889 16776
rect 16518 16745 16530 16748
rect 16472 16739 16530 16745
rect 18877 16745 18889 16748
rect 18923 16745 18935 16779
rect 18877 16739 18935 16745
rect 20349 16779 20407 16785
rect 20349 16745 20361 16779
rect 20395 16776 20407 16779
rect 20438 16776 20444 16788
rect 20395 16748 20444 16776
rect 20395 16745 20407 16748
rect 20349 16739 20407 16745
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 20714 16736 20720 16788
rect 20772 16776 20778 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 20772 16748 21281 16776
rect 20772 16736 20778 16748
rect 21269 16745 21281 16748
rect 21315 16745 21327 16779
rect 21269 16739 21327 16745
rect 21634 16736 21640 16788
rect 21692 16736 21698 16788
rect 23109 16779 23167 16785
rect 23109 16745 23121 16779
rect 23155 16776 23167 16779
rect 23566 16776 23572 16788
rect 23155 16748 23572 16776
rect 23155 16745 23167 16748
rect 23109 16739 23167 16745
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 24213 16779 24271 16785
rect 24213 16745 24225 16779
rect 24259 16745 24271 16779
rect 24213 16739 24271 16745
rect 14384 16708 14412 16736
rect 13004 16680 14412 16708
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 3973 16575 4031 16581
rect 3973 16572 3985 16575
rect 3467 16544 3985 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 3973 16541 3985 16544
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 4430 16532 4436 16584
rect 4488 16532 4494 16584
rect 4522 16532 4528 16584
rect 4580 16532 4586 16584
rect 6914 16572 6920 16584
rect 6118 16544 6920 16572
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 4157 16507 4215 16513
rect 4157 16473 4169 16507
rect 4203 16473 4215 16507
rect 4157 16467 4215 16473
rect 4172 16436 4200 16467
rect 4246 16464 4252 16516
rect 4304 16504 4310 16516
rect 4341 16507 4399 16513
rect 4341 16504 4353 16507
rect 4304 16476 4353 16504
rect 4304 16464 4310 16476
rect 4341 16473 4353 16476
rect 4387 16473 4399 16507
rect 4341 16467 4399 16473
rect 4540 16436 4568 16532
rect 4985 16507 5043 16513
rect 4985 16504 4997 16507
rect 4632 16476 4997 16504
rect 4632 16445 4660 16476
rect 4985 16473 4997 16476
rect 5031 16473 5043 16507
rect 4985 16467 5043 16473
rect 6362 16464 6368 16516
rect 6420 16504 6426 16516
rect 10689 16507 10747 16513
rect 6420 16476 6592 16504
rect 6420 16464 6426 16476
rect 4172 16408 4568 16436
rect 4617 16439 4675 16445
rect 4617 16405 4629 16439
rect 4663 16405 4675 16439
rect 4617 16399 4675 16405
rect 5994 16396 6000 16448
rect 6052 16436 6058 16448
rect 6564 16445 6592 16476
rect 10689 16473 10701 16507
rect 10735 16504 10747 16507
rect 10778 16504 10784 16516
rect 10735 16476 10784 16504
rect 10735 16473 10747 16476
rect 10689 16467 10747 16473
rect 10778 16464 10784 16476
rect 10836 16464 10842 16516
rect 10888 16476 11178 16504
rect 6457 16439 6515 16445
rect 6457 16436 6469 16439
rect 6052 16408 6469 16436
rect 6052 16396 6058 16408
rect 6457 16405 6469 16408
rect 6503 16405 6515 16439
rect 6457 16399 6515 16405
rect 6549 16439 6607 16445
rect 6549 16405 6561 16439
rect 6595 16405 6607 16439
rect 6549 16399 6607 16405
rect 8938 16396 8944 16448
rect 8996 16396 9002 16448
rect 10134 16396 10140 16448
rect 10192 16436 10198 16448
rect 10888 16436 10916 16476
rect 10192 16408 10916 16436
rect 10192 16396 10198 16408
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 12347 16436 12375 16535
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 13004 16581 13032 16680
rect 13909 16643 13967 16649
rect 13909 16609 13921 16643
rect 13955 16640 13967 16643
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13955 16612 14105 16640
rect 13955 16609 13967 16612
rect 13909 16603 13967 16609
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14568 16640 14596 16736
rect 18598 16668 18604 16720
rect 18656 16708 18662 16720
rect 18785 16711 18843 16717
rect 18785 16708 18797 16711
rect 18656 16680 18797 16708
rect 18656 16668 18662 16680
rect 18785 16677 18797 16680
rect 18831 16677 18843 16711
rect 18785 16671 18843 16677
rect 18984 16680 19932 16708
rect 15565 16643 15623 16649
rect 15565 16640 15577 16643
rect 14568 16612 15577 16640
rect 14093 16603 14151 16609
rect 15565 16609 15577 16612
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 15841 16643 15899 16649
rect 15841 16609 15853 16643
rect 15887 16640 15899 16643
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 15887 16612 16221 16640
rect 15887 16609 15899 16612
rect 15841 16603 15899 16609
rect 16209 16609 16221 16612
rect 16255 16640 16267 16643
rect 16574 16640 16580 16652
rect 16255 16612 16580 16640
rect 16255 16609 16267 16612
rect 16209 16603 16267 16609
rect 12897 16575 12955 16581
rect 12897 16572 12909 16575
rect 12584 16544 12909 16572
rect 12584 16532 12590 16544
rect 12897 16541 12909 16544
rect 12943 16541 12955 16575
rect 12897 16535 12955 16541
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16541 13047 16575
rect 12989 16535 13047 16541
rect 13556 16476 14320 16504
rect 13556 16448 13584 16476
rect 12618 16436 12624 16448
rect 11020 16408 12624 16436
rect 11020 16396 11026 16408
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 12710 16396 12716 16448
rect 12768 16396 12774 16448
rect 13262 16396 13268 16448
rect 13320 16396 13326 16448
rect 13538 16396 13544 16448
rect 13596 16396 13602 16448
rect 14292 16436 14320 16476
rect 14826 16464 14832 16516
rect 14884 16464 14890 16516
rect 15856 16504 15884 16603
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 17957 16643 18015 16649
rect 17957 16609 17969 16643
rect 18003 16640 18015 16643
rect 18141 16643 18199 16649
rect 18141 16640 18153 16643
rect 18003 16612 18153 16640
rect 18003 16609 18015 16612
rect 17957 16603 18015 16609
rect 18141 16609 18153 16612
rect 18187 16609 18199 16643
rect 18141 16603 18199 16609
rect 18690 16600 18696 16652
rect 18748 16640 18754 16652
rect 18984 16640 19012 16680
rect 19334 16640 19340 16652
rect 18748 16612 19012 16640
rect 19076 16612 19340 16640
rect 18748 16600 18754 16612
rect 18322 16532 18328 16584
rect 18380 16572 18386 16584
rect 18782 16572 18788 16584
rect 18380 16544 18788 16572
rect 18380 16532 18386 16544
rect 18782 16532 18788 16544
rect 18840 16572 18846 16584
rect 19076 16581 19104 16612
rect 19334 16600 19340 16612
rect 19392 16640 19398 16652
rect 19392 16612 19840 16640
rect 19392 16600 19398 16612
rect 19812 16584 19840 16612
rect 19904 16584 19932 16680
rect 20806 16668 20812 16720
rect 20864 16668 20870 16720
rect 21085 16711 21143 16717
rect 21085 16677 21097 16711
rect 21131 16677 21143 16711
rect 21085 16671 21143 16677
rect 20824 16640 20852 16668
rect 20732 16612 20852 16640
rect 21100 16640 21128 16671
rect 21542 16668 21548 16720
rect 21600 16708 21606 16720
rect 21821 16711 21879 16717
rect 21821 16708 21833 16711
rect 21600 16680 21833 16708
rect 21600 16668 21606 16680
rect 21821 16677 21833 16680
rect 21867 16677 21879 16711
rect 21821 16671 21879 16677
rect 22097 16711 22155 16717
rect 22097 16677 22109 16711
rect 22143 16708 22155 16711
rect 22922 16708 22928 16720
rect 22143 16680 22928 16708
rect 22143 16677 22155 16680
rect 22097 16671 22155 16677
rect 22922 16668 22928 16680
rect 22980 16668 22986 16720
rect 24228 16708 24256 16739
rect 24946 16736 24952 16788
rect 25004 16776 25010 16788
rect 25133 16779 25191 16785
rect 25133 16776 25145 16779
rect 25004 16748 25145 16776
rect 25004 16736 25010 16748
rect 25133 16745 25145 16748
rect 25179 16745 25191 16779
rect 25133 16739 25191 16745
rect 25498 16708 25504 16720
rect 23492 16680 24256 16708
rect 24826 16680 25504 16708
rect 21726 16640 21732 16652
rect 21100 16612 21732 16640
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 18840 16544 18889 16572
rect 18840 16532 18846 16544
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 19061 16575 19119 16581
rect 19061 16541 19073 16575
rect 19107 16541 19119 16575
rect 19061 16535 19119 16541
rect 19242 16532 19248 16584
rect 19300 16532 19306 16584
rect 19794 16532 19800 16584
rect 19852 16532 19858 16584
rect 19886 16532 19892 16584
rect 19944 16572 19950 16584
rect 19981 16575 20039 16581
rect 19981 16572 19993 16575
rect 19944 16544 19993 16572
rect 19944 16532 19950 16544
rect 19981 16541 19993 16544
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 20165 16575 20223 16581
rect 20165 16541 20177 16575
rect 20211 16572 20223 16575
rect 20732 16572 20760 16612
rect 21726 16600 21732 16612
rect 21784 16600 21790 16652
rect 21910 16600 21916 16652
rect 21968 16640 21974 16652
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 21968 16612 22201 16640
rect 21968 16600 21974 16612
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 22189 16603 22247 16609
rect 22317 16643 22375 16649
rect 22317 16609 22329 16643
rect 22363 16640 22375 16643
rect 22554 16640 22560 16652
rect 22363 16612 22560 16640
rect 22363 16609 22375 16612
rect 22317 16603 22375 16609
rect 22554 16600 22560 16612
rect 22612 16600 22618 16652
rect 22646 16600 22652 16652
rect 22704 16600 22710 16652
rect 22830 16600 22836 16652
rect 22888 16600 22894 16652
rect 20211 16544 20760 16572
rect 20809 16575 20867 16581
rect 20211 16541 20223 16544
rect 20165 16535 20223 16541
rect 20809 16541 20821 16575
rect 20855 16572 20867 16575
rect 20898 16572 20904 16584
rect 20855 16544 20904 16572
rect 20855 16541 20867 16544
rect 20809 16535 20867 16541
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 20990 16532 20996 16584
rect 21048 16572 21054 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 21048 16544 21097 16572
rect 21048 16532 21054 16544
rect 21085 16541 21097 16544
rect 21131 16572 21143 16575
rect 21177 16575 21235 16581
rect 21177 16572 21189 16575
rect 21131 16544 21189 16572
rect 21131 16541 21143 16544
rect 21085 16535 21143 16541
rect 21177 16541 21189 16544
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 15764 16476 15884 16504
rect 15764 16436 15792 16476
rect 17494 16464 17500 16516
rect 17552 16464 17558 16516
rect 21192 16504 21220 16535
rect 22002 16532 22008 16584
rect 22060 16532 22066 16584
rect 22465 16575 22523 16581
rect 22465 16572 22477 16575
rect 22388 16544 22477 16572
rect 22388 16516 22416 16544
rect 22465 16541 22477 16544
rect 22511 16541 22523 16575
rect 22848 16572 22876 16600
rect 23017 16575 23075 16581
rect 23017 16572 23029 16575
rect 22848 16544 23029 16572
rect 22465 16535 22523 16541
rect 23017 16541 23029 16544
rect 23063 16541 23075 16575
rect 23017 16535 23075 16541
rect 23293 16575 23351 16581
rect 23293 16541 23305 16575
rect 23339 16572 23351 16575
rect 23492 16572 23520 16680
rect 23934 16600 23940 16652
rect 23992 16640 23998 16652
rect 24826 16640 24854 16680
rect 25498 16668 25504 16680
rect 25556 16668 25562 16720
rect 23992 16612 24854 16640
rect 23992 16600 23998 16612
rect 25038 16600 25044 16652
rect 25096 16600 25102 16652
rect 25777 16643 25835 16649
rect 25777 16609 25789 16643
rect 25823 16640 25835 16643
rect 25958 16640 25964 16652
rect 25823 16612 25964 16640
rect 25823 16609 25835 16612
rect 25777 16603 25835 16609
rect 25958 16600 25964 16612
rect 26016 16600 26022 16652
rect 23339 16544 23520 16572
rect 23753 16575 23811 16581
rect 23339 16541 23351 16544
rect 23293 16535 23351 16541
rect 23753 16541 23765 16575
rect 23799 16574 23811 16575
rect 24397 16575 24455 16581
rect 23799 16572 23888 16574
rect 24397 16572 24409 16575
rect 23799 16546 24409 16572
rect 23799 16541 23811 16546
rect 23860 16544 24409 16546
rect 23753 16535 23811 16541
rect 24397 16541 24409 16544
rect 24443 16541 24455 16575
rect 24397 16535 24455 16541
rect 25317 16575 25375 16581
rect 25317 16541 25329 16575
rect 25363 16572 25375 16575
rect 25363 16544 25820 16572
rect 25363 16541 25375 16544
rect 25317 16535 25375 16541
rect 21192 16476 21772 16504
rect 14292 16408 15792 16436
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 19889 16439 19947 16445
rect 19889 16436 19901 16439
rect 19576 16408 19901 16436
rect 19576 16396 19582 16408
rect 19889 16405 19901 16408
rect 19935 16405 19947 16439
rect 19889 16399 19947 16405
rect 20898 16396 20904 16448
rect 20956 16396 20962 16448
rect 21744 16436 21772 16476
rect 22370 16464 22376 16516
rect 22428 16464 22434 16516
rect 22738 16464 22744 16516
rect 22796 16504 22802 16516
rect 22833 16507 22891 16513
rect 22833 16504 22845 16507
rect 22796 16476 22845 16504
rect 22796 16464 22802 16476
rect 22833 16473 22845 16476
rect 22879 16504 22891 16507
rect 22922 16504 22928 16516
rect 22879 16476 22928 16504
rect 22879 16473 22891 16476
rect 22833 16467 22891 16473
rect 22922 16464 22928 16476
rect 22980 16464 22986 16516
rect 23382 16464 23388 16516
rect 23440 16464 23446 16516
rect 23474 16464 23480 16516
rect 23532 16464 23538 16516
rect 23566 16464 23572 16516
rect 23624 16513 23630 16516
rect 23624 16507 23653 16513
rect 23641 16473 23653 16507
rect 23624 16467 23653 16473
rect 23845 16507 23903 16513
rect 23845 16473 23857 16507
rect 23891 16473 23903 16507
rect 23845 16467 23903 16473
rect 23624 16464 23630 16467
rect 22756 16436 22784 16464
rect 21744 16408 22784 16436
rect 23106 16396 23112 16448
rect 23164 16436 23170 16448
rect 23860 16436 23888 16467
rect 24026 16464 24032 16516
rect 24084 16464 24090 16516
rect 25406 16464 25412 16516
rect 25464 16464 25470 16516
rect 25498 16464 25504 16516
rect 25556 16504 25562 16516
rect 25682 16513 25688 16516
rect 25639 16507 25688 16513
rect 25556 16476 25601 16504
rect 25556 16464 25562 16476
rect 25639 16473 25651 16507
rect 25685 16473 25688 16507
rect 25639 16467 25688 16473
rect 25682 16464 25688 16467
rect 25740 16464 25746 16516
rect 25792 16504 25820 16544
rect 25866 16532 25872 16584
rect 25924 16532 25930 16584
rect 25961 16507 26019 16513
rect 25961 16504 25973 16507
rect 25792 16476 25973 16504
rect 25961 16473 25973 16476
rect 26007 16473 26019 16507
rect 25961 16467 26019 16473
rect 23164 16408 23888 16436
rect 23164 16396 23170 16408
rect 1104 16346 26656 16368
rect 1104 16294 7298 16346
rect 7350 16294 7362 16346
rect 7414 16294 7426 16346
rect 7478 16294 7490 16346
rect 7542 16294 7554 16346
rect 7606 16294 13646 16346
rect 13698 16294 13710 16346
rect 13762 16294 13774 16346
rect 13826 16294 13838 16346
rect 13890 16294 13902 16346
rect 13954 16294 19994 16346
rect 20046 16294 20058 16346
rect 20110 16294 20122 16346
rect 20174 16294 20186 16346
rect 20238 16294 20250 16346
rect 20302 16294 26342 16346
rect 26394 16294 26406 16346
rect 26458 16294 26470 16346
rect 26522 16294 26534 16346
rect 26586 16294 26598 16346
rect 26650 16294 26656 16346
rect 1104 16272 26656 16294
rect 3970 16192 3976 16244
rect 4028 16232 4034 16244
rect 5629 16235 5687 16241
rect 4028 16204 5488 16232
rect 4028 16192 4034 16204
rect 3142 16164 3148 16176
rect 3082 16136 3148 16164
rect 3142 16124 3148 16136
rect 3200 16164 3206 16176
rect 3988 16164 4016 16192
rect 5460 16164 5488 16204
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 5810 16232 5816 16244
rect 5675 16204 5816 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 5997 16235 6055 16241
rect 5997 16201 6009 16235
rect 6043 16232 6055 16235
rect 6454 16232 6460 16244
rect 6043 16204 6460 16232
rect 6043 16201 6055 16204
rect 5997 16195 6055 16201
rect 6454 16192 6460 16204
rect 6512 16192 6518 16244
rect 8938 16232 8944 16244
rect 7944 16204 8944 16232
rect 3200 16136 4016 16164
rect 5382 16136 5856 16164
rect 3200 16124 3206 16136
rect 5718 16056 5724 16108
rect 5776 16056 5782 16108
rect 5828 16096 5856 16136
rect 6270 16124 6276 16176
rect 6328 16164 6334 16176
rect 6365 16167 6423 16173
rect 6365 16164 6377 16167
rect 6328 16136 6377 16164
rect 6328 16124 6334 16136
rect 6365 16133 6377 16136
rect 6411 16133 6423 16167
rect 6365 16127 6423 16133
rect 6914 16124 6920 16176
rect 6972 16124 6978 16176
rect 7006 16124 7012 16176
rect 7064 16164 7070 16176
rect 7944 16173 7972 16204
rect 8938 16192 8944 16204
rect 8996 16192 9002 16244
rect 9585 16235 9643 16241
rect 9585 16201 9597 16235
rect 9631 16232 9643 16235
rect 10226 16232 10232 16244
rect 9631 16204 10232 16232
rect 9631 16201 9643 16204
rect 9585 16195 9643 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 11238 16192 11244 16244
rect 11296 16192 11302 16244
rect 12894 16192 12900 16244
rect 12952 16232 12958 16244
rect 13446 16232 13452 16244
rect 12952 16204 13452 16232
rect 12952 16192 12958 16204
rect 13446 16192 13452 16204
rect 13504 16232 13510 16244
rect 18417 16235 18475 16241
rect 13504 16204 15976 16232
rect 13504 16192 13510 16204
rect 7101 16167 7159 16173
rect 7101 16164 7113 16167
rect 7064 16136 7113 16164
rect 7064 16124 7070 16136
rect 7101 16133 7113 16136
rect 7147 16164 7159 16167
rect 7929 16167 7987 16173
rect 7147 16136 7696 16164
rect 7147 16133 7159 16136
rect 7101 16127 7159 16133
rect 6932 16096 6960 16124
rect 7466 16096 7472 16108
rect 5828 16068 7472 16096
rect 7466 16056 7472 16068
rect 7524 16056 7530 16108
rect 7668 16105 7696 16136
rect 7929 16133 7941 16167
rect 7975 16133 7987 16167
rect 11256 16164 11284 16192
rect 12710 16164 12716 16176
rect 11256 16136 11376 16164
rect 7929 16127 7987 16133
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 7653 16099 7711 16105
rect 10042 16100 10048 16108
rect 7653 16065 7665 16099
rect 7699 16065 7711 16099
rect 9968 16096 10048 16100
rect 9062 16072 10048 16096
rect 9062 16068 9982 16072
rect 7653 16059 7711 16065
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 16028 1639 16031
rect 1627 16000 1716 16028
rect 1627 15997 1639 16000
rect 1581 15991 1639 15997
rect 1688 15904 1716 16000
rect 1854 15988 1860 16040
rect 1912 15988 1918 16040
rect 3418 15988 3424 16040
rect 3476 16028 3482 16040
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 3476 16000 3617 16028
rect 3476 15988 3482 16000
rect 3605 15997 3617 16000
rect 3651 15997 3663 16031
rect 3605 15991 3663 15997
rect 3881 16031 3939 16037
rect 3881 15997 3893 16031
rect 3927 15997 3939 16031
rect 3881 15991 3939 15997
rect 4157 16031 4215 16037
rect 4157 15997 4169 16031
rect 4203 16028 4215 16031
rect 4246 16028 4252 16040
rect 4203 16000 4252 16028
rect 4203 15997 4215 16000
rect 4157 15991 4215 15997
rect 1670 15852 1676 15904
rect 1728 15892 1734 15904
rect 3896 15892 3924 15991
rect 4246 15988 4252 16000
rect 4304 16028 4310 16040
rect 5997 16031 6055 16037
rect 4304 16000 5856 16028
rect 4304 15988 4310 16000
rect 5828 15969 5856 16000
rect 5997 15997 6009 16031
rect 6043 16028 6055 16031
rect 6454 16028 6460 16040
rect 6043 16000 6460 16028
rect 6043 15997 6055 16000
rect 5997 15991 6055 15997
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 7576 16028 7604 16059
rect 10042 16056 10048 16072
rect 10100 16056 10106 16108
rect 11348 16105 11376 16136
rect 11716 16136 12716 16164
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 9766 16028 9772 16040
rect 7576 16000 9772 16028
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11716 16028 11744 16136
rect 12710 16124 12716 16136
rect 12768 16124 12774 16176
rect 14826 16124 14832 16176
rect 14884 16124 14890 16176
rect 12066 16056 12072 16108
rect 12124 16096 12130 16108
rect 12529 16099 12587 16105
rect 12529 16096 12541 16099
rect 12124 16068 12541 16096
rect 12124 16056 12130 16068
rect 12529 16065 12541 16068
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 15470 16056 15476 16108
rect 15528 16096 15534 16108
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15528 16068 15761 16096
rect 15528 16056 15534 16068
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 11103 16000 11744 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 12894 15988 12900 16040
rect 12952 15988 12958 16040
rect 13538 15988 13544 16040
rect 13596 15988 13602 16040
rect 13814 15988 13820 16040
rect 13872 15988 13878 16040
rect 15948 16037 15976 16204
rect 18417 16201 18429 16235
rect 18463 16232 18475 16235
rect 18598 16232 18604 16244
rect 18463 16204 18604 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 18598 16192 18604 16204
rect 18656 16232 18662 16244
rect 19242 16232 19248 16244
rect 18656 16204 19248 16232
rect 18656 16192 18662 16204
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19613 16235 19671 16241
rect 19613 16201 19625 16235
rect 19659 16201 19671 16235
rect 19613 16195 19671 16201
rect 17494 16124 17500 16176
rect 17552 16124 17558 16176
rect 19260 16164 19288 16192
rect 19628 16164 19656 16195
rect 19794 16192 19800 16244
rect 19852 16192 19858 16244
rect 19886 16192 19892 16244
rect 19944 16232 19950 16244
rect 19981 16235 20039 16241
rect 19981 16232 19993 16235
rect 19944 16204 19993 16232
rect 19944 16192 19950 16204
rect 19981 16201 19993 16204
rect 20027 16201 20039 16235
rect 19981 16195 20039 16201
rect 20898 16192 20904 16244
rect 20956 16232 20962 16244
rect 22370 16232 22376 16244
rect 20956 16204 22376 16232
rect 20956 16192 20962 16204
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 23014 16192 23020 16244
rect 23072 16192 23078 16244
rect 23293 16235 23351 16241
rect 23293 16201 23305 16235
rect 23339 16232 23351 16235
rect 23382 16232 23388 16244
rect 23339 16204 23388 16232
rect 23339 16201 23351 16204
rect 23293 16195 23351 16201
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 24026 16192 24032 16244
rect 24084 16192 24090 16244
rect 24946 16232 24952 16244
rect 24872 16204 24952 16232
rect 19260 16136 19380 16164
rect 19628 16136 20208 16164
rect 16390 16056 16396 16108
rect 16448 16056 16454 16108
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16632 16068 16681 16096
rect 16632 16056 16638 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 18414 16056 18420 16108
rect 18472 16096 18478 16108
rect 19352 16105 19380 16136
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18472 16068 19073 16096
rect 18472 16056 18478 16068
rect 19061 16065 19073 16068
rect 19107 16096 19119 16099
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 19107 16068 19257 16096
rect 19107 16065 19119 16068
rect 19061 16059 19119 16065
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19337 16099 19395 16105
rect 19337 16065 19349 16099
rect 19383 16065 19395 16099
rect 19337 16059 19395 16065
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 20180 16105 20208 16136
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 19576 16068 19901 16096
rect 19576 16056 19582 16068
rect 19889 16065 19901 16068
rect 19935 16065 19947 16099
rect 19889 16059 19947 16065
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16065 20223 16099
rect 23032 16096 23060 16192
rect 23474 16124 23480 16176
rect 23532 16164 23538 16176
rect 23750 16164 23756 16176
rect 23532 16136 23756 16164
rect 23532 16124 23538 16136
rect 23750 16124 23756 16136
rect 23808 16124 23814 16176
rect 23109 16099 23167 16105
rect 23109 16096 23121 16099
rect 23032 16068 23121 16096
rect 20165 16059 20223 16065
rect 23109 16065 23121 16068
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16096 23351 16099
rect 24044 16096 24072 16192
rect 23339 16068 24072 16096
rect 23339 16065 23351 16068
rect 23293 16059 23351 16065
rect 15841 16031 15899 16037
rect 15841 16028 15853 16031
rect 15580 16000 15853 16028
rect 5813 15963 5871 15969
rect 5813 15929 5825 15963
rect 5859 15960 5871 15963
rect 7377 15963 7435 15969
rect 7377 15960 7389 15963
rect 5859 15932 7389 15960
rect 5859 15929 5871 15932
rect 5813 15923 5871 15929
rect 7377 15929 7389 15932
rect 7423 15929 7435 15963
rect 7377 15923 7435 15929
rect 9401 15963 9459 15969
rect 9401 15929 9413 15963
rect 9447 15960 9459 15963
rect 9674 15960 9680 15972
rect 9447 15932 9680 15960
rect 9447 15929 9459 15932
rect 9401 15923 9459 15929
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 15381 15963 15439 15969
rect 15381 15960 15393 15963
rect 14844 15932 15393 15960
rect 5534 15892 5540 15904
rect 1728 15864 5540 15892
rect 1728 15852 1734 15864
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 11974 15852 11980 15904
rect 12032 15852 12038 15904
rect 13449 15895 13507 15901
rect 13449 15861 13461 15895
rect 13495 15892 13507 15895
rect 13906 15892 13912 15904
rect 13495 15864 13912 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 14844 15892 14872 15932
rect 15381 15929 15393 15932
rect 15427 15929 15439 15963
rect 15381 15923 15439 15929
rect 14056 15864 14872 15892
rect 14056 15852 14062 15864
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 15580 15892 15608 16000
rect 15841 15997 15853 16000
rect 15887 15997 15899 16031
rect 15841 15991 15899 15997
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 15997 15991 16031
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 15933 15991 15991 15997
rect 16684 16000 16957 16028
rect 16684 15972 16712 16000
rect 16945 15997 16957 16000
rect 16991 15997 17003 16031
rect 16945 15991 17003 15997
rect 22002 15988 22008 16040
rect 22060 16028 22066 16040
rect 23308 16028 23336 16059
rect 24578 16056 24584 16108
rect 24636 16056 24642 16108
rect 24872 16105 24900 16204
rect 24946 16192 24952 16204
rect 25004 16192 25010 16244
rect 25041 16235 25099 16241
rect 25041 16201 25053 16235
rect 25087 16232 25099 16235
rect 25406 16232 25412 16244
rect 25087 16204 25412 16232
rect 25087 16201 25099 16204
rect 25041 16195 25099 16201
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 25498 16192 25504 16244
rect 25556 16232 25562 16244
rect 25556 16204 26188 16232
rect 25556 16192 25562 16204
rect 25130 16164 25136 16176
rect 24964 16136 25136 16164
rect 24857 16099 24915 16105
rect 24857 16065 24869 16099
rect 24903 16065 24915 16099
rect 24857 16059 24915 16065
rect 22060 16000 23336 16028
rect 24673 16031 24731 16037
rect 22060 15988 22066 16000
rect 24673 15997 24685 16031
rect 24719 15997 24731 16031
rect 24673 15991 24731 15997
rect 24765 16031 24823 16037
rect 24765 15997 24777 16031
rect 24811 16028 24823 16031
rect 24964 16028 24992 16136
rect 25130 16124 25136 16136
rect 25188 16164 25194 16176
rect 25317 16167 25375 16173
rect 25317 16164 25329 16167
rect 25188 16136 25329 16164
rect 25188 16124 25194 16136
rect 25317 16133 25329 16136
rect 25363 16133 25375 16167
rect 25317 16127 25375 16133
rect 25590 16124 25596 16176
rect 25648 16164 25654 16176
rect 26160 16173 26188 16204
rect 25929 16167 25987 16173
rect 25929 16164 25941 16167
rect 25648 16136 25941 16164
rect 25648 16124 25654 16136
rect 25929 16133 25941 16136
rect 25975 16133 25987 16167
rect 25929 16127 25987 16133
rect 26145 16167 26203 16173
rect 26145 16133 26157 16167
rect 26191 16133 26203 16167
rect 26145 16127 26203 16133
rect 25038 16056 25044 16108
rect 25096 16056 25102 16108
rect 25406 16056 25412 16108
rect 25464 16056 25470 16108
rect 25501 16099 25559 16105
rect 25501 16065 25513 16099
rect 25547 16065 25559 16099
rect 25501 16059 25559 16065
rect 24811 16000 24992 16028
rect 25056 16028 25084 16056
rect 25516 16028 25544 16059
rect 25056 16000 25544 16028
rect 24811 15997 24823 16000
rect 24765 15991 24823 15997
rect 16206 15920 16212 15972
rect 16264 15920 16270 15972
rect 16666 15920 16672 15972
rect 16724 15920 16730 15972
rect 22922 15920 22928 15972
rect 22980 15960 22986 15972
rect 24688 15960 24716 15991
rect 25133 15963 25191 15969
rect 25133 15960 25145 15963
rect 22980 15932 25145 15960
rect 22980 15920 22986 15932
rect 25133 15929 25145 15932
rect 25179 15929 25191 15963
rect 25866 15960 25872 15972
rect 25133 15923 25191 15929
rect 25700 15932 25872 15960
rect 15344 15864 15608 15892
rect 15344 15852 15350 15864
rect 18506 15852 18512 15904
rect 18564 15852 18570 15904
rect 19426 15852 19432 15904
rect 19484 15852 19490 15904
rect 24578 15852 24584 15904
rect 24636 15892 24642 15904
rect 25314 15892 25320 15904
rect 24636 15864 25320 15892
rect 24636 15852 24642 15864
rect 25314 15852 25320 15864
rect 25372 15852 25378 15904
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 25700 15901 25728 15932
rect 25866 15920 25872 15932
rect 25924 15960 25930 15972
rect 25924 15932 26004 15960
rect 25924 15920 25930 15932
rect 25685 15895 25743 15901
rect 25685 15892 25697 15895
rect 25464 15864 25697 15892
rect 25464 15852 25470 15864
rect 25685 15861 25697 15864
rect 25731 15861 25743 15895
rect 25685 15855 25743 15861
rect 25774 15852 25780 15904
rect 25832 15852 25838 15904
rect 25976 15901 26004 15932
rect 25961 15895 26019 15901
rect 25961 15861 25973 15895
rect 26007 15861 26019 15895
rect 25961 15855 26019 15861
rect 1104 15802 26496 15824
rect 1104 15750 4124 15802
rect 4176 15750 4188 15802
rect 4240 15750 4252 15802
rect 4304 15750 4316 15802
rect 4368 15750 4380 15802
rect 4432 15750 10472 15802
rect 10524 15750 10536 15802
rect 10588 15750 10600 15802
rect 10652 15750 10664 15802
rect 10716 15750 10728 15802
rect 10780 15750 16820 15802
rect 16872 15750 16884 15802
rect 16936 15750 16948 15802
rect 17000 15750 17012 15802
rect 17064 15750 17076 15802
rect 17128 15750 23168 15802
rect 23220 15750 23232 15802
rect 23284 15750 23296 15802
rect 23348 15750 23360 15802
rect 23412 15750 23424 15802
rect 23476 15750 26496 15802
rect 1104 15728 26496 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 2133 15691 2191 15697
rect 2133 15688 2145 15691
rect 1912 15660 2145 15688
rect 1912 15648 1918 15660
rect 2133 15657 2145 15660
rect 2179 15657 2191 15691
rect 2133 15651 2191 15657
rect 3053 15691 3111 15697
rect 3053 15657 3065 15691
rect 3099 15688 3111 15691
rect 3142 15688 3148 15700
rect 3099 15660 3148 15688
rect 3099 15657 3111 15660
rect 3053 15651 3111 15657
rect 3142 15648 3148 15660
rect 3200 15648 3206 15700
rect 3421 15691 3479 15697
rect 3421 15657 3433 15691
rect 3467 15657 3479 15691
rect 3421 15651 3479 15657
rect 3436 15620 3464 15651
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 5776 15660 6285 15688
rect 5776 15648 5782 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 7742 15688 7748 15700
rect 6273 15651 6331 15657
rect 6380 15660 7748 15688
rect 6380 15620 6408 15660
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10192 15660 11836 15688
rect 10192 15648 10198 15660
rect 3436 15592 6408 15620
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 2314 15444 2320 15496
rect 2372 15444 2378 15496
rect 3145 15487 3203 15493
rect 3145 15453 3157 15487
rect 3191 15484 3203 15487
rect 3436 15484 3464 15592
rect 5442 15512 5448 15564
rect 5500 15512 5506 15564
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 6730 15552 6736 15564
rect 5592 15524 6736 15552
rect 5592 15512 5598 15524
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15552 8539 15555
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8527 15524 8953 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 9674 15512 9680 15564
rect 9732 15512 9738 15564
rect 10413 15555 10471 15561
rect 10413 15521 10425 15555
rect 10459 15552 10471 15555
rect 11238 15552 11244 15564
rect 10459 15524 11244 15552
rect 10459 15521 10471 15524
rect 10413 15515 10471 15521
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 3191 15456 3464 15484
rect 3605 15487 3663 15493
rect 3191 15453 3203 15456
rect 3145 15447 3203 15453
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 3620 15416 3648 15447
rect 4890 15444 4896 15496
rect 4948 15484 4954 15496
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 4948 15456 5273 15484
rect 4948 15444 4954 15456
rect 5261 15453 5273 15456
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 5353 15487 5411 15493
rect 5353 15453 5365 15487
rect 5399 15484 5411 15487
rect 6362 15484 6368 15496
rect 5399 15456 6368 15484
rect 5399 15453 5411 15456
rect 5353 15447 5411 15453
rect 6362 15444 6368 15456
rect 6420 15444 6426 15496
rect 6454 15444 6460 15496
rect 6512 15444 6518 15496
rect 6638 15444 6644 15496
rect 6696 15444 6702 15496
rect 11808 15484 11836 15660
rect 12894 15648 12900 15700
rect 12952 15688 12958 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 12952 15660 13001 15688
rect 12952 15648 12958 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 12989 15651 13047 15657
rect 13262 15648 13268 15700
rect 13320 15648 13326 15700
rect 13538 15648 13544 15700
rect 13596 15648 13602 15700
rect 13725 15691 13783 15697
rect 13725 15657 13737 15691
rect 13771 15688 13783 15691
rect 13814 15688 13820 15700
rect 13771 15660 13820 15688
rect 13771 15657 13783 15660
rect 13725 15651 13783 15657
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 13906 15648 13912 15700
rect 13964 15648 13970 15700
rect 14550 15648 14556 15700
rect 14608 15688 14614 15700
rect 15010 15688 15016 15700
rect 14608 15660 15016 15688
rect 14608 15648 14614 15660
rect 15010 15648 15016 15660
rect 15068 15688 15074 15700
rect 15841 15691 15899 15697
rect 15841 15688 15853 15691
rect 15068 15660 15853 15688
rect 15068 15648 15074 15660
rect 15841 15657 15853 15660
rect 15887 15657 15899 15691
rect 15841 15651 15899 15657
rect 16666 15648 16672 15700
rect 16724 15648 16730 15700
rect 18506 15648 18512 15700
rect 18564 15648 18570 15700
rect 21082 15648 21088 15700
rect 21140 15688 21146 15700
rect 21269 15691 21327 15697
rect 21269 15688 21281 15691
rect 21140 15660 21281 15688
rect 21140 15648 21146 15660
rect 21269 15657 21281 15660
rect 21315 15657 21327 15691
rect 21269 15651 21327 15657
rect 12161 15555 12219 15561
rect 12161 15521 12173 15555
rect 12207 15552 12219 15555
rect 12805 15555 12863 15561
rect 12805 15552 12817 15555
rect 12207 15524 12817 15552
rect 12207 15521 12219 15524
rect 12161 15515 12219 15521
rect 12805 15521 12817 15524
rect 12851 15521 12863 15555
rect 12805 15515 12863 15521
rect 12618 15484 12624 15496
rect 11808 15470 12624 15484
rect 11822 15456 12624 15470
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15484 13231 15487
rect 13280 15484 13308 15648
rect 13556 15552 13584 15648
rect 13924 15620 13952 15648
rect 16684 15620 16712 15648
rect 16761 15623 16819 15629
rect 16761 15620 16773 15623
rect 13924 15592 14228 15620
rect 16684 15592 16773 15620
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 13556 15524 14105 15552
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 14200 15552 14228 15592
rect 16761 15589 16773 15592
rect 16807 15589 16819 15623
rect 16761 15583 16819 15589
rect 16945 15623 17003 15629
rect 16945 15589 16957 15623
rect 16991 15589 17003 15623
rect 16945 15583 17003 15589
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 14200 15524 14381 15552
rect 14093 15515 14151 15521
rect 14369 15521 14381 15524
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 14826 15512 14832 15564
rect 14884 15552 14890 15564
rect 15562 15552 15568 15564
rect 14884 15524 15568 15552
rect 14884 15512 14890 15524
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 13219 15456 13308 15484
rect 13219 15453 13231 15456
rect 13173 15447 13231 15453
rect 13446 15444 13452 15496
rect 13504 15444 13510 15496
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15484 13967 15487
rect 13998 15484 14004 15496
rect 13955 15456 14004 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 13998 15444 14004 15456
rect 14056 15444 14062 15496
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15484 16635 15487
rect 16960 15484 16988 15583
rect 17589 15555 17647 15561
rect 17589 15521 17601 15555
rect 17635 15552 17647 15555
rect 18322 15552 18328 15564
rect 17635 15524 18328 15552
rect 17635 15521 17647 15524
rect 17589 15515 17647 15521
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 18524 15552 18552 15648
rect 19521 15555 19579 15561
rect 18524 15524 18736 15552
rect 16623 15456 16988 15484
rect 18340 15484 18368 15512
rect 18340 15456 18552 15484
rect 16623 15453 16635 15456
rect 16577 15447 16635 15453
rect 6549 15419 6607 15425
rect 3344 15388 5028 15416
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 3344 15348 3372 15388
rect 1627 15320 3372 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 4890 15308 4896 15360
rect 4948 15308 4954 15360
rect 5000 15348 5028 15388
rect 6549 15385 6561 15419
rect 6595 15416 6607 15419
rect 7009 15419 7067 15425
rect 7009 15416 7021 15419
rect 6595 15388 7021 15416
rect 6595 15385 6607 15388
rect 6549 15379 6607 15385
rect 7009 15385 7021 15388
rect 7055 15385 7067 15419
rect 7009 15379 7067 15385
rect 7466 15376 7472 15428
rect 7524 15376 7530 15428
rect 10689 15419 10747 15425
rect 8312 15388 10456 15416
rect 8312 15348 8340 15388
rect 5000 15320 8340 15348
rect 9585 15351 9643 15357
rect 9585 15317 9597 15351
rect 9631 15348 9643 15351
rect 10134 15348 10140 15360
rect 9631 15320 10140 15348
rect 9631 15317 9643 15320
rect 9585 15311 9643 15317
rect 10134 15308 10140 15320
rect 10192 15308 10198 15360
rect 10318 15308 10324 15360
rect 10376 15308 10382 15360
rect 10428 15348 10456 15388
rect 10689 15385 10701 15419
rect 10735 15416 10747 15419
rect 10962 15416 10968 15428
rect 10735 15388 10968 15416
rect 10735 15385 10747 15388
rect 10689 15379 10747 15385
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 11992 15388 14780 15416
rect 11992 15348 12020 15388
rect 10428 15320 12020 15348
rect 12250 15308 12256 15360
rect 12308 15308 12314 15360
rect 13357 15351 13415 15357
rect 13357 15317 13369 15351
rect 13403 15348 13415 15351
rect 14550 15348 14556 15360
rect 13403 15320 14556 15348
rect 13403 15317 13415 15320
rect 13357 15311 13415 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 14752 15348 14780 15388
rect 14826 15376 14832 15428
rect 14884 15376 14890 15428
rect 17313 15419 17371 15425
rect 17313 15385 17325 15419
rect 17359 15416 17371 15419
rect 18414 15416 18420 15428
rect 17359 15388 18420 15416
rect 17359 15385 17371 15388
rect 17313 15379 17371 15385
rect 18414 15376 18420 15388
rect 18472 15376 18478 15428
rect 18524 15416 18552 15456
rect 18598 15444 18604 15496
rect 18656 15444 18662 15496
rect 18708 15493 18736 15524
rect 19521 15521 19533 15555
rect 19567 15552 19579 15555
rect 19886 15552 19892 15564
rect 19567 15524 19892 15552
rect 19567 15521 19579 15524
rect 19521 15515 19579 15521
rect 19886 15512 19892 15524
rect 19944 15512 19950 15564
rect 20898 15552 20904 15564
rect 20640 15524 20904 15552
rect 18693 15487 18751 15493
rect 18693 15453 18705 15487
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 19242 15444 19248 15496
rect 19300 15444 19306 15496
rect 20640 15470 20668 15524
rect 20898 15512 20904 15524
rect 20956 15552 20962 15564
rect 21100 15552 21128 15648
rect 20956 15524 21128 15552
rect 22465 15555 22523 15561
rect 20956 15512 20962 15524
rect 22465 15521 22477 15555
rect 22511 15521 22523 15555
rect 22465 15515 22523 15521
rect 22741 15555 22799 15561
rect 22741 15521 22753 15555
rect 22787 15552 22799 15555
rect 23106 15552 23112 15564
rect 22787 15524 23112 15552
rect 22787 15521 22799 15524
rect 22741 15515 22799 15521
rect 21174 15444 21180 15496
rect 21232 15444 21238 15496
rect 22370 15444 22376 15496
rect 22428 15444 22434 15496
rect 22480 15484 22508 15515
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 24578 15512 24584 15564
rect 24636 15512 24642 15564
rect 25774 15552 25780 15564
rect 24688 15524 25780 15552
rect 23934 15484 23940 15496
rect 22480 15456 23940 15484
rect 23934 15444 23940 15456
rect 23992 15484 23998 15496
rect 24596 15484 24624 15512
rect 24688 15493 24716 15524
rect 25774 15512 25780 15524
rect 25832 15512 25838 15564
rect 23992 15456 24624 15484
rect 24673 15487 24731 15493
rect 23992 15444 23998 15456
rect 24673 15453 24685 15487
rect 24719 15453 24731 15487
rect 24673 15447 24731 15453
rect 24946 15444 24952 15496
rect 25004 15444 25010 15496
rect 26050 15444 26056 15496
rect 26108 15444 26114 15496
rect 19610 15416 19616 15428
rect 18524 15388 19616 15416
rect 19610 15376 19616 15388
rect 19668 15376 19674 15428
rect 24210 15376 24216 15428
rect 24268 15416 24274 15428
rect 26068 15416 26096 15444
rect 24268 15388 26096 15416
rect 24268 15376 24274 15388
rect 15194 15348 15200 15360
rect 14752 15320 15200 15348
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 17405 15351 17463 15357
rect 17405 15317 17417 15351
rect 17451 15348 17463 15351
rect 17957 15351 18015 15357
rect 17957 15348 17969 15351
rect 17451 15320 17969 15348
rect 17451 15317 17463 15320
rect 17405 15311 17463 15317
rect 17957 15317 17969 15320
rect 18003 15317 18015 15351
rect 17957 15311 18015 15317
rect 18782 15308 18788 15360
rect 18840 15308 18846 15360
rect 20993 15351 21051 15357
rect 20993 15317 21005 15351
rect 21039 15348 21051 15351
rect 21082 15348 21088 15360
rect 21039 15320 21088 15348
rect 21039 15317 21051 15320
rect 20993 15311 21051 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 24486 15308 24492 15360
rect 24544 15308 24550 15360
rect 24857 15351 24915 15357
rect 24857 15317 24869 15351
rect 24903 15348 24915 15351
rect 25409 15351 25467 15357
rect 25409 15348 25421 15351
rect 24903 15320 25421 15348
rect 24903 15317 24915 15320
rect 24857 15311 24915 15317
rect 25409 15317 25421 15320
rect 25455 15317 25467 15351
rect 25409 15311 25467 15317
rect 1104 15258 26656 15280
rect 1104 15206 7298 15258
rect 7350 15206 7362 15258
rect 7414 15206 7426 15258
rect 7478 15206 7490 15258
rect 7542 15206 7554 15258
rect 7606 15206 13646 15258
rect 13698 15206 13710 15258
rect 13762 15206 13774 15258
rect 13826 15206 13838 15258
rect 13890 15206 13902 15258
rect 13954 15206 19994 15258
rect 20046 15206 20058 15258
rect 20110 15206 20122 15258
rect 20174 15206 20186 15258
rect 20238 15206 20250 15258
rect 20302 15206 26342 15258
rect 26394 15206 26406 15258
rect 26458 15206 26470 15258
rect 26522 15206 26534 15258
rect 26586 15206 26598 15258
rect 26650 15206 26656 15258
rect 1104 15184 26656 15206
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 6512 15116 6561 15144
rect 6512 15104 6518 15116
rect 6549 15113 6561 15116
rect 6595 15113 6607 15147
rect 9217 15147 9275 15153
rect 9217 15144 9229 15147
rect 6549 15107 6607 15113
rect 6656 15116 9229 15144
rect 3142 15076 3148 15088
rect 3082 15048 3148 15076
rect 3142 15036 3148 15048
rect 3200 15036 3206 15088
rect 6656 15017 6684 15116
rect 9217 15113 9229 15116
rect 9263 15113 9275 15147
rect 9217 15107 9275 15113
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 9732 15116 10057 15144
rect 9732 15104 9738 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 10045 15107 10103 15113
rect 10318 15104 10324 15156
rect 10376 15104 10382 15156
rect 10410 15104 10416 15156
rect 10468 15104 10474 15156
rect 10870 15104 10876 15156
rect 10928 15104 10934 15156
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 11885 15147 11943 15153
rect 11885 15113 11897 15147
rect 11931 15144 11943 15147
rect 12250 15144 12256 15156
rect 11931 15116 12256 15144
rect 11931 15113 11943 15116
rect 11885 15107 11943 15113
rect 8878 15048 10088 15076
rect 10060 15020 10088 15048
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 6788 14980 7389 15008
rect 6788 14968 6794 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 9953 15011 10011 15017
rect 9953 15008 9965 15011
rect 7377 14971 7435 14977
rect 9048 14980 9965 15008
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14940 1639 14943
rect 1857 14943 1915 14949
rect 1627 14912 1716 14940
rect 1627 14909 1639 14912
rect 1581 14903 1639 14909
rect 1688 14816 1716 14912
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 2406 14940 2412 14952
rect 1903 14912 2412 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3292 14912 3617 14940
rect 3292 14900 3298 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 7650 14900 7656 14952
rect 7708 14900 7714 14952
rect 8754 14832 8760 14884
rect 8812 14872 8818 14884
rect 9048 14872 9076 14980
rect 9953 14977 9965 14980
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 10042 14968 10048 15020
rect 10100 14968 10106 15020
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10229 15011 10287 15017
rect 10229 15008 10241 15011
rect 10192 14980 10241 15008
rect 10192 14968 10198 14980
rect 10229 14977 10241 14980
rect 10275 14977 10287 15011
rect 10336 15008 10364 15104
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10336 14980 10517 15008
rect 10229 14971 10287 14977
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 15008 11115 15011
rect 11532 15008 11560 15107
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 17494 15144 17500 15156
rect 17144 15116 17500 15144
rect 13446 15076 13452 15088
rect 12452 15048 13452 15076
rect 12345 15011 12403 15017
rect 12345 15008 12357 15011
rect 11103 14980 11560 15008
rect 11992 14980 12357 15008
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 9582 14940 9588 14952
rect 8812 14844 9076 14872
rect 9140 14912 9588 14940
rect 8812 14832 8818 14844
rect 1670 14764 1676 14816
rect 1728 14764 1734 14816
rect 8662 14764 8668 14816
rect 8720 14804 8726 14816
rect 9140 14813 9168 14912
rect 9582 14900 9588 14912
rect 9640 14940 9646 14952
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 9640 14912 9781 14940
rect 9640 14900 9646 14912
rect 9769 14909 9781 14912
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 11992 14949 12020 14980
rect 12345 14977 12357 14980
rect 12391 15008 12403 15011
rect 12452 15008 12480 15048
rect 13446 15036 13452 15048
rect 13504 15036 13510 15088
rect 12391 14980 12480 15008
rect 12391 14977 12403 14980
rect 12345 14971 12403 14977
rect 12526 14968 12532 15020
rect 12584 14968 12590 15020
rect 13814 14968 13820 15020
rect 13872 14968 13878 15020
rect 17144 15017 17172 15116
rect 17494 15104 17500 15116
rect 17552 15144 17558 15156
rect 19242 15144 19248 15156
rect 17552 15116 19248 15144
rect 17552 15104 17558 15116
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 22370 15144 22376 15156
rect 19444 15116 22376 15144
rect 17954 15036 17960 15088
rect 18012 15036 18018 15088
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 19334 14968 19340 15020
rect 19392 14968 19398 15020
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 11572 14912 11989 14940
rect 11572 14900 11578 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 12066 14900 12072 14952
rect 12124 14900 12130 14952
rect 17402 14900 17408 14952
rect 17460 14900 17466 14952
rect 18874 14900 18880 14952
rect 18932 14940 18938 14952
rect 19444 14940 19472 15116
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 22830 15104 22836 15156
rect 22888 15144 22894 15156
rect 23658 15144 23664 15156
rect 22888 15116 23664 15144
rect 22888 15104 22894 15116
rect 23658 15104 23664 15116
rect 23716 15144 23722 15156
rect 24213 15147 24271 15153
rect 23716 15116 24072 15144
rect 23716 15104 23722 15116
rect 19889 15079 19947 15085
rect 19889 15076 19901 15079
rect 18932 14912 19472 14940
rect 19536 15048 19901 15076
rect 18932 14900 18938 14912
rect 19536 14881 19564 15048
rect 19889 15045 19901 15048
rect 19935 15045 19947 15079
rect 19889 15039 19947 15045
rect 20898 15036 20904 15088
rect 20956 15036 20962 15088
rect 22278 15036 22284 15088
rect 22336 15036 22342 15088
rect 22646 15036 22652 15088
rect 22704 15076 22710 15088
rect 23109 15079 23167 15085
rect 23109 15076 23121 15079
rect 22704 15048 23121 15076
rect 22704 15036 22710 15048
rect 23109 15045 23121 15048
rect 23155 15045 23167 15079
rect 23109 15039 23167 15045
rect 23842 15036 23848 15088
rect 23900 15036 23906 15088
rect 22296 15008 22324 15036
rect 24044 15017 24072 15116
rect 24213 15113 24225 15147
rect 24259 15144 24271 15147
rect 24946 15144 24952 15156
rect 24259 15116 24952 15144
rect 24259 15113 24271 15116
rect 24213 15107 24271 15113
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 26050 15104 26056 15156
rect 26108 15104 26114 15156
rect 24486 15036 24492 15088
rect 24544 15076 24550 15088
rect 24581 15079 24639 15085
rect 24581 15076 24593 15079
rect 24544 15048 24593 15076
rect 24544 15036 24550 15048
rect 24581 15045 24593 15048
rect 24627 15045 24639 15079
rect 24581 15039 24639 15045
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 24912 15048 25070 15076
rect 24912 15036 24918 15048
rect 22373 15011 22431 15017
rect 22373 15008 22385 15011
rect 22296 14980 22385 15008
rect 22373 14977 22385 14980
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 14977 23443 15011
rect 23385 14971 23443 14977
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 15008 23811 15011
rect 24029 15011 24087 15017
rect 23799 14980 23980 15008
rect 23799 14977 23811 14980
rect 23753 14971 23811 14977
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 19521 14875 19579 14881
rect 19521 14841 19533 14875
rect 19567 14841 19579 14875
rect 19521 14835 19579 14841
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 8720 14776 9137 14804
rect 8720 14764 8726 14776
rect 9125 14773 9137 14776
rect 9171 14773 9183 14807
rect 9125 14767 9183 14773
rect 9950 14764 9956 14816
rect 10008 14804 10014 14816
rect 10597 14807 10655 14813
rect 10597 14804 10609 14807
rect 10008 14776 10609 14804
rect 10008 14764 10014 14776
rect 10597 14773 10609 14776
rect 10643 14773 10655 14807
rect 10597 14767 10655 14773
rect 12342 14764 12348 14816
rect 12400 14764 12406 14816
rect 15102 14764 15108 14816
rect 15160 14764 15166 14816
rect 19628 14804 19656 14903
rect 23014 14900 23020 14952
rect 23072 14900 23078 14952
rect 23293 14943 23351 14949
rect 23293 14909 23305 14943
rect 23339 14909 23351 14943
rect 23400 14940 23428 14971
rect 23400 14912 23888 14940
rect 23293 14903 23351 14909
rect 23308 14872 23336 14903
rect 23658 14872 23664 14884
rect 23308 14844 23664 14872
rect 23658 14832 23664 14844
rect 23716 14832 23722 14884
rect 23860 14816 23888 14912
rect 23952 14872 23980 14980
rect 24029 14977 24041 15011
rect 24075 15008 24087 15011
rect 24118 15008 24124 15020
rect 24075 14980 24124 15008
rect 24075 14977 24087 14980
rect 24029 14971 24087 14977
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 25590 14968 25596 15020
rect 25648 14968 25654 15020
rect 24302 14900 24308 14952
rect 24360 14900 24366 14952
rect 25222 14940 25228 14952
rect 24412 14912 25228 14940
rect 24412 14872 24440 14912
rect 25222 14900 25228 14912
rect 25280 14940 25286 14952
rect 25608 14940 25636 14968
rect 25280 14912 25636 14940
rect 25280 14900 25286 14912
rect 23952 14844 24440 14872
rect 19886 14804 19892 14816
rect 19628 14776 19892 14804
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 21358 14764 21364 14816
rect 21416 14764 21422 14816
rect 23106 14764 23112 14816
rect 23164 14764 23170 14816
rect 23566 14764 23572 14816
rect 23624 14764 23630 14816
rect 23842 14764 23848 14816
rect 23900 14764 23906 14816
rect 24118 14764 24124 14816
rect 24176 14804 24182 14816
rect 25130 14804 25136 14816
rect 24176 14776 25136 14804
rect 24176 14764 24182 14776
rect 25130 14764 25136 14776
rect 25188 14804 25194 14816
rect 25682 14804 25688 14816
rect 25188 14776 25688 14804
rect 25188 14764 25194 14776
rect 25682 14764 25688 14776
rect 25740 14764 25746 14816
rect 1104 14714 26496 14736
rect 1104 14662 4124 14714
rect 4176 14662 4188 14714
rect 4240 14662 4252 14714
rect 4304 14662 4316 14714
rect 4368 14662 4380 14714
rect 4432 14662 10472 14714
rect 10524 14662 10536 14714
rect 10588 14662 10600 14714
rect 10652 14662 10664 14714
rect 10716 14662 10728 14714
rect 10780 14662 16820 14714
rect 16872 14662 16884 14714
rect 16936 14662 16948 14714
rect 17000 14662 17012 14714
rect 17064 14662 17076 14714
rect 17128 14662 23168 14714
rect 23220 14662 23232 14714
rect 23284 14662 23296 14714
rect 23348 14662 23360 14714
rect 23412 14662 23424 14714
rect 23476 14662 26496 14714
rect 1104 14640 26496 14662
rect 2314 14560 2320 14612
rect 2372 14560 2378 14612
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 6696 14572 7604 14600
rect 6696 14560 6702 14572
rect 7576 14532 7604 14572
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7745 14603 7803 14609
rect 7745 14600 7757 14603
rect 7708 14572 7757 14600
rect 7708 14560 7714 14572
rect 7745 14569 7757 14572
rect 7791 14569 7803 14603
rect 7745 14563 7803 14569
rect 7944 14572 8340 14600
rect 7944 14532 7972 14572
rect 7576 14504 7972 14532
rect 8021 14535 8079 14541
rect 8021 14501 8033 14535
rect 8067 14501 8079 14535
rect 8021 14495 8079 14501
rect 2961 14467 3019 14473
rect 2961 14464 2973 14467
rect 2148 14436 2973 14464
rect 2148 14405 2176 14436
rect 2961 14433 2973 14436
rect 3007 14464 3019 14467
rect 4706 14464 4712 14476
rect 3007 14436 4712 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14365 2283 14399
rect 2225 14359 2283 14365
rect 1946 14288 1952 14340
rect 2004 14288 2010 14340
rect 2240 14328 2268 14359
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 3329 14399 3387 14405
rect 3329 14396 3341 14399
rect 3292 14368 3341 14396
rect 3292 14356 3298 14368
rect 3329 14365 3341 14368
rect 3375 14365 3387 14399
rect 3329 14359 3387 14365
rect 3418 14356 3424 14408
rect 3476 14396 3482 14408
rect 3620 14405 3648 14436
rect 4706 14424 4712 14436
rect 4764 14464 4770 14476
rect 5442 14464 5448 14476
rect 4764 14436 5448 14464
rect 4764 14424 4770 14436
rect 5442 14424 5448 14436
rect 5500 14464 5506 14476
rect 5500 14436 5580 14464
rect 5500 14424 5506 14436
rect 5552 14405 5580 14436
rect 3605 14399 3663 14405
rect 3605 14396 3617 14399
rect 3476 14368 3617 14396
rect 3476 14356 3482 14368
rect 3605 14365 3617 14368
rect 3651 14365 3663 14399
rect 3605 14359 3663 14365
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14365 5411 14399
rect 5353 14359 5411 14365
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14396 5595 14399
rect 5583 14368 5672 14396
rect 5583 14365 5595 14368
rect 5537 14359 5595 14365
rect 3050 14328 3056 14340
rect 2240 14300 3056 14328
rect 3050 14288 3056 14300
rect 3108 14328 3114 14340
rect 3513 14331 3571 14337
rect 3513 14328 3525 14331
rect 3108 14300 3525 14328
rect 3108 14288 3114 14300
rect 3513 14297 3525 14300
rect 3559 14328 3571 14331
rect 4798 14328 4804 14340
rect 3559 14300 4804 14328
rect 3559 14297 3571 14300
rect 3513 14291 3571 14297
rect 2222 14220 2228 14272
rect 2280 14220 2286 14272
rect 2682 14220 2688 14272
rect 2740 14220 2746 14272
rect 2777 14263 2835 14269
rect 2777 14229 2789 14263
rect 2823 14260 2835 14263
rect 2866 14260 2872 14272
rect 2823 14232 2872 14260
rect 2823 14229 2835 14232
rect 2777 14223 2835 14229
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 3142 14220 3148 14272
rect 3200 14220 3206 14272
rect 3528 14260 3556 14291
rect 4798 14288 4804 14300
rect 4856 14328 4862 14340
rect 5368 14328 5396 14359
rect 5644 14328 5672 14368
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 5994 14396 6000 14408
rect 5776 14368 6000 14396
rect 5776 14356 5782 14368
rect 5994 14356 6000 14368
rect 6052 14396 6058 14408
rect 6733 14399 6791 14405
rect 6733 14396 6745 14399
rect 6052 14368 6745 14396
rect 6052 14356 6058 14368
rect 6733 14365 6745 14368
rect 6779 14365 6791 14399
rect 6733 14359 6791 14365
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 8036 14396 8064 14495
rect 8312 14464 8340 14572
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 12342 14609 12348 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 9640 14572 10241 14600
rect 9640 14560 9646 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 10229 14563 10287 14569
rect 12332 14603 12348 14609
rect 12332 14569 12344 14603
rect 12332 14563 12348 14569
rect 12342 14560 12348 14563
rect 12400 14560 12406 14612
rect 14921 14603 14979 14609
rect 14921 14569 14933 14603
rect 14967 14600 14979 14603
rect 15010 14600 15016 14612
rect 14967 14572 15016 14600
rect 14967 14569 14979 14572
rect 14921 14563 14979 14569
rect 15010 14560 15016 14572
rect 15068 14560 15074 14612
rect 16390 14560 16396 14612
rect 16448 14560 16454 14612
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 17589 14603 17647 14609
rect 17589 14600 17601 14603
rect 17460 14572 17601 14600
rect 17460 14560 17466 14572
rect 17589 14569 17601 14572
rect 17635 14569 17647 14603
rect 17589 14563 17647 14569
rect 18874 14560 18880 14612
rect 18932 14560 18938 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 20165 14603 20223 14609
rect 20165 14600 20177 14603
rect 19392 14572 20177 14600
rect 19392 14560 19398 14572
rect 20165 14569 20177 14572
rect 20211 14569 20223 14603
rect 20165 14563 20223 14569
rect 22830 14560 22836 14612
rect 22888 14560 22894 14612
rect 23750 14600 23756 14612
rect 23400 14572 23756 14600
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 10597 14535 10655 14541
rect 10597 14532 10609 14535
rect 9824 14504 10609 14532
rect 9824 14492 9830 14504
rect 10597 14501 10609 14504
rect 10643 14501 10655 14535
rect 10597 14495 10655 14501
rect 14553 14535 14611 14541
rect 14553 14501 14565 14535
rect 14599 14532 14611 14535
rect 16408 14532 16436 14560
rect 14599 14504 16436 14532
rect 14599 14501 14611 14504
rect 14553 14495 14611 14501
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 18693 14535 18751 14541
rect 18693 14532 18705 14535
rect 18472 14504 18705 14532
rect 18472 14492 18478 14504
rect 18693 14501 18705 14504
rect 18739 14501 18751 14535
rect 18693 14495 18751 14501
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8312 14436 8585 14464
rect 8573 14433 8585 14436
rect 8619 14464 8631 14467
rect 8754 14464 8760 14476
rect 8619 14436 8760 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11296 14436 12081 14464
rect 11296 14424 11302 14436
rect 12069 14433 12081 14436
rect 12115 14464 12127 14467
rect 14829 14467 14887 14473
rect 12115 14436 14228 14464
rect 12115 14433 12127 14436
rect 12069 14427 12127 14433
rect 7975 14368 8064 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 8352 14368 9505 14396
rect 8352 14356 8358 14368
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 9674 14356 9680 14408
rect 9732 14396 9738 14408
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 9732 14368 10241 14396
rect 9732 14356 9738 14368
rect 10229 14365 10241 14368
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 10318 14356 10324 14408
rect 10376 14356 10382 14408
rect 6822 14328 6828 14340
rect 4856 14300 5580 14328
rect 5644 14300 6828 14328
rect 4856 14288 4862 14300
rect 5552 14272 5580 14300
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 9769 14331 9827 14337
rect 9769 14297 9781 14331
rect 9815 14328 9827 14331
rect 9858 14328 9864 14340
rect 9815 14300 9864 14328
rect 9815 14297 9827 14300
rect 9769 14291 9827 14297
rect 9858 14288 9864 14300
rect 9916 14328 9922 14340
rect 10134 14328 10140 14340
rect 9916 14300 10140 14328
rect 9916 14288 9922 14300
rect 10134 14288 10140 14300
rect 10192 14328 10198 14340
rect 10192 14300 12434 14328
rect 10192 14288 10198 14300
rect 12406 14272 12434 14300
rect 12618 14288 12624 14340
rect 12676 14328 12682 14340
rect 12676 14300 12834 14328
rect 12676 14288 12682 14300
rect 14200 14272 14228 14436
rect 14829 14433 14841 14467
rect 14875 14464 14887 14467
rect 15286 14464 15292 14476
rect 14875 14436 15292 14464
rect 14875 14433 14887 14436
rect 14829 14427 14887 14433
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 18892 14464 18920 14560
rect 22186 14492 22192 14544
rect 22244 14532 22250 14544
rect 23400 14541 23428 14572
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 23842 14560 23848 14612
rect 23900 14560 23906 14612
rect 24026 14560 24032 14612
rect 24084 14560 24090 14612
rect 23385 14535 23443 14541
rect 22244 14504 23244 14532
rect 22244 14492 22250 14504
rect 18524 14436 18920 14464
rect 20809 14467 20867 14473
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14396 14979 14399
rect 15930 14396 15936 14408
rect 14967 14368 15936 14396
rect 14967 14365 14979 14368
rect 14921 14359 14979 14365
rect 15930 14356 15936 14368
rect 15988 14396 15994 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15988 14368 16129 14396
rect 15988 14356 15994 14368
rect 16117 14365 16129 14368
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14396 17555 14399
rect 17586 14396 17592 14408
rect 17543 14368 17592 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 16592 14328 16620 14359
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 18524 14405 18552 14436
rect 20809 14433 20821 14467
rect 20855 14464 20867 14467
rect 21358 14464 21364 14476
rect 20855 14436 21364 14464
rect 20855 14433 20867 14436
rect 20809 14427 20867 14433
rect 21358 14424 21364 14436
rect 21416 14464 21422 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 21416 14436 22293 14464
rect 21416 14424 21422 14436
rect 22281 14433 22293 14436
rect 22327 14464 22339 14467
rect 22465 14467 22523 14473
rect 22465 14464 22477 14467
rect 22327 14436 22477 14464
rect 22327 14433 22339 14436
rect 22281 14427 22339 14433
rect 22465 14433 22477 14436
rect 22511 14433 22523 14467
rect 22465 14427 22523 14433
rect 23014 14424 23020 14476
rect 23072 14424 23078 14476
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18325 14399 18383 14405
rect 18325 14396 18337 14399
rect 18279 14368 18337 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18325 14365 18337 14368
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14365 18567 14399
rect 18509 14359 18567 14365
rect 18601 14399 18659 14405
rect 18601 14365 18613 14399
rect 18647 14365 18659 14399
rect 18601 14359 18659 14365
rect 14700 14300 16620 14328
rect 18616 14328 18644 14359
rect 18782 14356 18788 14408
rect 18840 14396 18846 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 18840 14368 19257 14396
rect 18840 14356 18846 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 19610 14396 19616 14408
rect 19475 14368 19616 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 19610 14356 19616 14368
rect 19668 14396 19674 14408
rect 20622 14396 20628 14408
rect 19668 14368 20628 14396
rect 19668 14356 19674 14368
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 21082 14356 21088 14408
rect 21140 14396 21146 14408
rect 23216 14405 23244 14504
rect 23385 14501 23397 14535
rect 23431 14501 23443 14535
rect 24044 14532 24072 14560
rect 23385 14495 23443 14501
rect 23860 14504 24072 14532
rect 23584 14436 23796 14464
rect 23584 14408 23612 14436
rect 21545 14399 21603 14405
rect 21545 14396 21557 14399
rect 21140 14368 21557 14396
rect 21140 14356 21146 14368
rect 21545 14365 21557 14368
rect 21591 14365 21603 14399
rect 21545 14359 21603 14365
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14396 23259 14399
rect 23247 14368 23336 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 19518 14328 19524 14340
rect 18616 14300 19524 14328
rect 14700 14288 14706 14300
rect 19518 14288 19524 14300
rect 19576 14288 19582 14340
rect 20533 14331 20591 14337
rect 20533 14297 20545 14331
rect 20579 14328 20591 14331
rect 20993 14331 21051 14337
rect 20993 14328 21005 14331
rect 20579 14300 21005 14328
rect 20579 14297 20591 14300
rect 20533 14291 20591 14297
rect 20993 14297 21005 14300
rect 21039 14297 21051 14331
rect 20993 14291 21051 14297
rect 22664 14272 22692 14359
rect 23308 14328 23336 14368
rect 23566 14356 23572 14408
rect 23624 14356 23630 14408
rect 23768 14405 23796 14436
rect 23860 14405 23888 14504
rect 24949 14467 25007 14473
rect 24949 14464 24961 14467
rect 24044 14436 24961 14464
rect 23753 14399 23811 14405
rect 23753 14365 23765 14399
rect 23799 14365 23811 14399
rect 23753 14359 23811 14365
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14365 23903 14399
rect 23845 14359 23903 14365
rect 24044 14340 24072 14436
rect 24949 14433 24961 14436
rect 24995 14433 25007 14467
rect 24949 14427 25007 14433
rect 24121 14399 24179 14405
rect 24121 14365 24133 14399
rect 24167 14396 24179 14399
rect 24210 14396 24216 14408
rect 24167 14368 24216 14396
rect 24167 14365 24179 14368
rect 24121 14359 24179 14365
rect 24210 14356 24216 14368
rect 24268 14396 24274 14408
rect 25225 14399 25283 14405
rect 25225 14396 25237 14399
rect 24268 14368 25237 14396
rect 24268 14356 24274 14368
rect 25225 14365 25237 14368
rect 25271 14365 25283 14399
rect 25225 14359 25283 14365
rect 25406 14356 25412 14408
rect 25464 14356 25470 14408
rect 23937 14331 23995 14337
rect 23308 14300 23612 14328
rect 3602 14260 3608 14272
rect 3528 14232 3608 14260
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 5350 14220 5356 14272
rect 5408 14220 5414 14272
rect 5534 14220 5540 14272
rect 5592 14220 5598 14272
rect 7374 14220 7380 14272
rect 7432 14220 7438 14272
rect 8386 14220 8392 14272
rect 8444 14220 8450 14272
rect 8478 14220 8484 14272
rect 8536 14220 8542 14272
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8812 14232 8953 14260
rect 8812 14220 8818 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 10042 14220 10048 14272
rect 10100 14220 10106 14272
rect 12406 14232 12440 14272
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 13817 14263 13875 14269
rect 13817 14229 13829 14263
rect 13863 14260 13875 14263
rect 14090 14260 14096 14272
rect 13863 14232 14096 14260
rect 13863 14229 13875 14232
rect 13817 14223 13875 14229
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 14182 14220 14188 14272
rect 14240 14220 14246 14272
rect 15470 14220 15476 14272
rect 15528 14260 15534 14272
rect 15565 14263 15623 14269
rect 15565 14260 15577 14263
rect 15528 14232 15577 14260
rect 15528 14220 15534 14232
rect 15565 14229 15577 14232
rect 15611 14229 15623 14263
rect 15565 14223 15623 14229
rect 16666 14220 16672 14272
rect 16724 14220 16730 14272
rect 16850 14220 16856 14272
rect 16908 14220 16914 14272
rect 19334 14220 19340 14272
rect 19392 14220 19398 14272
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 21729 14263 21787 14269
rect 21729 14260 21741 14263
rect 20956 14232 21741 14260
rect 20956 14220 20962 14232
rect 21729 14229 21741 14232
rect 21775 14229 21787 14263
rect 21729 14223 21787 14229
rect 22646 14220 22652 14272
rect 22704 14220 22710 14272
rect 23584 14269 23612 14300
rect 23937 14297 23949 14331
rect 23983 14328 23995 14331
rect 24026 14328 24032 14340
rect 23983 14300 24032 14328
rect 23983 14297 23995 14300
rect 23937 14291 23995 14297
rect 24026 14288 24032 14300
rect 24084 14288 24090 14340
rect 24857 14331 24915 14337
rect 24857 14297 24869 14331
rect 24903 14328 24915 14331
rect 24946 14328 24952 14340
rect 24903 14300 24952 14328
rect 24903 14297 24915 14300
rect 24857 14291 24915 14297
rect 24946 14288 24952 14300
rect 25004 14288 25010 14340
rect 23569 14263 23627 14269
rect 23569 14229 23581 14263
rect 23615 14229 23627 14263
rect 23569 14223 23627 14229
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 24762 14220 24768 14272
rect 24820 14220 24826 14272
rect 25498 14220 25504 14272
rect 25556 14260 25562 14272
rect 25593 14263 25651 14269
rect 25593 14260 25605 14263
rect 25556 14232 25605 14260
rect 25556 14220 25562 14232
rect 25593 14229 25605 14232
rect 25639 14229 25651 14263
rect 25593 14223 25651 14229
rect 1104 14170 26656 14192
rect 1104 14118 7298 14170
rect 7350 14118 7362 14170
rect 7414 14118 7426 14170
rect 7478 14118 7490 14170
rect 7542 14118 7554 14170
rect 7606 14118 13646 14170
rect 13698 14118 13710 14170
rect 13762 14118 13774 14170
rect 13826 14118 13838 14170
rect 13890 14118 13902 14170
rect 13954 14118 19994 14170
rect 20046 14118 20058 14170
rect 20110 14118 20122 14170
rect 20174 14118 20186 14170
rect 20238 14118 20250 14170
rect 20302 14118 26342 14170
rect 26394 14118 26406 14170
rect 26458 14118 26470 14170
rect 26522 14118 26534 14170
rect 26586 14118 26598 14170
rect 26650 14118 26656 14170
rect 1104 14096 26656 14118
rect 1946 14016 1952 14068
rect 2004 14016 2010 14068
rect 2222 14016 2228 14068
rect 2280 14016 2286 14068
rect 2317 14059 2375 14065
rect 2317 14025 2329 14059
rect 2363 14056 2375 14059
rect 2406 14056 2412 14068
rect 2363 14028 2412 14056
rect 2363 14025 2375 14028
rect 2317 14019 2375 14025
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 3142 14056 3148 14068
rect 2608 14028 3148 14056
rect 1964 13852 1992 14016
rect 2240 13920 2268 14016
rect 2608 13997 2636 14028
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 3418 14016 3424 14068
rect 3476 14016 3482 14068
rect 5350 14056 5356 14068
rect 5092 14028 5356 14056
rect 2593 13991 2651 13997
rect 2593 13957 2605 13991
rect 2639 13957 2651 13991
rect 2593 13951 2651 13957
rect 3602 13948 3608 14000
rect 3660 13988 3666 14000
rect 4801 13991 4859 13997
rect 3660 13960 4568 13988
rect 3660 13948 3666 13960
rect 2501 13923 2559 13929
rect 2501 13920 2513 13923
rect 2240 13892 2513 13920
rect 2501 13889 2513 13892
rect 2547 13889 2559 13923
rect 2501 13883 2559 13889
rect 2682 13880 2688 13932
rect 2740 13880 2746 13932
rect 2866 13929 2872 13932
rect 2823 13923 2872 13929
rect 2823 13889 2835 13923
rect 2869 13889 2872 13923
rect 2823 13883 2872 13889
rect 2866 13880 2872 13883
rect 2924 13920 2930 13932
rect 2924 13892 3096 13920
rect 2924 13880 2930 13892
rect 2961 13855 3019 13861
rect 2961 13852 2973 13855
rect 1964 13824 2973 13852
rect 2961 13821 2973 13824
rect 3007 13821 3019 13855
rect 3068 13852 3096 13892
rect 3234 13880 3240 13932
rect 3292 13880 3298 13932
rect 4540 13929 4568 13960
rect 4801 13957 4813 13991
rect 4847 13988 4859 13991
rect 4847 13960 5028 13988
rect 4847 13957 4859 13960
rect 4801 13951 4859 13957
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13920 3387 13923
rect 4525 13923 4583 13929
rect 3375 13892 3648 13920
rect 3375 13889 3387 13892
rect 3329 13883 3387 13889
rect 3620 13864 3648 13892
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 4525 13883 4583 13889
rect 3068 13824 3372 13852
rect 2961 13815 3019 13821
rect 2976 13784 3004 13815
rect 3344 13784 3372 13824
rect 3602 13812 3608 13864
rect 3660 13812 3666 13864
rect 4706 13812 4712 13864
rect 4764 13852 4770 13864
rect 4801 13855 4859 13861
rect 4801 13852 4813 13855
rect 4764 13824 4813 13852
rect 4764 13812 4770 13824
rect 4801 13821 4813 13824
rect 4847 13821 4859 13855
rect 5000 13852 5028 13960
rect 5092 13929 5120 14028
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 5592 14028 6009 14056
rect 5592 14016 5598 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 5997 14019 6055 14025
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 15378 14056 15384 14068
rect 6788 14028 8984 14056
rect 6788 14016 6794 14028
rect 5261 13991 5319 13997
rect 5261 13957 5273 13991
rect 5307 13988 5319 13991
rect 7098 13988 7104 14000
rect 5307 13960 7104 13988
rect 5307 13957 5319 13960
rect 5261 13951 5319 13957
rect 7098 13948 7104 13960
rect 7156 13948 7162 14000
rect 8665 13991 8723 13997
rect 8665 13957 8677 13991
rect 8711 13988 8723 13991
rect 8754 13988 8760 14000
rect 8711 13960 8760 13988
rect 8711 13957 8723 13960
rect 8665 13951 8723 13957
rect 8754 13948 8760 13960
rect 8812 13948 8818 14000
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5166 13880 5172 13932
rect 5224 13880 5230 13932
rect 5350 13880 5356 13932
rect 5408 13929 5414 13932
rect 5408 13923 5437 13929
rect 5425 13889 5437 13923
rect 5408 13883 5437 13889
rect 5408 13880 5414 13883
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 8956 13929 8984 14028
rect 14108 14028 15384 14056
rect 11974 13948 11980 14000
rect 12032 13948 12038 14000
rect 13449 13991 13507 13997
rect 13449 13988 13461 13991
rect 13096 13960 13461 13988
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5644 13892 5825 13920
rect 5000 13844 5304 13852
rect 5000 13824 5488 13844
rect 4801 13815 4859 13821
rect 5276 13816 5488 13824
rect 5460 13784 5488 13816
rect 5644 13784 5672 13892
rect 5813 13889 5825 13892
rect 5859 13889 5871 13923
rect 5813 13883 5871 13889
rect 6089 13923 6147 13929
rect 6089 13889 6101 13923
rect 6135 13889 6147 13923
rect 8941 13923 8999 13929
rect 6089 13883 6147 13889
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 6104 13852 6132 13883
rect 5960 13824 6132 13852
rect 7576 13852 7604 13906
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9125 13923 9183 13929
rect 9125 13920 9137 13923
rect 8987 13892 9137 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9125 13889 9137 13892
rect 9171 13889 9183 13923
rect 9125 13883 9183 13889
rect 10042 13852 10048 13864
rect 7576 13824 10048 13852
rect 5960 13812 5966 13824
rect 10042 13812 10048 13824
rect 10100 13852 10106 13864
rect 10520 13852 10548 13906
rect 11514 13880 11520 13932
rect 11572 13880 11578 13932
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13920 11759 13923
rect 11992 13920 12020 13948
rect 13096 13929 13124 13960
rect 13449 13957 13461 13960
rect 13495 13957 13507 13991
rect 13449 13951 13507 13957
rect 11747 13892 12020 13920
rect 13081 13923 13139 13929
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 13081 13889 13093 13923
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 14108 13920 14136 14028
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 15930 14016 15936 14068
rect 15988 14016 15994 14068
rect 16393 14059 16451 14065
rect 16393 14025 16405 14059
rect 16439 14056 16451 14059
rect 16666 14056 16672 14068
rect 16439 14028 16672 14056
rect 16439 14025 16451 14028
rect 16393 14019 16451 14025
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 16850 14016 16856 14068
rect 16908 14016 16914 14068
rect 19242 14016 19248 14068
rect 19300 14016 19306 14068
rect 23934 14056 23940 14068
rect 23492 14028 23940 14056
rect 16868 13988 16896 14016
rect 16224 13960 16896 13988
rect 19260 13988 19288 14016
rect 19260 13960 19380 13988
rect 13403 13892 14136 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 12618 13852 12624 13864
rect 10100 13824 12624 13852
rect 10100 13812 10106 13824
rect 12618 13812 12624 13824
rect 12676 13812 12682 13864
rect 13280 13852 13308 13883
rect 14182 13880 14188 13932
rect 14240 13880 14246 13932
rect 15562 13880 15568 13932
rect 15620 13880 15626 13932
rect 16224 13929 16252 13960
rect 16209 13923 16267 13929
rect 16209 13889 16221 13923
rect 16255 13889 16267 13923
rect 16209 13883 16267 13889
rect 16485 13923 16543 13929
rect 16485 13889 16497 13923
rect 16531 13920 16543 13923
rect 16531 13892 17908 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 13280 13824 14044 13852
rect 2976 13756 3280 13784
rect 3344 13756 5396 13784
rect 5460 13756 5672 13784
rect 3252 13728 3280 13756
rect 5368 13728 5396 13756
rect 10870 13744 10876 13796
rect 10928 13784 10934 13796
rect 13906 13784 13912 13796
rect 10928 13756 13912 13784
rect 10928 13744 10934 13756
rect 13906 13744 13912 13756
rect 13964 13744 13970 13796
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 3053 13719 3111 13725
rect 3053 13716 3065 13719
rect 2832 13688 3065 13716
rect 2832 13676 2838 13688
rect 3053 13685 3065 13688
rect 3099 13685 3111 13719
rect 3053 13679 3111 13685
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 4614 13716 4620 13728
rect 3292 13688 4620 13716
rect 3292 13676 3298 13688
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 4893 13719 4951 13725
rect 4893 13685 4905 13719
rect 4939 13716 4951 13719
rect 4982 13716 4988 13728
rect 4939 13688 4988 13716
rect 4939 13685 4951 13688
rect 4893 13679 4951 13685
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 5350 13676 5356 13728
rect 5408 13676 5414 13728
rect 5626 13676 5632 13728
rect 5684 13676 5690 13728
rect 7006 13676 7012 13728
rect 7064 13716 7070 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 7064 13688 7205 13716
rect 7064 13676 7070 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 7193 13679 7251 13685
rect 9122 13676 9128 13728
rect 9180 13716 9186 13728
rect 9382 13719 9440 13725
rect 9382 13716 9394 13719
rect 9180 13688 9394 13716
rect 9180 13676 9186 13688
rect 9382 13685 9394 13688
rect 9428 13685 9440 13719
rect 9382 13679 9440 13685
rect 11606 13676 11612 13728
rect 11664 13676 11670 13728
rect 12894 13676 12900 13728
rect 12952 13676 12958 13728
rect 14016 13716 14044 13824
rect 14090 13812 14096 13864
rect 14148 13812 14154 13864
rect 14458 13812 14464 13864
rect 14516 13812 14522 13864
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13852 16083 13855
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16071 13824 16681 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 17880 13852 17908 13892
rect 17954 13880 17960 13932
rect 18012 13880 18018 13932
rect 19352 13929 19380 13960
rect 20806 13948 20812 14000
rect 20864 13948 20870 14000
rect 23014 13988 23020 14000
rect 22388 13960 23020 13988
rect 19337 13923 19395 13929
rect 19337 13889 19349 13923
rect 19383 13889 19395 13923
rect 22186 13920 22192 13932
rect 19337 13883 19395 13889
rect 21008 13892 22192 13920
rect 18046 13852 18052 13864
rect 17880 13824 18052 13852
rect 16669 13815 16727 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19705 13855 19763 13861
rect 19107 13824 19288 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 19260 13784 19288 13824
rect 19705 13821 19717 13855
rect 19751 13852 19763 13855
rect 19886 13852 19892 13864
rect 19751 13824 19892 13852
rect 19751 13821 19763 13824
rect 19705 13815 19763 13821
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13852 20131 13855
rect 20438 13852 20444 13864
rect 20119 13824 20444 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 20622 13812 20628 13864
rect 20680 13852 20686 13864
rect 21008 13852 21036 13892
rect 22186 13880 22192 13892
rect 22244 13880 22250 13932
rect 22388 13929 22416 13960
rect 23014 13948 23020 13960
rect 23072 13948 23078 14000
rect 23492 13929 23520 14028
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 24121 14059 24179 14065
rect 24121 14025 24133 14059
rect 24167 14056 24179 14059
rect 24762 14056 24768 14068
rect 24167 14028 24768 14056
rect 24167 14025 24179 14028
rect 24121 14019 24179 14025
rect 24762 14016 24768 14028
rect 24820 14016 24826 14068
rect 23658 13948 23664 14000
rect 23716 13948 23722 14000
rect 25498 13988 25504 14000
rect 23952 13960 25504 13988
rect 22373 13923 22431 13929
rect 22373 13889 22385 13923
rect 22419 13889 22431 13923
rect 22373 13883 22431 13889
rect 23477 13923 23535 13929
rect 23477 13889 23489 13923
rect 23523 13889 23535 13923
rect 23477 13883 23535 13889
rect 23569 13923 23627 13929
rect 23569 13889 23581 13923
rect 23615 13920 23627 13923
rect 23676 13920 23704 13948
rect 23952 13932 23980 13960
rect 23615 13892 23704 13920
rect 23615 13889 23627 13892
rect 23569 13883 23627 13889
rect 22388 13852 22416 13883
rect 23934 13880 23940 13932
rect 23992 13880 23998 13932
rect 24780 13929 24808 13960
rect 25498 13948 25504 13960
rect 25556 13948 25562 14000
rect 24029 13923 24087 13929
rect 24029 13889 24041 13923
rect 24075 13920 24087 13923
rect 24213 13923 24271 13929
rect 24075 13892 24164 13920
rect 24075 13889 24087 13892
rect 24029 13883 24087 13889
rect 22646 13852 22652 13864
rect 20680 13824 21036 13852
rect 22066 13824 22416 13852
rect 22480 13824 22652 13852
rect 20680 13812 20686 13824
rect 19334 13784 19340 13796
rect 19260 13756 19340 13784
rect 19334 13744 19340 13756
rect 19392 13744 19398 13796
rect 21726 13744 21732 13796
rect 21784 13784 21790 13796
rect 22066 13784 22094 13824
rect 21784 13756 22094 13784
rect 22281 13787 22339 13793
rect 21784 13744 21790 13756
rect 22281 13753 22293 13787
rect 22327 13784 22339 13787
rect 22480 13784 22508 13824
rect 22646 13812 22652 13824
rect 22704 13852 22710 13864
rect 24136 13852 24164 13892
rect 24213 13889 24225 13923
rect 24259 13889 24271 13923
rect 24213 13883 24271 13889
rect 24765 13923 24823 13929
rect 24765 13889 24777 13923
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 22704 13824 24164 13852
rect 24228 13852 24256 13883
rect 24854 13880 24860 13932
rect 24912 13880 24918 13932
rect 24946 13880 24952 13932
rect 25004 13920 25010 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 25004 13892 25053 13920
rect 25004 13880 25010 13892
rect 25041 13889 25053 13892
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 24673 13855 24731 13861
rect 24673 13852 24685 13855
rect 24228 13824 24685 13852
rect 22704 13812 22710 13824
rect 22327 13756 22508 13784
rect 24136 13784 24164 13824
rect 24673 13821 24685 13824
rect 24719 13852 24731 13855
rect 25222 13852 25228 13864
rect 24719 13824 25228 13852
rect 24719 13821 24731 13824
rect 24673 13815 24731 13821
rect 25222 13812 25228 13824
rect 25280 13812 25286 13864
rect 24854 13784 24860 13796
rect 24136 13756 24860 13784
rect 22327 13753 22339 13756
rect 22281 13747 22339 13753
rect 24854 13744 24860 13756
rect 24912 13744 24918 13796
rect 14550 13716 14556 13728
rect 14016 13688 14556 13716
rect 14550 13676 14556 13688
rect 14608 13676 14614 13728
rect 17310 13676 17316 13728
rect 17368 13676 17374 13728
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 19242 13716 19248 13728
rect 17644 13688 19248 13716
rect 17644 13676 17650 13688
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 21358 13676 21364 13728
rect 21416 13716 21422 13728
rect 21499 13719 21557 13725
rect 21499 13716 21511 13719
rect 21416 13688 21511 13716
rect 21416 13676 21422 13688
rect 21499 13685 21511 13688
rect 21545 13685 21557 13719
rect 21499 13679 21557 13685
rect 22646 13676 22652 13728
rect 22704 13716 22710 13728
rect 23201 13719 23259 13725
rect 23201 13716 23213 13719
rect 22704 13688 23213 13716
rect 22704 13676 22710 13688
rect 23201 13685 23213 13688
rect 23247 13685 23259 13719
rect 23201 13679 23259 13685
rect 23569 13719 23627 13725
rect 23569 13685 23581 13719
rect 23615 13716 23627 13719
rect 23842 13716 23848 13728
rect 23615 13688 23848 13716
rect 23615 13685 23627 13688
rect 23569 13679 23627 13685
rect 23842 13676 23848 13688
rect 23900 13716 23906 13728
rect 24026 13716 24032 13728
rect 23900 13688 24032 13716
rect 23900 13676 23906 13688
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 25038 13676 25044 13728
rect 25096 13676 25102 13728
rect 1104 13626 26496 13648
rect 1104 13574 4124 13626
rect 4176 13574 4188 13626
rect 4240 13574 4252 13626
rect 4304 13574 4316 13626
rect 4368 13574 4380 13626
rect 4432 13574 10472 13626
rect 10524 13574 10536 13626
rect 10588 13574 10600 13626
rect 10652 13574 10664 13626
rect 10716 13574 10728 13626
rect 10780 13574 16820 13626
rect 16872 13574 16884 13626
rect 16936 13574 16948 13626
rect 17000 13574 17012 13626
rect 17064 13574 17076 13626
rect 17128 13574 23168 13626
rect 23220 13574 23232 13626
rect 23284 13574 23296 13626
rect 23348 13574 23360 13626
rect 23412 13574 23424 13626
rect 23476 13574 26496 13626
rect 1104 13552 26496 13574
rect 2682 13472 2688 13524
rect 2740 13512 2746 13524
rect 3237 13515 3295 13521
rect 3237 13512 3249 13515
rect 2740 13484 3249 13512
rect 2740 13472 2746 13484
rect 3237 13481 3249 13484
rect 3283 13481 3295 13515
rect 3237 13475 3295 13481
rect 3510 13472 3516 13524
rect 3568 13512 3574 13524
rect 5074 13512 5080 13524
rect 3568 13484 5080 13512
rect 3568 13472 3574 13484
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 5166 13472 5172 13524
rect 5224 13512 5230 13524
rect 6362 13512 6368 13524
rect 5224 13484 6368 13512
rect 5224 13472 5230 13484
rect 6362 13472 6368 13484
rect 6420 13512 6426 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 6420 13484 7205 13512
rect 6420 13472 6426 13484
rect 7193 13481 7205 13484
rect 7239 13481 7251 13515
rect 7193 13475 7251 13481
rect 8021 13515 8079 13521
rect 8021 13481 8033 13515
rect 8067 13512 8079 13515
rect 8202 13512 8208 13524
rect 8067 13484 8208 13512
rect 8067 13481 8079 13484
rect 8021 13475 8079 13481
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 8386 13472 8392 13524
rect 8444 13512 8450 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8444 13484 8953 13512
rect 8444 13472 8450 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 14553 13515 14611 13521
rect 14553 13512 14565 13515
rect 14516 13484 14565 13512
rect 14516 13472 14522 13484
rect 14553 13481 14565 13484
rect 14599 13481 14611 13515
rect 14553 13475 14611 13481
rect 15378 13472 15384 13524
rect 15436 13472 15442 13524
rect 15488 13484 17632 13512
rect 3145 13447 3203 13453
rect 3145 13413 3157 13447
rect 3191 13444 3203 13447
rect 3602 13444 3608 13456
rect 3191 13416 3608 13444
rect 3191 13413 3203 13416
rect 3145 13407 3203 13413
rect 3602 13404 3608 13416
rect 3660 13444 3666 13456
rect 4430 13444 4436 13456
rect 3660 13416 4436 13444
rect 3660 13404 3666 13416
rect 4430 13404 4436 13416
rect 4488 13404 4494 13456
rect 8297 13447 8355 13453
rect 8297 13413 8309 13447
rect 8343 13444 8355 13447
rect 9677 13447 9735 13453
rect 9677 13444 9689 13447
rect 8343 13416 9689 13444
rect 8343 13413 8355 13416
rect 8297 13407 8355 13413
rect 9677 13413 9689 13416
rect 9723 13444 9735 13447
rect 9858 13444 9864 13456
rect 9723 13416 9864 13444
rect 9723 13413 9735 13416
rect 9677 13407 9735 13413
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13376 1734 13388
rect 4709 13379 4767 13385
rect 4709 13376 4721 13379
rect 1728 13348 4721 13376
rect 1728 13336 1734 13348
rect 4709 13345 4721 13348
rect 4755 13345 4767 13379
rect 4709 13339 4767 13345
rect 4982 13336 4988 13388
rect 5040 13336 5046 13388
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 5592 13348 6745 13376
rect 5592 13336 5598 13348
rect 6733 13345 6745 13348
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 3418 13268 3424 13320
rect 3476 13268 3482 13320
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13277 3663 13311
rect 3605 13271 3663 13277
rect 1670 13200 1676 13252
rect 1728 13200 1734 13252
rect 2958 13240 2964 13252
rect 2898 13212 2964 13240
rect 2958 13200 2964 13212
rect 3016 13240 3022 13252
rect 3510 13240 3516 13252
rect 3016 13212 3516 13240
rect 3016 13200 3022 13212
rect 3510 13200 3516 13212
rect 3568 13200 3574 13252
rect 3620 13240 3648 13271
rect 4430 13268 4436 13320
rect 4488 13268 4494 13320
rect 6748 13308 6776 13339
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 7064 13348 8248 13376
rect 7064 13336 7070 13348
rect 8220 13317 8248 13348
rect 8386 13336 8392 13388
rect 8444 13336 8450 13388
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 9766 13376 9772 13388
rect 9631 13348 9772 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 9766 13336 9772 13348
rect 9824 13376 9830 13388
rect 10318 13376 10324 13388
rect 9824 13348 10324 13376
rect 9824 13336 9830 13348
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 11296 13348 11345 13376
rect 11296 13336 11302 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 11664 13348 11713 13376
rect 11664 13336 11670 13348
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 12894 13336 12900 13388
rect 12952 13376 12958 13388
rect 13265 13379 13323 13385
rect 13265 13376 13277 13379
rect 12952 13348 13277 13376
rect 12952 13336 12958 13348
rect 13265 13345 13277 13348
rect 13311 13345 13323 13379
rect 13265 13339 13323 13345
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14642 13376 14648 13388
rect 13964 13348 14648 13376
rect 13964 13336 13970 13348
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 8205 13311 8263 13317
rect 6748 13280 7052 13308
rect 4706 13240 4712 13252
rect 3620 13212 4712 13240
rect 4706 13200 4712 13212
rect 4764 13200 4770 13252
rect 5074 13200 5080 13252
rect 5132 13240 5138 13252
rect 5132 13212 5474 13240
rect 5132 13200 5138 13212
rect 6822 13200 6828 13252
rect 6880 13200 6886 13252
rect 7024 13249 7052 13280
rect 8205 13277 8217 13311
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 8938 13308 8944 13320
rect 8527 13280 8944 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 8938 13268 8944 13280
rect 8996 13308 9002 13320
rect 9950 13308 9956 13320
rect 8996 13280 9956 13308
rect 8996 13268 9002 13280
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 10870 13308 10876 13320
rect 10643 13280 10876 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 15194 13268 15200 13320
rect 15252 13268 15258 13320
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 15488 13317 15516 13484
rect 17604 13456 17632 13484
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 18233 13515 18291 13521
rect 18233 13512 18245 13515
rect 18104 13484 18245 13512
rect 18104 13472 18110 13484
rect 18233 13481 18245 13484
rect 18279 13481 18291 13515
rect 18233 13475 18291 13481
rect 18325 13515 18383 13521
rect 18325 13481 18337 13515
rect 18371 13512 18383 13515
rect 18414 13512 18420 13524
rect 18371 13484 18420 13512
rect 18371 13481 18383 13484
rect 18325 13475 18383 13481
rect 17586 13404 17592 13456
rect 17644 13404 17650 13456
rect 15703 13379 15761 13385
rect 15703 13345 15715 13379
rect 15749 13376 15761 13379
rect 17129 13379 17187 13385
rect 15749 13348 17080 13376
rect 15749 13345 15761 13348
rect 15703 13339 15761 13345
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 15344 13280 15485 13308
rect 15344 13268 15350 13280
rect 15473 13277 15485 13280
rect 15519 13277 15531 13311
rect 17052 13308 17080 13348
rect 17129 13345 17141 13379
rect 17175 13376 17187 13379
rect 17310 13376 17316 13388
rect 17175 13348 17316 13376
rect 17175 13345 17187 13348
rect 17129 13339 17187 13345
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 17494 13336 17500 13388
rect 17552 13336 17558 13388
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17052 13280 17601 13308
rect 15473 13271 15531 13277
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 18248 13308 18276 13475
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 20438 13472 20444 13524
rect 20496 13472 20502 13524
rect 20622 13472 20628 13524
rect 20680 13472 20686 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 23845 13515 23903 13521
rect 23845 13512 23857 13515
rect 23716 13484 23857 13512
rect 23716 13472 23722 13484
rect 23845 13481 23857 13484
rect 23891 13481 23903 13515
rect 23845 13475 23903 13481
rect 24210 13472 24216 13524
rect 24268 13512 24274 13524
rect 24486 13512 24492 13524
rect 24268 13484 24492 13512
rect 24268 13472 24274 13484
rect 24486 13472 24492 13484
rect 24544 13512 24550 13524
rect 25685 13515 25743 13521
rect 25685 13512 25697 13515
rect 24544 13484 25697 13512
rect 24544 13472 24550 13484
rect 25685 13481 25697 13484
rect 25731 13481 25743 13515
rect 25685 13475 25743 13481
rect 18432 13444 18460 13472
rect 18432 13416 19840 13444
rect 18969 13379 19027 13385
rect 18969 13345 18981 13379
rect 19015 13376 19027 13379
rect 19518 13376 19524 13388
rect 19015 13348 19524 13376
rect 19015 13345 19027 13348
rect 18969 13339 19027 13345
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 19812 13317 19840 13416
rect 20640 13376 20668 13472
rect 25409 13447 25467 13453
rect 25409 13444 25421 13447
rect 24688 13416 25421 13444
rect 21358 13376 21364 13388
rect 20364 13348 20668 13376
rect 21100 13348 21364 13376
rect 20364 13317 20392 13348
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 18248 13280 19441 13308
rect 17589 13271 17647 13277
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13277 20407 13311
rect 20349 13271 20407 13277
rect 20533 13311 20591 13317
rect 20533 13277 20545 13311
rect 20579 13308 20591 13311
rect 20898 13308 20904 13320
rect 20579 13280 20904 13308
rect 20579 13277 20591 13280
rect 20533 13271 20591 13277
rect 7009 13243 7067 13249
rect 7009 13209 7021 13243
rect 7055 13209 7067 13243
rect 7009 13203 7067 13209
rect 12618 13200 12624 13252
rect 12676 13200 12682 13252
rect 13004 13212 14228 13240
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 3200 13144 3801 13172
rect 3200 13132 3206 13144
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 4982 13172 4988 13184
rect 4672 13144 4988 13172
rect 4672 13132 4678 13144
rect 4982 13132 4988 13144
rect 5040 13172 5046 13184
rect 5902 13172 5908 13184
rect 5040 13144 5908 13172
rect 5040 13132 5046 13144
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11241 13175 11299 13181
rect 11241 13172 11253 13175
rect 11204 13144 11253 13172
rect 11204 13132 11210 13144
rect 11241 13141 11253 13144
rect 11287 13172 11299 13175
rect 13004 13172 13032 13212
rect 13170 13181 13176 13184
rect 11287 13144 13032 13172
rect 13127 13175 13176 13181
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 13127 13141 13139 13175
rect 13173 13141 13176 13175
rect 13127 13135 13176 13141
rect 13170 13132 13176 13135
rect 13228 13132 13234 13184
rect 13909 13175 13967 13181
rect 13909 13141 13921 13175
rect 13955 13172 13967 13175
rect 14090 13172 14096 13184
rect 13955 13144 14096 13172
rect 13955 13141 13967 13144
rect 13909 13135 13967 13141
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 14200 13172 14228 13212
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 19521 13243 19579 13249
rect 19521 13240 19533 13243
rect 15620 13212 16146 13240
rect 17420 13212 19533 13240
rect 15620 13200 15626 13212
rect 17420 13172 17448 13212
rect 19521 13209 19533 13212
rect 19567 13209 19579 13243
rect 19521 13203 19579 13209
rect 19613 13243 19671 13249
rect 19613 13209 19625 13243
rect 19659 13240 19671 13243
rect 20364 13240 20392 13271
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 21100 13317 21128 13348
rect 21358 13336 21364 13348
rect 21416 13336 21422 13388
rect 23842 13336 23848 13388
rect 23900 13376 23906 13388
rect 23900 13348 24532 13376
rect 23900 13336 23906 13348
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 23477 13311 23535 13317
rect 23477 13277 23489 13311
rect 23523 13308 23535 13311
rect 24394 13308 24400 13320
rect 23523 13280 24400 13308
rect 23523 13277 23535 13280
rect 23477 13271 23535 13277
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 20438 13240 20444 13252
rect 19659 13212 20444 13240
rect 19659 13209 19671 13212
rect 19613 13203 19671 13209
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 24026 13200 24032 13252
rect 24084 13200 24090 13252
rect 24210 13200 24216 13252
rect 24268 13200 24274 13252
rect 14200 13144 17448 13172
rect 19242 13132 19248 13184
rect 19300 13132 19306 13184
rect 19794 13132 19800 13184
rect 19852 13172 19858 13184
rect 20993 13175 21051 13181
rect 20993 13172 21005 13175
rect 19852 13144 21005 13172
rect 19852 13132 19858 13144
rect 20993 13141 21005 13144
rect 21039 13141 21051 13175
rect 20993 13135 21051 13141
rect 23014 13132 23020 13184
rect 23072 13172 23078 13184
rect 23293 13175 23351 13181
rect 23293 13172 23305 13175
rect 23072 13144 23305 13172
rect 23072 13132 23078 13144
rect 23293 13141 23305 13144
rect 23339 13141 23351 13175
rect 23293 13135 23351 13141
rect 24118 13132 24124 13184
rect 24176 13172 24182 13184
rect 24397 13175 24455 13181
rect 24397 13172 24409 13175
rect 24176 13144 24409 13172
rect 24176 13132 24182 13144
rect 24397 13141 24409 13144
rect 24443 13141 24455 13175
rect 24504 13172 24532 13348
rect 24578 13268 24584 13320
rect 24636 13308 24642 13320
rect 24688 13308 24716 13416
rect 25409 13413 25421 13416
rect 25455 13413 25467 13447
rect 25409 13407 25467 13413
rect 25501 13447 25559 13453
rect 25501 13413 25513 13447
rect 25547 13413 25559 13447
rect 25501 13407 25559 13413
rect 24636 13280 24716 13308
rect 24636 13268 24642 13280
rect 24946 13268 24952 13320
rect 25004 13268 25010 13320
rect 25038 13268 25044 13320
rect 25096 13268 25102 13320
rect 25516 13308 25544 13407
rect 25148 13280 25544 13308
rect 24670 13200 24676 13252
rect 24728 13200 24734 13252
rect 24762 13200 24768 13252
rect 24820 13200 24826 13252
rect 24964 13240 24992 13268
rect 25148 13240 25176 13280
rect 26142 13268 26148 13320
rect 26200 13268 26206 13320
rect 24964 13212 25176 13240
rect 25222 13200 25228 13252
rect 25280 13200 25286 13252
rect 25498 13200 25504 13252
rect 25556 13240 25562 13252
rect 25664 13243 25722 13249
rect 25664 13240 25676 13243
rect 25556 13212 25676 13240
rect 25556 13200 25562 13212
rect 25664 13209 25676 13212
rect 25710 13209 25722 13243
rect 25664 13203 25722 13209
rect 25869 13243 25927 13249
rect 25869 13209 25881 13243
rect 25915 13209 25927 13243
rect 25869 13203 25927 13209
rect 25884 13172 25912 13203
rect 24504 13144 25912 13172
rect 24397 13135 24455 13141
rect 25958 13132 25964 13184
rect 26016 13132 26022 13184
rect 1104 13082 26656 13104
rect 1104 13030 7298 13082
rect 7350 13030 7362 13082
rect 7414 13030 7426 13082
rect 7478 13030 7490 13082
rect 7542 13030 7554 13082
rect 7606 13030 13646 13082
rect 13698 13030 13710 13082
rect 13762 13030 13774 13082
rect 13826 13030 13838 13082
rect 13890 13030 13902 13082
rect 13954 13030 19994 13082
rect 20046 13030 20058 13082
rect 20110 13030 20122 13082
rect 20174 13030 20186 13082
rect 20238 13030 20250 13082
rect 20302 13030 26342 13082
rect 26394 13030 26406 13082
rect 26458 13030 26470 13082
rect 26522 13030 26534 13082
rect 26586 13030 26598 13082
rect 26650 13030 26656 13082
rect 1104 13008 26656 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 2317 12971 2375 12977
rect 2317 12968 2329 12971
rect 1728 12940 2329 12968
rect 1728 12928 1734 12940
rect 2317 12937 2329 12940
rect 2363 12937 2375 12971
rect 3053 12971 3111 12977
rect 3053 12968 3065 12971
rect 2317 12931 2375 12937
rect 2746 12940 3065 12968
rect 2593 12903 2651 12909
rect 2593 12869 2605 12903
rect 2639 12900 2651 12903
rect 2746 12900 2774 12940
rect 3053 12937 3065 12940
rect 3099 12937 3111 12971
rect 3053 12931 3111 12937
rect 4890 12928 4896 12980
rect 4948 12928 4954 12980
rect 7006 12968 7012 12980
rect 6196 12940 7012 12968
rect 2866 12909 2872 12912
rect 2639 12872 2774 12900
rect 2823 12903 2872 12909
rect 2639 12869 2651 12872
rect 2593 12863 2651 12869
rect 2823 12869 2835 12903
rect 2869 12869 2872 12903
rect 2823 12863 2872 12869
rect 2866 12860 2872 12863
rect 2924 12860 2930 12912
rect 4908 12900 4936 12928
rect 5626 12900 5632 12912
rect 3344 12872 3832 12900
rect 4908 12872 5120 12900
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 2516 12628 2544 12795
rect 2682 12792 2688 12844
rect 2740 12792 2746 12844
rect 3344 12832 3372 12872
rect 3804 12841 3832 12872
rect 2792 12804 3372 12832
rect 3789 12835 3847 12841
rect 2792 12776 2820 12804
rect 3789 12801 3801 12835
rect 3835 12801 3847 12835
rect 3789 12795 3847 12801
rect 4775 12835 4833 12841
rect 4775 12801 4787 12835
rect 4821 12832 4833 12835
rect 4821 12801 4844 12832
rect 4775 12795 4844 12801
rect 2774 12724 2780 12776
rect 2832 12724 2838 12776
rect 2961 12767 3019 12773
rect 2961 12733 2973 12767
rect 3007 12764 3019 12767
rect 3142 12764 3148 12776
rect 3007 12736 3148 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 3234 12724 3240 12776
rect 3292 12724 3298 12776
rect 3326 12724 3332 12776
rect 3384 12724 3390 12776
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 3050 12656 3056 12708
rect 3108 12696 3114 12708
rect 3436 12696 3464 12727
rect 3510 12724 3516 12776
rect 3568 12724 3574 12776
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 4816 12764 4844 12795
rect 4890 12792 4896 12844
rect 4948 12792 4954 12844
rect 4982 12792 4988 12844
rect 5040 12792 5046 12844
rect 5092 12841 5120 12872
rect 5184 12872 5632 12900
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5184 12764 5212 12872
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12832 5595 12835
rect 6196 12832 6224 12940
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 7561 12971 7619 12977
rect 7561 12968 7573 12971
rect 7156 12940 7573 12968
rect 7156 12928 7162 12940
rect 7561 12937 7573 12940
rect 7607 12937 7619 12971
rect 7561 12931 7619 12937
rect 9033 12971 9091 12977
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 9122 12968 9128 12980
rect 9079 12940 9128 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9309 12971 9367 12977
rect 9309 12937 9321 12971
rect 9355 12968 9367 12971
rect 9766 12968 9772 12980
rect 9355 12940 9772 12968
rect 9355 12937 9367 12940
rect 9309 12931 9367 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 15427 12971 15485 12977
rect 15427 12968 15439 12971
rect 14608 12940 15439 12968
rect 14608 12928 14614 12940
rect 15427 12937 15439 12940
rect 15473 12937 15485 12971
rect 17954 12968 17960 12980
rect 15427 12931 15485 12937
rect 15580 12940 17960 12968
rect 15580 12912 15608 12940
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 9214 12900 9220 12912
rect 6328 12872 9220 12900
rect 6328 12860 6334 12872
rect 9214 12860 9220 12872
rect 9272 12860 9278 12912
rect 12434 12860 12440 12912
rect 12492 12860 12498 12912
rect 15562 12900 15568 12912
rect 15042 12872 15568 12900
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 17402 12900 17408 12912
rect 16868 12872 17408 12900
rect 5583 12804 6224 12832
rect 6365 12835 6423 12841
rect 5583 12801 5595 12804
rect 5537 12795 5595 12801
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 4816 12736 5212 12764
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12733 5503 12767
rect 5445 12727 5503 12733
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 6380 12764 6408 12795
rect 6638 12792 6644 12844
rect 6696 12792 6702 12844
rect 8846 12792 8852 12844
rect 8904 12792 8910 12844
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12801 9183 12835
rect 9125 12795 9183 12801
rect 5951 12736 6408 12764
rect 6457 12767 6515 12773
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 6457 12733 6469 12767
rect 6503 12733 6515 12767
rect 6457 12727 6515 12733
rect 3881 12699 3939 12705
rect 3881 12696 3893 12699
rect 3108 12668 3464 12696
rect 3528 12668 3893 12696
rect 3108 12656 3114 12668
rect 3528 12628 3556 12668
rect 3881 12665 3893 12668
rect 3927 12665 3939 12699
rect 3881 12659 3939 12665
rect 4430 12656 4436 12708
rect 4488 12696 4494 12708
rect 5460 12696 5488 12727
rect 5534 12696 5540 12708
rect 4488 12668 5540 12696
rect 4488 12656 4494 12668
rect 5534 12656 5540 12668
rect 5592 12656 5598 12708
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 6472 12696 6500 12727
rect 8110 12724 8116 12776
rect 8168 12724 8174 12776
rect 8864 12764 8892 12792
rect 9140 12764 9168 12795
rect 9674 12792 9680 12844
rect 9732 12792 9738 12844
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12832 14059 12835
rect 14090 12832 14096 12844
rect 14047 12804 14096 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 16868 12841 16896 12872
rect 17402 12860 17408 12872
rect 17460 12860 17466 12912
rect 17512 12900 17540 12940
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 19242 12928 19248 12980
rect 19300 12928 19306 12980
rect 23842 12928 23848 12980
rect 23900 12968 23906 12980
rect 23900 12940 24072 12968
rect 23900 12928 23906 12940
rect 17512 12872 17618 12900
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 8864 12736 9168 12764
rect 10042 12724 10048 12776
rect 10100 12764 10106 12776
rect 10781 12767 10839 12773
rect 10781 12764 10793 12767
rect 10100 12736 10793 12764
rect 10100 12724 10106 12736
rect 10781 12733 10793 12736
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 11112 12736 11621 12764
rect 11112 12724 11118 12736
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 6052 12668 6500 12696
rect 6052 12656 6058 12668
rect 2516 12600 3556 12628
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5626 12628 5632 12640
rect 5307 12600 5632 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 6362 12588 6368 12640
rect 6420 12588 6426 12640
rect 6822 12588 6828 12640
rect 6880 12588 6886 12640
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 10134 12628 10140 12640
rect 8996 12600 10140 12628
rect 8996 12588 9002 12600
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 11624 12628 11652 12727
rect 11882 12724 11888 12776
rect 11940 12724 11946 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 12912 12736 13645 12764
rect 12912 12628 12940 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 19260 12764 19288 12928
rect 21545 12903 21603 12909
rect 21545 12900 21557 12903
rect 20180 12872 21557 12900
rect 20180 12841 20208 12872
rect 21545 12869 21557 12872
rect 21591 12869 21603 12903
rect 21545 12863 21603 12869
rect 23934 12860 23940 12912
rect 23992 12860 23998 12912
rect 24044 12909 24072 12940
rect 24670 12928 24676 12980
rect 24728 12928 24734 12980
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 25317 12971 25375 12977
rect 25317 12968 25329 12971
rect 24820 12940 25329 12968
rect 24820 12928 24826 12940
rect 25317 12937 25329 12940
rect 25363 12937 25375 12971
rect 25317 12931 25375 12937
rect 24029 12903 24087 12909
rect 24029 12869 24041 12903
rect 24075 12869 24087 12903
rect 24029 12863 24087 12869
rect 24167 12903 24225 12909
rect 24167 12869 24179 12903
rect 24213 12900 24225 12903
rect 24578 12900 24584 12912
rect 24213 12872 24584 12900
rect 24213 12869 24225 12872
rect 24167 12863 24225 12869
rect 24578 12860 24584 12872
rect 24636 12860 24642 12912
rect 24688 12900 24716 12928
rect 25501 12903 25559 12909
rect 25501 12900 25513 12903
rect 24688 12872 25513 12900
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 20438 12792 20444 12844
rect 20496 12792 20502 12844
rect 20898 12792 20904 12844
rect 20956 12792 20962 12844
rect 21177 12835 21235 12841
rect 21177 12801 21189 12835
rect 21223 12801 21235 12835
rect 21177 12795 21235 12801
rect 21361 12835 21419 12841
rect 21361 12801 21373 12835
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 17175 12736 19288 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 19426 12724 19432 12776
rect 19484 12724 19490 12776
rect 20625 12767 20683 12773
rect 20625 12733 20637 12767
rect 20671 12764 20683 12767
rect 20806 12764 20812 12776
rect 20671 12736 20812 12764
rect 20671 12733 20683 12736
rect 20625 12727 20683 12733
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 18601 12699 18659 12705
rect 18601 12665 18613 12699
rect 18647 12696 18659 12699
rect 19444 12696 19472 12724
rect 18647 12668 19472 12696
rect 21192 12696 21220 12795
rect 21376 12764 21404 12795
rect 21450 12792 21456 12844
rect 21508 12792 21514 12844
rect 21637 12835 21695 12841
rect 21637 12801 21649 12835
rect 21683 12832 21695 12835
rect 21726 12832 21732 12844
rect 21683 12804 21732 12832
rect 21683 12801 21695 12804
rect 21637 12795 21695 12801
rect 21726 12792 21732 12804
rect 21784 12792 21790 12844
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 22152 12804 23213 12832
rect 22152 12792 22158 12804
rect 23201 12801 23213 12804
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23566 12792 23572 12844
rect 23624 12792 23630 12844
rect 23845 12835 23903 12841
rect 23845 12801 23857 12835
rect 23891 12832 23903 12835
rect 25038 12832 25044 12844
rect 23891 12804 25044 12832
rect 23891 12801 23903 12804
rect 23845 12795 23903 12801
rect 25038 12792 25044 12804
rect 25096 12792 25102 12844
rect 25130 12792 25136 12844
rect 25188 12832 25194 12844
rect 25424 12841 25452 12872
rect 25501 12869 25513 12872
rect 25547 12869 25559 12903
rect 25501 12863 25559 12869
rect 25225 12835 25283 12841
rect 25225 12832 25237 12835
rect 25188 12804 25237 12832
rect 25188 12792 25194 12804
rect 25225 12801 25237 12804
rect 25271 12801 25283 12835
rect 25225 12795 25283 12801
rect 25409 12835 25467 12841
rect 25409 12801 25421 12835
rect 25455 12832 25467 12835
rect 26050 12832 26056 12844
rect 25455 12804 25489 12832
rect 25608 12804 26056 12832
rect 25455 12801 25467 12804
rect 25409 12795 25467 12801
rect 21542 12764 21548 12776
rect 21376 12736 21548 12764
rect 21542 12724 21548 12736
rect 21600 12724 21606 12776
rect 24026 12724 24032 12776
rect 24084 12724 24090 12776
rect 24305 12767 24363 12773
rect 24305 12733 24317 12767
rect 24351 12764 24363 12767
rect 24397 12767 24455 12773
rect 24397 12764 24409 12767
rect 24351 12736 24409 12764
rect 24351 12733 24363 12736
rect 24305 12727 24363 12733
rect 24397 12733 24409 12736
rect 24443 12733 24455 12767
rect 24397 12727 24455 12733
rect 24486 12724 24492 12776
rect 24544 12764 24550 12776
rect 24949 12767 25007 12773
rect 24949 12764 24961 12767
rect 24544 12736 24961 12764
rect 24544 12724 24550 12736
rect 24949 12733 24961 12736
rect 24995 12733 25007 12767
rect 25608 12764 25636 12804
rect 26050 12792 26056 12804
rect 26108 12832 26114 12844
rect 26145 12835 26203 12841
rect 26145 12832 26157 12835
rect 26108 12804 26157 12832
rect 26108 12792 26114 12804
rect 26145 12801 26157 12804
rect 26191 12801 26203 12835
rect 26145 12795 26203 12801
rect 24949 12727 25007 12733
rect 25424 12736 25636 12764
rect 22646 12696 22652 12708
rect 21192 12668 22652 12696
rect 18647 12665 18659 12668
rect 18601 12659 18659 12665
rect 22646 12656 22652 12668
rect 22704 12656 22710 12708
rect 24044 12696 24072 12724
rect 25424 12696 25452 12736
rect 24044 12668 25452 12696
rect 11624 12600 12940 12628
rect 12986 12588 12992 12640
rect 13044 12628 13050 12640
rect 13357 12631 13415 12637
rect 13357 12628 13369 12631
rect 13044 12600 13369 12628
rect 13044 12588 13050 12600
rect 13357 12597 13369 12600
rect 13403 12597 13415 12631
rect 13357 12591 13415 12597
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 20714 12588 20720 12640
rect 20772 12588 20778 12640
rect 21910 12588 21916 12640
rect 21968 12588 21974 12640
rect 23658 12588 23664 12640
rect 23716 12588 23722 12640
rect 1104 12538 26496 12560
rect 1104 12486 4124 12538
rect 4176 12486 4188 12538
rect 4240 12486 4252 12538
rect 4304 12486 4316 12538
rect 4368 12486 4380 12538
rect 4432 12486 10472 12538
rect 10524 12486 10536 12538
rect 10588 12486 10600 12538
rect 10652 12486 10664 12538
rect 10716 12486 10728 12538
rect 10780 12486 16820 12538
rect 16872 12486 16884 12538
rect 16936 12486 16948 12538
rect 17000 12486 17012 12538
rect 17064 12486 17076 12538
rect 17128 12486 23168 12538
rect 23220 12486 23232 12538
rect 23284 12486 23296 12538
rect 23348 12486 23360 12538
rect 23412 12486 23424 12538
rect 23476 12486 26496 12538
rect 1104 12464 26496 12486
rect 4982 12384 4988 12436
rect 5040 12384 5046 12436
rect 6270 12384 6276 12436
rect 6328 12384 6334 12436
rect 6638 12424 6644 12436
rect 6380 12396 6644 12424
rect 5261 12359 5319 12365
rect 5261 12325 5273 12359
rect 5307 12356 5319 12359
rect 6380 12356 6408 12396
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 11940 12396 12265 12424
rect 11940 12384 11946 12396
rect 12253 12393 12265 12396
rect 12299 12393 12311 12427
rect 12253 12387 12311 12393
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12424 13783 12427
rect 14274 12424 14280 12436
rect 13771 12396 14280 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 15194 12424 15200 12436
rect 14599 12396 15200 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 19242 12384 19248 12436
rect 19300 12424 19306 12436
rect 20898 12424 20904 12436
rect 19300 12396 20904 12424
rect 19300 12384 19306 12396
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 23842 12384 23848 12436
rect 23900 12424 23906 12436
rect 24213 12427 24271 12433
rect 24213 12424 24225 12427
rect 23900 12396 24225 12424
rect 23900 12384 23906 12396
rect 24213 12393 24225 12396
rect 24259 12393 24271 12427
rect 24213 12387 24271 12393
rect 26050 12384 26056 12436
rect 26108 12424 26114 12436
rect 26145 12427 26203 12433
rect 26145 12424 26157 12427
rect 26108 12396 26157 12424
rect 26108 12384 26114 12396
rect 26145 12393 26157 12396
rect 26191 12393 26203 12427
rect 26145 12387 26203 12393
rect 5307 12328 6408 12356
rect 6457 12359 6515 12365
rect 5307 12325 5319 12328
rect 5261 12319 5319 12325
rect 6457 12325 6469 12359
rect 6503 12356 6515 12359
rect 7742 12356 7748 12368
rect 6503 12328 7748 12356
rect 6503 12325 6515 12328
rect 6457 12319 6515 12325
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 11572 12328 14964 12356
rect 11572 12316 11578 12328
rect 3973 12291 4031 12297
rect 3973 12257 3985 12291
rect 4019 12288 4031 12291
rect 4614 12288 4620 12300
rect 4019 12260 4620 12288
rect 4019 12257 4031 12260
rect 3973 12251 4031 12257
rect 4614 12248 4620 12260
rect 4672 12288 4678 12300
rect 4985 12291 5043 12297
rect 4985 12288 4997 12291
rect 4672 12260 4997 12288
rect 4672 12248 4678 12260
rect 4985 12257 4997 12260
rect 5031 12257 5043 12291
rect 9217 12291 9275 12297
rect 4985 12251 5043 12257
rect 8128 12260 8708 12288
rect 8128 12232 8156 12260
rect 3878 12180 3884 12232
rect 3936 12180 3942 12232
rect 4522 12180 4528 12232
rect 4580 12220 4586 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4580 12192 4721 12220
rect 4580 12180 4586 12192
rect 4709 12189 4721 12192
rect 4755 12220 4767 12223
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 4755 12192 5365 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 5353 12189 5365 12192
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12220 5779 12223
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 5767 12192 6101 12220
rect 5767 12189 5779 12192
rect 5721 12183 5779 12189
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 5813 12155 5871 12161
rect 5813 12152 5825 12155
rect 5684 12124 5825 12152
rect 5684 12112 5690 12124
rect 5813 12121 5825 12124
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 6288 12152 6316 12183
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 6822 12220 6828 12232
rect 6604 12192 6828 12220
rect 6604 12180 6610 12192
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 6932 12152 6960 12183
rect 7098 12180 7104 12232
rect 7156 12180 7162 12232
rect 8110 12180 8116 12232
rect 8168 12180 8174 12232
rect 8680 12229 8708 12260
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 9490 12288 9496 12300
rect 9263 12260 9496 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 9490 12248 9496 12260
rect 9548 12288 9554 12300
rect 11054 12288 11060 12300
rect 9548 12260 11060 12288
rect 9548 12248 9554 12260
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12189 8723 12223
rect 8665 12183 8723 12189
rect 6052 12124 6316 12152
rect 6748 12124 6960 12152
rect 8496 12152 8524 12183
rect 9582 12180 9588 12232
rect 9640 12180 9646 12232
rect 12452 12229 12480 12328
rect 12621 12291 12679 12297
rect 12621 12257 12633 12291
rect 12667 12288 12679 12291
rect 12805 12291 12863 12297
rect 12805 12288 12817 12291
rect 12667 12260 12817 12288
rect 12667 12257 12679 12260
rect 12621 12251 12679 12257
rect 12805 12257 12817 12260
rect 12851 12257 12863 12291
rect 12805 12251 12863 12257
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 14608 12260 14872 12288
rect 14608 12248 14614 12260
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12189 11759 12223
rect 11701 12183 11759 12189
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 8496 12124 8800 12152
rect 6052 12112 6058 12124
rect 6748 12096 6776 12124
rect 8772 12096 8800 12124
rect 9306 12112 9312 12164
rect 9364 12112 9370 12164
rect 11011 12155 11069 12161
rect 9876 12124 9982 12152
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 6730 12084 6736 12096
rect 3476 12056 6736 12084
rect 3476 12044 3482 12056
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7006 12044 7012 12096
rect 7064 12044 7070 12096
rect 8570 12044 8576 12096
rect 8628 12044 8634 12096
rect 8754 12044 8760 12096
rect 8812 12044 8818 12096
rect 9324 12084 9352 12112
rect 9876 12084 9904 12124
rect 11011 12121 11023 12155
rect 11057 12152 11069 12155
rect 11238 12152 11244 12164
rect 11057 12124 11244 12152
rect 11057 12121 11069 12124
rect 11011 12115 11069 12121
rect 11238 12112 11244 12124
rect 11296 12152 11302 12164
rect 11716 12152 11744 12183
rect 12710 12180 12716 12232
rect 12768 12180 12774 12232
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 13170 12180 13176 12232
rect 13228 12180 13234 12232
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 14844 12229 14872 12260
rect 14936 12229 14964 12328
rect 15654 12316 15660 12368
rect 15712 12356 15718 12368
rect 20438 12356 20444 12368
rect 15712 12328 20444 12356
rect 15712 12316 15718 12328
rect 20438 12316 20444 12328
rect 20496 12316 20502 12368
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19392 12260 19441 12288
rect 19392 12248 19398 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 19886 12248 19892 12300
rect 19944 12288 19950 12300
rect 20533 12291 20591 12297
rect 20533 12288 20545 12291
rect 19944 12260 20545 12288
rect 19944 12248 19950 12260
rect 20533 12257 20545 12260
rect 20579 12288 20591 12291
rect 20898 12288 20904 12300
rect 20579 12260 20904 12288
rect 20579 12257 20591 12260
rect 20533 12251 20591 12257
rect 20898 12248 20904 12260
rect 20956 12288 20962 12300
rect 22465 12291 22523 12297
rect 22465 12288 22477 12291
rect 20956 12260 22477 12288
rect 20956 12248 20962 12260
rect 22465 12257 22477 12260
rect 22511 12288 22523 12291
rect 22738 12288 22744 12300
rect 22511 12260 22744 12288
rect 22511 12257 22523 12260
rect 22465 12251 22523 12257
rect 22738 12248 22744 12260
rect 22796 12288 22802 12300
rect 24302 12288 24308 12300
rect 22796 12260 24308 12288
rect 22796 12248 22802 12260
rect 24302 12248 24308 12260
rect 24360 12288 24366 12300
rect 24397 12291 24455 12297
rect 24397 12288 24409 12291
rect 24360 12260 24409 12288
rect 24360 12248 24366 12260
rect 24397 12257 24409 12260
rect 24443 12257 24455 12291
rect 24397 12251 24455 12257
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 14737 12223 14795 12229
rect 13771 12192 14228 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14200 12164 14228 12192
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12220 15163 12223
rect 15470 12220 15476 12232
rect 15151 12192 15476 12220
rect 15151 12189 15163 12192
rect 15105 12183 15163 12189
rect 11296 12124 11744 12152
rect 11296 12112 11302 12124
rect 14182 12112 14188 12164
rect 14240 12112 14246 12164
rect 14752 12152 14780 12183
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 16390 12180 16396 12232
rect 16448 12220 16454 12232
rect 19242 12220 19248 12232
rect 16448 12192 19248 12220
rect 16448 12180 16454 12192
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19518 12180 19524 12232
rect 19576 12180 19582 12232
rect 19610 12180 19616 12232
rect 19668 12180 19674 12232
rect 19702 12180 19708 12232
rect 19760 12180 19766 12232
rect 19794 12180 19800 12232
rect 19852 12220 19858 12232
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 19852 12192 20269 12220
rect 19852 12180 19858 12192
rect 20257 12189 20269 12192
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 15194 12152 15200 12164
rect 14752 12124 15200 12152
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 19812 12152 19840 12180
rect 15580 12124 19840 12152
rect 15580 12096 15608 12124
rect 20456 12096 20484 12183
rect 21818 12180 21824 12232
rect 21876 12220 21882 12232
rect 21876 12192 22508 12220
rect 21876 12180 21882 12192
rect 20806 12112 20812 12164
rect 20864 12112 20870 12164
rect 21542 12112 21548 12164
rect 21600 12112 21606 12164
rect 9324 12056 9904 12084
rect 10502 12044 10508 12096
rect 10560 12084 10566 12096
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 10560 12056 11161 12084
rect 10560 12044 10566 12056
rect 11149 12053 11161 12056
rect 11195 12053 11207 12087
rect 11149 12047 11207 12053
rect 13909 12087 13967 12093
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14458 12084 14464 12096
rect 13955 12056 14464 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 15562 12044 15568 12096
rect 15620 12044 15626 12096
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 19334 12084 19340 12096
rect 16356 12056 19340 12084
rect 16356 12044 16362 12056
rect 19334 12044 19340 12056
rect 19392 12084 19398 12096
rect 19702 12084 19708 12096
rect 19392 12056 19708 12084
rect 19392 12044 19398 12056
rect 19702 12044 19708 12056
rect 19760 12044 19766 12096
rect 19886 12044 19892 12096
rect 19944 12044 19950 12096
rect 20254 12044 20260 12096
rect 20312 12084 20318 12096
rect 20349 12087 20407 12093
rect 20349 12084 20361 12087
rect 20312 12056 20361 12084
rect 20312 12044 20318 12056
rect 20349 12053 20361 12056
rect 20395 12053 20407 12087
rect 20349 12047 20407 12053
rect 20438 12044 20444 12096
rect 20496 12044 20502 12096
rect 21174 12044 21180 12096
rect 21232 12084 21238 12096
rect 21726 12084 21732 12096
rect 21232 12056 21732 12084
rect 21232 12044 21238 12056
rect 21726 12044 21732 12056
rect 21784 12084 21790 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 21784 12056 22293 12084
rect 21784 12044 21790 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 22480 12084 22508 12192
rect 22741 12155 22799 12161
rect 22741 12121 22753 12155
rect 22787 12152 22799 12155
rect 23014 12152 23020 12164
rect 22787 12124 23020 12152
rect 22787 12121 22799 12124
rect 22741 12115 22799 12121
rect 23014 12112 23020 12124
rect 23072 12112 23078 12164
rect 23750 12112 23756 12164
rect 23808 12112 23814 12164
rect 24118 12112 24124 12164
rect 24176 12152 24182 12164
rect 24673 12155 24731 12161
rect 24673 12152 24685 12155
rect 24176 12124 24685 12152
rect 24176 12112 24182 12124
rect 24673 12121 24685 12124
rect 24719 12121 24731 12155
rect 24673 12115 24731 12121
rect 24780 12124 25162 12152
rect 23474 12084 23480 12096
rect 22480 12056 23480 12084
rect 22281 12047 22339 12053
rect 23474 12044 23480 12056
rect 23532 12084 23538 12096
rect 24780 12084 24808 12124
rect 23532 12056 24808 12084
rect 23532 12044 23538 12056
rect 1104 11994 26656 12016
rect 1104 11942 7298 11994
rect 7350 11942 7362 11994
rect 7414 11942 7426 11994
rect 7478 11942 7490 11994
rect 7542 11942 7554 11994
rect 7606 11942 13646 11994
rect 13698 11942 13710 11994
rect 13762 11942 13774 11994
rect 13826 11942 13838 11994
rect 13890 11942 13902 11994
rect 13954 11942 19994 11994
rect 20046 11942 20058 11994
rect 20110 11942 20122 11994
rect 20174 11942 20186 11994
rect 20238 11942 20250 11994
rect 20302 11942 26342 11994
rect 26394 11942 26406 11994
rect 26458 11942 26470 11994
rect 26522 11942 26534 11994
rect 26586 11942 26598 11994
rect 26650 11942 26656 11994
rect 1104 11920 26656 11942
rect 3510 11880 3516 11892
rect 2792 11852 3516 11880
rect 2792 11753 2820 11852
rect 3510 11840 3516 11852
rect 3568 11880 3574 11892
rect 3568 11852 3832 11880
rect 3568 11840 3574 11852
rect 2866 11772 2872 11824
rect 2924 11772 2930 11824
rect 3804 11812 3832 11852
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 4856 11852 5856 11880
rect 4856 11840 4862 11852
rect 3973 11815 4031 11821
rect 3973 11812 3985 11815
rect 3804 11784 3985 11812
rect 3973 11781 3985 11784
rect 4019 11781 4031 11815
rect 3973 11775 4031 11781
rect 4157 11815 4215 11821
rect 4157 11781 4169 11815
rect 4203 11812 4215 11815
rect 5828 11812 5856 11852
rect 7098 11840 7104 11892
rect 7156 11880 7162 11892
rect 9217 11883 9275 11889
rect 7156 11852 7328 11880
rect 7156 11840 7162 11852
rect 7300 11812 7328 11852
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 9306 11880 9312 11892
rect 9263 11852 9312 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 9640 11852 10057 11880
rect 9640 11840 9646 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10045 11843 10103 11849
rect 10502 11840 10508 11892
rect 10560 11840 10566 11892
rect 11149 11883 11207 11889
rect 11149 11849 11161 11883
rect 11195 11880 11207 11883
rect 11238 11880 11244 11892
rect 11195 11852 11244 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12768 11852 12909 11880
rect 12768 11840 12774 11852
rect 12897 11849 12909 11852
rect 12943 11849 12955 11883
rect 12897 11843 12955 11849
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 15470 11880 15476 11892
rect 13044 11852 15476 11880
rect 13044 11840 13050 11852
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15654 11840 15660 11892
rect 15712 11840 15718 11892
rect 17773 11883 17831 11889
rect 17773 11849 17785 11883
rect 17819 11880 17831 11883
rect 18138 11880 18144 11892
rect 17819 11852 18144 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 18138 11840 18144 11852
rect 18196 11880 18202 11892
rect 18196 11852 18828 11880
rect 18196 11840 18202 11852
rect 8846 11812 8852 11824
rect 4203 11784 5304 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 5276 11756 5304 11784
rect 5828 11784 6684 11812
rect 7300 11784 7406 11812
rect 8496 11784 8852 11812
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 3237 11747 3295 11753
rect 3237 11744 3249 11747
rect 3191 11716 3249 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3237 11713 3249 11716
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 2976 11608 3004 11707
rect 3878 11704 3884 11756
rect 3936 11704 3942 11756
rect 4430 11704 4436 11756
rect 4488 11704 4494 11756
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4764 11716 4813 11744
rect 4764 11704 4770 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 4816 11676 4844 11707
rect 4982 11704 4988 11756
rect 5040 11704 5046 11756
rect 5258 11704 5264 11756
rect 5316 11704 5322 11756
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5552 11676 5580 11707
rect 5718 11704 5724 11756
rect 5776 11704 5782 11756
rect 5828 11753 5856 11784
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11744 6055 11747
rect 6546 11744 6552 11756
rect 6043 11716 6552 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 6656 11744 6684 11784
rect 8496 11756 8524 11784
rect 8846 11772 8852 11784
rect 8904 11812 8910 11824
rect 8904 11784 9628 11812
rect 8904 11772 8910 11784
rect 6656 11716 6960 11744
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 4816 11648 5917 11676
rect 5905 11645 5917 11648
rect 5951 11676 5963 11679
rect 6362 11676 6368 11688
rect 5951 11648 6368 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 6822 11676 6828 11688
rect 6687 11648 6828 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 6932 11676 6960 11716
rect 7006 11704 7012 11756
rect 7064 11704 7070 11756
rect 8478 11704 8484 11756
rect 8536 11704 8542 11756
rect 8938 11704 8944 11756
rect 8996 11704 9002 11756
rect 9600 11753 9628 11784
rect 9674 11772 9680 11824
rect 9732 11772 9738 11824
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9766 11704 9772 11756
rect 9824 11704 9830 11756
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10520 11744 10548 11840
rect 13004 11812 13032 11840
rect 14182 11812 14188 11824
rect 12820 11784 13032 11812
rect 14016 11784 14188 11812
rect 9999 11716 10548 11744
rect 10965 11747 11023 11753
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10965 11713 10977 11747
rect 11011 11744 11023 11747
rect 11146 11744 11152 11756
rect 11011 11716 11152 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 12820 11753 12848 11784
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11744 13047 11747
rect 13170 11744 13176 11756
rect 13035 11716 13176 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 8110 11676 8116 11688
rect 6932 11648 8116 11676
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 8956 11676 8984 11704
rect 10042 11676 10048 11688
rect 8312 11648 8984 11676
rect 9416 11648 10048 11676
rect 3050 11608 3056 11620
rect 2976 11580 3056 11608
rect 3050 11568 3056 11580
rect 3108 11608 3114 11620
rect 4341 11611 4399 11617
rect 4341 11608 4353 11611
rect 3108 11580 4353 11608
rect 3108 11568 3114 11580
rect 4341 11577 4353 11580
rect 4387 11577 4399 11611
rect 4341 11571 4399 11577
rect 4430 11568 4436 11620
rect 4488 11608 4494 11620
rect 4488 11580 6684 11608
rect 4488 11568 4494 11580
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2593 11543 2651 11549
rect 2593 11540 2605 11543
rect 2188 11512 2605 11540
rect 2188 11500 2194 11512
rect 2593 11509 2605 11512
rect 2639 11509 2651 11543
rect 2593 11503 2651 11509
rect 3142 11500 3148 11552
rect 3200 11540 3206 11552
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 3200 11512 4629 11540
rect 3200 11500 3206 11512
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 4985 11543 5043 11549
rect 4985 11509 4997 11543
rect 5031 11540 5043 11543
rect 5074 11540 5080 11552
rect 5031 11512 5080 11540
rect 5031 11509 5043 11512
rect 4985 11503 5043 11509
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5316 11512 5365 11540
rect 5316 11500 5322 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 6656 11540 6684 11580
rect 8312 11540 8340 11648
rect 9214 11568 9220 11620
rect 9272 11568 9278 11620
rect 9416 11617 9444 11648
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10735 11648 10793 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 9401 11611 9459 11617
rect 9401 11577 9413 11611
rect 9447 11577 9459 11611
rect 11256 11608 11284 11707
rect 13170 11704 13176 11716
rect 13228 11744 13234 11756
rect 13538 11744 13544 11756
rect 13228 11716 13544 11744
rect 13228 11704 13234 11716
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 14016 11753 14044 11784
rect 14182 11772 14188 11784
rect 14240 11812 14246 11824
rect 14240 11784 14320 11812
rect 14240 11772 14246 11784
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 9401 11571 9459 11577
rect 9646 11580 11284 11608
rect 13832 11608 13860 11707
rect 14090 11704 14096 11756
rect 14148 11704 14154 11756
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11645 14243 11679
rect 14185 11639 14243 11645
rect 14090 11608 14096 11620
rect 13832 11580 14096 11608
rect 6656 11512 8340 11540
rect 8435 11543 8493 11549
rect 5353 11503 5411 11509
rect 8435 11509 8447 11543
rect 8481 11540 8493 11543
rect 8846 11540 8852 11552
rect 8481 11512 8852 11540
rect 8481 11509 8493 11512
rect 8435 11503 8493 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9232 11540 9260 11568
rect 9646 11540 9674 11580
rect 9232 11512 9674 11540
rect 11256 11540 11284 11580
rect 14090 11568 14096 11580
rect 14148 11568 14154 11620
rect 14200 11552 14228 11639
rect 14292 11608 14320 11784
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 15672 11812 15700 11840
rect 16390 11812 16396 11824
rect 14516 11784 14872 11812
rect 14516 11772 14522 11784
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 14642 11744 14648 11756
rect 14415 11716 14648 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 14844 11753 14872 11784
rect 15212 11784 15700 11812
rect 15764 11784 16396 11812
rect 14829 11747 14887 11753
rect 14829 11713 14841 11747
rect 14875 11713 14887 11747
rect 14829 11707 14887 11713
rect 14918 11704 14924 11756
rect 14976 11704 14982 11756
rect 15212 11753 15240 11784
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15028 11676 15056 11707
rect 15286 11704 15292 11756
rect 15344 11704 15350 11756
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15396 11676 15424 11707
rect 15562 11704 15568 11756
rect 15620 11704 15626 11756
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11744 15715 11747
rect 15764 11744 15792 11784
rect 16390 11772 16396 11784
rect 16448 11772 16454 11824
rect 17402 11772 17408 11824
rect 17460 11812 17466 11824
rect 18690 11812 18696 11824
rect 17460 11784 18696 11812
rect 17460 11772 17466 11784
rect 18690 11772 18696 11784
rect 18748 11772 18754 11824
rect 18800 11812 18828 11852
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 20073 11883 20131 11889
rect 20073 11880 20085 11883
rect 19576 11852 20085 11880
rect 19576 11840 19582 11852
rect 20073 11849 20085 11852
rect 20119 11849 20131 11883
rect 20073 11843 20131 11849
rect 20346 11840 20352 11892
rect 20404 11880 20410 11892
rect 20533 11883 20591 11889
rect 20533 11880 20545 11883
rect 20404 11852 20545 11880
rect 20404 11840 20410 11852
rect 20533 11849 20545 11852
rect 20579 11849 20591 11883
rect 20533 11843 20591 11849
rect 22738 11840 22744 11892
rect 22796 11840 22802 11892
rect 24397 11883 24455 11889
rect 24397 11849 24409 11883
rect 24443 11880 24455 11883
rect 24486 11880 24492 11892
rect 24443 11852 24492 11880
rect 24443 11849 24455 11852
rect 24397 11843 24455 11849
rect 24486 11840 24492 11852
rect 24544 11840 24550 11892
rect 20441 11815 20499 11821
rect 18800 11784 19932 11812
rect 15930 11753 15936 11756
rect 15703 11716 15792 11744
rect 15835 11747 15893 11753
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 15835 11713 15847 11747
rect 15881 11713 15893 11747
rect 15835 11707 15893 11713
rect 15923 11747 15936 11753
rect 15923 11713 15935 11747
rect 15988 11744 15994 11756
rect 16117 11747 16175 11753
rect 15988 11716 16023 11744
rect 15923 11707 15936 11713
rect 15672 11676 15700 11707
rect 15028 11648 15700 11676
rect 15856 11608 15884 11707
rect 15930 11704 15936 11707
rect 15988 11704 15994 11716
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16163 11716 16528 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16500 11688 16528 11716
rect 17218 11704 17224 11756
rect 17276 11744 17282 11756
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 17276 11716 17693 11744
rect 17276 11704 17282 11716
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 16482 11636 16488 11688
rect 16540 11636 16546 11688
rect 17880 11676 17908 11707
rect 17954 11704 17960 11756
rect 18012 11704 18018 11756
rect 19610 11704 19616 11756
rect 19668 11704 19674 11756
rect 19702 11704 19708 11756
rect 19760 11704 19766 11756
rect 19904 11753 19932 11784
rect 20441 11781 20453 11815
rect 20487 11812 20499 11815
rect 22756 11812 22784 11840
rect 20487 11784 22094 11812
rect 20487 11781 20499 11784
rect 20441 11775 20499 11781
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 21174 11704 21180 11756
rect 21232 11704 21238 11756
rect 18046 11676 18052 11688
rect 17880 11648 18052 11676
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18506 11636 18512 11688
rect 18564 11676 18570 11688
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 18564 11648 20729 11676
rect 18564 11636 18570 11648
rect 20717 11645 20729 11648
rect 20763 11676 20775 11679
rect 20763 11648 21312 11676
rect 20763 11645 20775 11648
rect 20717 11639 20775 11645
rect 20438 11608 20444 11620
rect 14292 11580 15332 11608
rect 15856 11580 20444 11608
rect 15304 11552 15332 11580
rect 20438 11568 20444 11580
rect 20496 11608 20502 11620
rect 21085 11611 21143 11617
rect 21085 11608 21097 11611
rect 20496 11580 21097 11608
rect 20496 11568 20502 11580
rect 21085 11577 21097 11580
rect 21131 11577 21143 11611
rect 21085 11571 21143 11577
rect 21284 11552 21312 11648
rect 14182 11540 14188 11552
rect 11256 11512 14188 11540
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14550 11500 14556 11552
rect 14608 11500 14614 11552
rect 14642 11500 14648 11552
rect 14700 11500 14706 11552
rect 15286 11500 15292 11552
rect 15344 11500 15350 11552
rect 15381 11543 15439 11549
rect 15381 11509 15393 11543
rect 15427 11540 15439 11543
rect 15562 11540 15568 11552
rect 15427 11512 15568 11540
rect 15427 11509 15439 11512
rect 15381 11503 15439 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 15654 11500 15660 11552
rect 15712 11500 15718 11552
rect 16022 11500 16028 11552
rect 16080 11500 16086 11552
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 18969 11543 19027 11549
rect 18969 11540 18981 11543
rect 18288 11512 18981 11540
rect 18288 11500 18294 11512
rect 18969 11509 18981 11512
rect 19015 11509 19027 11543
rect 18969 11503 19027 11509
rect 19610 11500 19616 11552
rect 19668 11540 19674 11552
rect 19705 11543 19763 11549
rect 19705 11540 19717 11543
rect 19668 11512 19717 11540
rect 19668 11500 19674 11512
rect 19705 11509 19717 11512
rect 19751 11509 19763 11543
rect 19705 11503 19763 11509
rect 21266 11500 21272 11552
rect 21324 11500 21330 11552
rect 22066 11540 22094 11784
rect 22664 11784 22784 11812
rect 22664 11753 22692 11784
rect 23474 11772 23480 11824
rect 23532 11772 23538 11824
rect 22649 11747 22707 11753
rect 22649 11713 22661 11747
rect 22695 11713 22707 11747
rect 22649 11707 22707 11713
rect 22925 11679 22983 11685
rect 22925 11645 22937 11679
rect 22971 11676 22983 11679
rect 23658 11676 23664 11688
rect 22971 11648 23664 11676
rect 22971 11645 22983 11648
rect 22925 11639 22983 11645
rect 23658 11636 23664 11648
rect 23716 11636 23722 11688
rect 25958 11568 25964 11620
rect 26016 11568 26022 11620
rect 25976 11540 26004 11568
rect 22066 11512 26004 11540
rect 1104 11450 26496 11472
rect 1104 11398 4124 11450
rect 4176 11398 4188 11450
rect 4240 11398 4252 11450
rect 4304 11398 4316 11450
rect 4368 11398 4380 11450
rect 4432 11398 10472 11450
rect 10524 11398 10536 11450
rect 10588 11398 10600 11450
rect 10652 11398 10664 11450
rect 10716 11398 10728 11450
rect 10780 11398 16820 11450
rect 16872 11398 16884 11450
rect 16936 11398 16948 11450
rect 17000 11398 17012 11450
rect 17064 11398 17076 11450
rect 17128 11398 23168 11450
rect 23220 11398 23232 11450
rect 23284 11398 23296 11450
rect 23348 11398 23360 11450
rect 23412 11398 23424 11450
rect 23476 11398 26496 11450
rect 1104 11376 26496 11398
rect 1660 11339 1718 11345
rect 1660 11305 1672 11339
rect 1706 11336 1718 11339
rect 2130 11336 2136 11348
rect 1706 11308 2136 11336
rect 1706 11305 1718 11308
rect 1660 11299 1718 11305
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2866 11296 2872 11348
rect 2924 11296 2930 11348
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3878 11336 3884 11348
rect 3191 11308 3884 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 1394 11160 1400 11212
rect 1452 11160 1458 11212
rect 2884 11132 2912 11296
rect 3252 11209 3280 11308
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 3973 11339 4031 11345
rect 3973 11305 3985 11339
rect 4019 11305 4031 11339
rect 3973 11299 4031 11305
rect 3418 11228 3424 11280
rect 3476 11268 3482 11280
rect 3988 11268 4016 11299
rect 4614 11296 4620 11348
rect 4672 11296 4678 11348
rect 4801 11339 4859 11345
rect 4801 11305 4813 11339
rect 4847 11336 4859 11339
rect 4982 11336 4988 11348
rect 4847 11308 4988 11336
rect 4847 11305 4859 11308
rect 4801 11299 4859 11305
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 5994 11296 6000 11348
rect 6052 11296 6058 11348
rect 8110 11336 8116 11348
rect 7760 11308 8116 11336
rect 4706 11268 4712 11280
rect 3476 11240 4016 11268
rect 4080 11240 4712 11268
rect 3476 11228 3482 11240
rect 3237 11203 3295 11209
rect 3237 11169 3249 11203
rect 3283 11169 3295 11203
rect 3237 11163 3295 11169
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4080 11200 4108 11240
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 4798 11200 4804 11212
rect 3936 11172 4108 11200
rect 4172 11172 4804 11200
rect 3936 11160 3942 11172
rect 3421 11135 3479 11141
rect 3421 11132 3433 11135
rect 2884 11104 3433 11132
rect 3421 11101 3433 11104
rect 3467 11101 3479 11135
rect 3421 11095 3479 11101
rect 3142 11064 3148 11076
rect 2898 11036 3148 11064
rect 3142 11024 3148 11036
rect 3200 11024 3206 11076
rect 3605 11067 3663 11073
rect 3605 11033 3617 11067
rect 3651 11064 3663 11067
rect 3694 11064 3700 11076
rect 3651 11036 3700 11064
rect 3651 11033 3663 11036
rect 3605 11027 3663 11033
rect 3694 11024 3700 11036
rect 3752 11064 3758 11076
rect 4172 11073 4200 11172
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 5000 11141 5028 11296
rect 5534 11228 5540 11280
rect 5592 11228 5598 11280
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 5184 11172 6469 11200
rect 5184 11141 5212 11172
rect 6457 11169 6469 11172
rect 6503 11169 6515 11203
rect 6457 11163 6515 11169
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11132 5411 11135
rect 5442 11132 5448 11144
rect 5399 11104 5448 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5718 11132 5724 11144
rect 5552 11104 5724 11132
rect 3941 11067 3999 11073
rect 3941 11064 3953 11067
rect 3752 11036 3953 11064
rect 3752 11024 3758 11036
rect 3941 11033 3953 11036
rect 3987 11033 3999 11067
rect 3941 11027 3999 11033
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11033 4215 11067
rect 4157 11027 4215 11033
rect 4433 11067 4491 11073
rect 4433 11033 4445 11067
rect 4479 11064 4491 11067
rect 4522 11064 4528 11076
rect 4479 11036 4528 11064
rect 4479 11033 4491 11036
rect 4433 11027 4491 11033
rect 3786 10956 3792 11008
rect 3844 10956 3850 11008
rect 3956 10996 3984 11027
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5552 11064 5580 11104
rect 5718 11092 5724 11104
rect 5776 11132 5782 11144
rect 5776 11104 6316 11132
rect 5776 11092 5782 11104
rect 5307 11036 5580 11064
rect 5629 11067 5687 11073
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5629 11033 5641 11067
rect 5675 11033 5687 11067
rect 5629 11027 5687 11033
rect 5813 11067 5871 11073
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 6178 11064 6184 11076
rect 5859 11036 6184 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 4338 10996 4344 11008
rect 3956 10968 4344 10996
rect 4338 10956 4344 10968
rect 4396 10996 4402 11008
rect 4633 10999 4691 11005
rect 4633 10996 4645 10999
rect 4396 10968 4645 10996
rect 4396 10956 4402 10968
rect 4633 10965 4645 10968
rect 4679 10965 4691 10999
rect 4633 10959 4691 10965
rect 5166 10956 5172 11008
rect 5224 10996 5230 11008
rect 5644 10996 5672 11027
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 6288 11064 6316 11104
rect 6362 11092 6368 11144
rect 6420 11092 6426 11144
rect 6549 11135 6607 11141
rect 6549 11101 6561 11135
rect 6595 11101 6607 11135
rect 7760 11132 7788 11308
rect 8110 11296 8116 11308
rect 8168 11336 8174 11348
rect 9674 11336 9680 11348
rect 8168 11308 9680 11336
rect 8168 11296 8174 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 14553 11339 14611 11345
rect 14553 11336 14565 11339
rect 9824 11308 14565 11336
rect 9824 11296 9830 11308
rect 14553 11305 14565 11308
rect 14599 11336 14611 11339
rect 15194 11336 15200 11348
rect 14599 11308 15200 11336
rect 14599 11305 14611 11308
rect 14553 11299 14611 11305
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 15838 11296 15844 11348
rect 15896 11336 15902 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 15896 11308 15945 11336
rect 15896 11296 15902 11308
rect 15933 11305 15945 11308
rect 15979 11305 15991 11339
rect 15933 11299 15991 11305
rect 16390 11296 16396 11348
rect 16448 11296 16454 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18012 11308 21680 11336
rect 18012 11296 18018 11308
rect 14645 11271 14703 11277
rect 14645 11268 14657 11271
rect 7852 11240 8892 11268
rect 7852 11209 7880 11240
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 8757 11203 8815 11209
rect 8757 11200 8769 11203
rect 8628 11172 8769 11200
rect 8628 11160 8634 11172
rect 8757 11169 8769 11172
rect 8803 11169 8815 11203
rect 8757 11163 8815 11169
rect 8864 11144 8892 11240
rect 9416 11240 14657 11268
rect 9416 11209 9444 11240
rect 14645 11237 14657 11240
rect 14691 11237 14703 11271
rect 16022 11268 16028 11280
rect 14645 11231 14703 11237
rect 15315 11240 16028 11268
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11169 9551 11203
rect 15315 11200 15343 11240
rect 15562 11200 15568 11212
rect 9493 11163 9551 11169
rect 14568 11172 15343 11200
rect 15396 11172 15568 11200
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7760 11104 8033 11132
rect 6549 11095 6607 11101
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 6564 11064 6592 11095
rect 8478 11092 8484 11144
rect 8536 11092 8542 11144
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11101 8723 11135
rect 8665 11095 8723 11101
rect 6288 11036 6592 11064
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 8680 11064 8708 11095
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 8904 11104 9321 11132
rect 8904 11092 8910 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 8251 11036 8708 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 9214 11024 9220 11076
rect 9272 11064 9278 11076
rect 9508 11064 9536 11163
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11132 14427 11135
rect 14458 11132 14464 11144
rect 14415 11104 14464 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 14568 11141 14596 11172
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 14734 11092 14740 11144
rect 14792 11141 14798 11144
rect 14792 11135 14841 11141
rect 14792 11101 14795 11135
rect 14829 11101 14841 11135
rect 14792 11095 14841 11101
rect 15196 11135 15254 11141
rect 15196 11101 15208 11135
rect 15242 11101 15254 11135
rect 15196 11095 15254 11101
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11132 15347 11135
rect 15396 11132 15424 11172
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15335 11104 15424 11132
rect 15488 11104 15761 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 14792 11092 14798 11095
rect 9272 11036 9536 11064
rect 9272 11024 9278 11036
rect 13538 11024 13544 11076
rect 13596 11064 13602 11076
rect 14921 11067 14979 11073
rect 14921 11064 14933 11067
rect 13596 11036 14933 11064
rect 13596 11024 13602 11036
rect 14921 11033 14933 11036
rect 14967 11033 14979 11067
rect 14921 11027 14979 11033
rect 15013 11067 15071 11073
rect 15013 11033 15025 11067
rect 15059 11064 15071 11067
rect 15211 11064 15239 11095
rect 15488 11076 15516 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15948 11132 15976 11240
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 18230 11268 18236 11280
rect 17512 11240 18236 11268
rect 17512 11141 17540 11240
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 18690 11228 18696 11280
rect 18748 11228 18754 11280
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 15948 11104 16221 11132
rect 15749 11095 15807 11101
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11101 17555 11135
rect 17604 11132 17632 11163
rect 17862 11160 17868 11212
rect 17920 11160 17926 11212
rect 18138 11200 18144 11212
rect 17972 11172 18144 11200
rect 17972 11132 18000 11172
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 18708 11200 18736 11228
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 18708 11172 19257 11200
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 19521 11203 19579 11209
rect 19521 11169 19533 11203
rect 19567 11200 19579 11203
rect 19610 11200 19616 11212
rect 19567 11172 19616 11200
rect 19567 11169 19579 11172
rect 19521 11163 19579 11169
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 21266 11160 21272 11212
rect 21324 11160 21330 11212
rect 21652 11144 21680 11308
rect 22738 11296 22744 11348
rect 22796 11296 22802 11348
rect 22465 11203 22523 11209
rect 22465 11169 22477 11203
rect 22511 11200 22523 11203
rect 22756 11200 22784 11296
rect 22511 11172 22784 11200
rect 22511 11169 22523 11172
rect 22465 11163 22523 11169
rect 17604 11104 18000 11132
rect 18233 11135 18291 11141
rect 17497 11095 17555 11101
rect 18233 11101 18245 11135
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 15470 11064 15476 11076
rect 15059 11036 15148 11064
rect 15211 11036 15476 11064
rect 15059 11033 15071 11036
rect 15013 11027 15071 11033
rect 5224 10968 5672 10996
rect 5224 10956 5230 10968
rect 8294 10956 8300 11008
rect 8352 10956 8358 11008
rect 8938 10956 8944 11008
rect 8996 10956 9002 11008
rect 15120 10996 15148 11036
rect 15470 11024 15476 11036
rect 15528 11024 15534 11076
rect 15565 11067 15623 11073
rect 15565 11033 15577 11067
rect 15611 11064 15623 11067
rect 16025 11067 16083 11073
rect 15611 11036 15982 11064
rect 15611 11033 15623 11036
rect 15565 11027 15623 11033
rect 15194 10996 15200 11008
rect 15120 10968 15200 10996
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 15381 10999 15439 11005
rect 15381 10996 15393 10999
rect 15344 10968 15393 10996
rect 15344 10956 15350 10968
rect 15381 10965 15393 10968
rect 15427 10965 15439 10999
rect 15954 10996 15982 11036
rect 16025 11033 16037 11067
rect 16071 11064 16083 11067
rect 16298 11064 16304 11076
rect 16071 11036 16304 11064
rect 16071 11033 16083 11036
rect 16025 11027 16083 11033
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 16482 11024 16488 11076
rect 16540 11024 16546 11076
rect 16666 11024 16672 11076
rect 16724 11024 16730 11076
rect 17218 11024 17224 11076
rect 17276 11024 17282 11076
rect 17236 10996 17264 11024
rect 15954 10968 17264 10996
rect 18248 10996 18276 11095
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11132 18751 11135
rect 19150 11132 19156 11144
rect 18739 11104 19156 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 21634 11092 21640 11144
rect 21692 11092 21698 11144
rect 18601 11067 18659 11073
rect 18601 11033 18613 11067
rect 18647 11064 18659 11067
rect 19794 11064 19800 11076
rect 18647 11036 19800 11064
rect 18647 11033 18659 11036
rect 18601 11027 18659 11033
rect 19794 11024 19800 11036
rect 19852 11024 19858 11076
rect 22094 11064 22100 11076
rect 19904 11036 20010 11064
rect 20824 11036 22100 11064
rect 18690 10996 18696 11008
rect 18248 10968 18696 10996
rect 15381 10959 15439 10965
rect 18690 10956 18696 10968
rect 18748 10996 18754 11008
rect 19518 10996 19524 11008
rect 18748 10968 19524 10996
rect 18748 10956 18754 10968
rect 19518 10956 19524 10968
rect 19576 10956 19582 11008
rect 19610 10956 19616 11008
rect 19668 10996 19674 11008
rect 19904 10996 19932 11036
rect 20824 10996 20852 11036
rect 22094 11024 22100 11036
rect 22152 11024 22158 11076
rect 19668 10968 20852 10996
rect 19668 10956 19674 10968
rect 1104 10906 26656 10928
rect 1104 10854 7298 10906
rect 7350 10854 7362 10906
rect 7414 10854 7426 10906
rect 7478 10854 7490 10906
rect 7542 10854 7554 10906
rect 7606 10854 13646 10906
rect 13698 10854 13710 10906
rect 13762 10854 13774 10906
rect 13826 10854 13838 10906
rect 13890 10854 13902 10906
rect 13954 10854 19994 10906
rect 20046 10854 20058 10906
rect 20110 10854 20122 10906
rect 20174 10854 20186 10906
rect 20238 10854 20250 10906
rect 20302 10854 26342 10906
rect 26394 10854 26406 10906
rect 26458 10854 26470 10906
rect 26522 10854 26534 10906
rect 26586 10854 26598 10906
rect 26650 10854 26656 10906
rect 1104 10832 26656 10854
rect 2593 10795 2651 10801
rect 2593 10761 2605 10795
rect 2639 10761 2651 10795
rect 2593 10755 2651 10761
rect 2961 10795 3019 10801
rect 2961 10761 2973 10795
rect 3007 10792 3019 10795
rect 3786 10792 3792 10804
rect 3007 10764 3792 10792
rect 3007 10761 3019 10764
rect 2961 10755 3019 10761
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2608 10656 2636 10755
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 4706 10752 4712 10804
rect 4764 10752 4770 10804
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5537 10795 5595 10801
rect 5316 10764 5488 10792
rect 5316 10752 5322 10764
rect 3050 10684 3056 10736
rect 3108 10684 3114 10736
rect 3510 10684 3516 10736
rect 3568 10724 3574 10736
rect 3568 10696 3832 10724
rect 3568 10684 3574 10696
rect 2363 10628 2636 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 3694 10616 3700 10668
rect 3752 10616 3758 10668
rect 3804 10665 3832 10696
rect 4250 10681 4308 10687
rect 4338 10684 4344 10736
rect 4396 10684 4402 10736
rect 4614 10733 4620 10736
rect 4571 10727 4620 10733
rect 4571 10693 4583 10727
rect 4617 10693 4620 10727
rect 4250 10678 4262 10681
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3878 10616 3884 10668
rect 3936 10616 3942 10668
rect 4080 10650 4262 10678
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10588 3295 10591
rect 4080 10588 4108 10650
rect 4250 10647 4262 10650
rect 4296 10647 4308 10681
rect 4250 10641 4308 10647
rect 4430 10640 4436 10692
rect 4488 10640 4494 10692
rect 4571 10687 4620 10693
rect 4614 10684 4620 10687
rect 4672 10684 4678 10736
rect 4724 10724 4752 10752
rect 5166 10724 5172 10736
rect 4724 10696 5172 10724
rect 5166 10684 5172 10696
rect 5224 10724 5230 10736
rect 5460 10724 5488 10764
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5718 10792 5724 10804
rect 5583 10764 5724 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 6914 10752 6920 10804
rect 6972 10752 6978 10804
rect 7377 10795 7435 10801
rect 7377 10761 7389 10795
rect 7423 10792 7435 10795
rect 8938 10792 8944 10804
rect 7423 10764 8944 10792
rect 7423 10761 7435 10764
rect 7377 10755 7435 10761
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 9732 10764 9781 10792
rect 9732 10752 9738 10764
rect 9769 10761 9781 10764
rect 9815 10792 9827 10795
rect 14645 10795 14703 10801
rect 14645 10792 14657 10795
rect 9815 10764 14657 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 14645 10761 14657 10764
rect 14691 10761 14703 10795
rect 14645 10755 14703 10761
rect 14737 10795 14795 10801
rect 14737 10761 14749 10795
rect 14783 10792 14795 10795
rect 15105 10795 15163 10801
rect 15105 10792 15117 10795
rect 14783 10764 15117 10792
rect 14783 10761 14795 10764
rect 14737 10755 14795 10761
rect 15105 10761 15117 10764
rect 15151 10761 15163 10795
rect 15105 10755 15163 10761
rect 15654 10752 15660 10804
rect 15712 10752 15718 10804
rect 16482 10752 16488 10804
rect 16540 10792 16546 10804
rect 18506 10792 18512 10804
rect 16540 10764 18512 10792
rect 16540 10752 16546 10764
rect 6549 10727 6607 10733
rect 6549 10724 6561 10727
rect 5224 10696 5396 10724
rect 5460 10696 6561 10724
rect 5224 10684 5230 10696
rect 5368 10665 5396 10696
rect 6549 10693 6561 10696
rect 6595 10693 6607 10727
rect 6549 10687 6607 10693
rect 6822 10684 6828 10736
rect 6880 10724 6886 10736
rect 6880 10696 8064 10724
rect 6880 10684 6886 10696
rect 5353 10659 5411 10665
rect 4433 10625 4445 10640
rect 4479 10625 4491 10640
rect 4433 10619 4491 10625
rect 4566 10628 5120 10656
rect 4566 10588 4594 10628
rect 5092 10600 5120 10628
rect 5353 10625 5365 10659
rect 5399 10625 5411 10659
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5353 10619 5411 10625
rect 5460 10628 6377 10656
rect 3283 10560 3372 10588
rect 4080 10560 4594 10588
rect 4709 10591 4767 10597
rect 3283 10557 3295 10560
rect 3237 10551 3295 10557
rect 3344 10520 3372 10560
rect 4709 10557 4721 10591
rect 4755 10588 4767 10591
rect 4801 10591 4859 10597
rect 4801 10588 4813 10591
rect 4755 10560 4813 10588
rect 4755 10557 4767 10560
rect 4709 10551 4767 10557
rect 4801 10557 4813 10560
rect 4847 10557 4859 10591
rect 4801 10551 4859 10557
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5460 10588 5488 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 7190 10616 7196 10668
rect 7248 10656 7254 10668
rect 8036 10665 8064 10696
rect 8294 10684 8300 10736
rect 8352 10684 8358 10736
rect 12345 10727 12403 10733
rect 12345 10693 12357 10727
rect 12391 10724 12403 10727
rect 12802 10724 12808 10736
rect 12391 10696 12808 10724
rect 12391 10693 12403 10696
rect 12345 10687 12403 10693
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 15378 10684 15384 10736
rect 15436 10684 15442 10736
rect 15672 10724 15700 10752
rect 16761 10727 16819 10733
rect 16761 10724 16773 10727
rect 15672 10696 15792 10724
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 7248 10628 7297 10656
rect 7248 10616 7254 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 9364 10628 9430 10656
rect 9364 10616 9370 10628
rect 10870 10616 10876 10668
rect 10928 10656 10934 10668
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 10928 10628 11161 10656
rect 10928 10616 10934 10628
rect 11149 10625 11161 10628
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12526 10656 12532 10668
rect 12483 10628 12532 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 5132 10560 5488 10588
rect 5132 10548 5138 10560
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6638 10588 6644 10600
rect 6236 10560 6644 10588
rect 6236 10548 6242 10560
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 12176 10588 12204 10619
rect 12526 10616 12532 10628
rect 12584 10656 12590 10668
rect 13170 10656 13176 10668
rect 12584 10628 13176 10656
rect 12584 10616 12590 10628
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 14734 10616 14740 10668
rect 14792 10656 14798 10668
rect 15284 10659 15342 10665
rect 15284 10656 15296 10659
rect 14792 10628 15296 10656
rect 14792 10616 14798 10628
rect 15284 10625 15296 10628
rect 15330 10625 15342 10659
rect 15284 10619 15342 10625
rect 12710 10588 12716 10600
rect 7607 10560 8156 10588
rect 12176 10560 12716 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 3602 10520 3608 10532
rect 3344 10492 3608 10520
rect 3602 10480 3608 10492
rect 3660 10520 3666 10532
rect 4430 10520 4436 10532
rect 3660 10492 4436 10520
rect 3660 10480 3666 10492
rect 4430 10480 4436 10492
rect 4488 10480 4494 10532
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 5442 10520 5448 10532
rect 4672 10492 5448 10520
rect 4672 10480 4678 10492
rect 5442 10480 5448 10492
rect 5500 10520 5506 10532
rect 6733 10523 6791 10529
rect 6733 10520 6745 10523
rect 5500 10492 6745 10520
rect 5500 10480 5506 10492
rect 6733 10489 6745 10492
rect 6779 10489 6791 10523
rect 6733 10483 6791 10489
rect 8128 10464 8156 10560
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 14829 10591 14887 10597
rect 14829 10588 14841 10591
rect 14240 10560 14841 10588
rect 14240 10548 14246 10560
rect 14829 10557 14841 10560
rect 14875 10557 14887 10591
rect 15304 10588 15332 10619
rect 15470 10616 15476 10668
rect 15528 10616 15534 10668
rect 15562 10616 15568 10668
rect 15620 10665 15626 10668
rect 15764 10665 15792 10696
rect 15856 10696 16773 10724
rect 15620 10659 15659 10665
rect 15647 10625 15659 10659
rect 15620 10619 15659 10625
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 15620 10616 15626 10619
rect 15856 10588 15884 10696
rect 16761 10693 16773 10696
rect 16807 10693 16819 10727
rect 16761 10687 16819 10693
rect 16390 10616 16396 10668
rect 16448 10616 16454 10668
rect 16666 10616 16672 10668
rect 16724 10616 16730 10668
rect 16960 10665 16988 10764
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 17862 10684 17868 10736
rect 17920 10684 17926 10736
rect 18322 10684 18328 10736
rect 18380 10684 18386 10736
rect 19518 10684 19524 10736
rect 19576 10724 19582 10736
rect 19613 10727 19671 10733
rect 19613 10724 19625 10727
rect 19576 10696 19625 10724
rect 19576 10684 19582 10696
rect 19613 10693 19625 10696
rect 19659 10693 19671 10727
rect 19613 10687 19671 10693
rect 19794 10684 19800 10736
rect 19852 10724 19858 10736
rect 20533 10727 20591 10733
rect 20533 10724 20545 10727
rect 19852 10696 20545 10724
rect 19852 10684 19858 10696
rect 20533 10693 20545 10696
rect 20579 10693 20591 10727
rect 20533 10687 20591 10693
rect 21634 10684 21640 10736
rect 21692 10724 21698 10736
rect 21821 10727 21879 10733
rect 21821 10724 21833 10727
rect 21692 10696 21833 10724
rect 21692 10684 21698 10696
rect 21821 10693 21833 10696
rect 21867 10693 21879 10727
rect 21821 10687 21879 10693
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 15304 10560 15884 10588
rect 16117 10591 16175 10597
rect 14829 10551 14887 10557
rect 15396 10532 15424 10560
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16298 10588 16304 10600
rect 16163 10560 16304 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 14642 10520 14648 10532
rect 9456 10492 14648 10520
rect 9456 10480 9462 10492
rect 14642 10480 14648 10492
rect 14700 10480 14706 10532
rect 15378 10480 15384 10532
rect 15436 10480 15442 10532
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 16684 10520 16712 10616
rect 16868 10588 16896 10619
rect 17402 10616 17408 10668
rect 17460 10656 17466 10668
rect 17589 10659 17647 10665
rect 17589 10656 17601 10659
rect 17460 10628 17601 10656
rect 17460 10616 17466 10628
rect 17589 10625 17601 10628
rect 17635 10625 17647 10659
rect 17589 10619 17647 10625
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19392 10628 19717 10656
rect 19392 10616 19398 10628
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 19886 10616 19892 10668
rect 19944 10616 19950 10668
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10656 20315 10659
rect 20346 10656 20352 10668
rect 20303 10628 20352 10656
rect 20303 10625 20315 10628
rect 20257 10619 20315 10625
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 16868 10560 17080 10588
rect 15620 10492 16712 10520
rect 15620 10480 15626 10492
rect 2130 10412 2136 10464
rect 2188 10412 2194 10464
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10452 4123 10455
rect 4522 10452 4528 10464
rect 4111 10424 4528 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 8110 10412 8116 10464
rect 8168 10412 8174 10464
rect 10962 10412 10968 10464
rect 11020 10412 11026 10464
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 12124 10424 12173 10452
rect 12124 10412 12130 10424
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 14274 10412 14280 10464
rect 14332 10412 14338 10464
rect 15838 10412 15844 10464
rect 15896 10412 15902 10464
rect 16301 10455 16359 10461
rect 16301 10421 16313 10455
rect 16347 10452 16359 10455
rect 16482 10452 16488 10464
rect 16347 10424 16488 10452
rect 16347 10421 16359 10424
rect 16301 10415 16359 10421
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 17052 10461 17080 10560
rect 18322 10548 18328 10600
rect 18380 10588 18386 10600
rect 19610 10588 19616 10600
rect 18380 10560 19616 10588
rect 18380 10548 18386 10560
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 22554 10548 22560 10600
rect 22612 10548 22618 10600
rect 17037 10455 17095 10461
rect 17037 10421 17049 10455
rect 17083 10452 17095 10455
rect 17218 10452 17224 10464
rect 17083 10424 17224 10452
rect 17083 10421 17095 10424
rect 17037 10415 17095 10421
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 19242 10452 19248 10464
rect 18104 10424 19248 10452
rect 18104 10412 18110 10424
rect 19242 10412 19248 10424
rect 19300 10452 19306 10464
rect 19797 10455 19855 10461
rect 19797 10452 19809 10455
rect 19300 10424 19809 10452
rect 19300 10412 19306 10424
rect 19797 10421 19809 10424
rect 19843 10421 19855 10455
rect 19797 10415 19855 10421
rect 1104 10362 26496 10384
rect 1104 10310 4124 10362
rect 4176 10310 4188 10362
rect 4240 10310 4252 10362
rect 4304 10310 4316 10362
rect 4368 10310 4380 10362
rect 4432 10310 10472 10362
rect 10524 10310 10536 10362
rect 10588 10310 10600 10362
rect 10652 10310 10664 10362
rect 10716 10310 10728 10362
rect 10780 10310 16820 10362
rect 16872 10310 16884 10362
rect 16936 10310 16948 10362
rect 17000 10310 17012 10362
rect 17064 10310 17076 10362
rect 17128 10310 23168 10362
rect 23220 10310 23232 10362
rect 23284 10310 23296 10362
rect 23348 10310 23360 10362
rect 23412 10310 23424 10362
rect 23476 10310 26496 10362
rect 1104 10288 26496 10310
rect 1752 10251 1810 10257
rect 1752 10217 1764 10251
rect 1798 10248 1810 10251
rect 2130 10248 2136 10260
rect 1798 10220 2136 10248
rect 1798 10217 1810 10220
rect 1752 10211 1810 10217
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3602 10248 3608 10260
rect 3283 10220 3608 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4522 10208 4528 10260
rect 4580 10208 4586 10260
rect 5156 10251 5214 10257
rect 5156 10217 5168 10251
rect 5202 10248 5214 10251
rect 5534 10248 5540 10260
rect 5202 10220 5540 10248
rect 5202 10217 5214 10220
rect 5156 10211 5214 10217
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 6638 10208 6644 10260
rect 6696 10208 6702 10260
rect 9398 10208 9404 10260
rect 9456 10208 9462 10260
rect 9490 10208 9496 10260
rect 9548 10208 9554 10260
rect 10962 10208 10968 10260
rect 11020 10208 11026 10260
rect 15562 10208 15568 10260
rect 15620 10208 15626 10260
rect 15838 10208 15844 10260
rect 15896 10208 15902 10260
rect 15930 10208 15936 10260
rect 15988 10248 15994 10260
rect 16390 10248 16396 10260
rect 15988 10220 16396 10248
rect 15988 10208 15994 10220
rect 16390 10208 16396 10220
rect 16448 10248 16454 10260
rect 16485 10251 16543 10257
rect 16485 10248 16497 10251
rect 16448 10220 16497 10248
rect 16448 10208 16454 10220
rect 16485 10217 16497 10220
rect 16531 10217 16543 10251
rect 16485 10211 16543 10217
rect 18509 10251 18567 10257
rect 18509 10217 18521 10251
rect 18555 10248 18567 10251
rect 19702 10248 19708 10260
rect 18555 10220 19708 10248
rect 18555 10217 18567 10220
rect 18509 10211 18567 10217
rect 1394 10072 1400 10124
rect 1452 10112 1458 10124
rect 1489 10115 1547 10121
rect 1489 10112 1501 10115
rect 1452 10084 1501 10112
rect 1452 10072 1458 10084
rect 1489 10081 1501 10084
rect 1535 10112 1547 10115
rect 1854 10112 1860 10124
rect 1535 10084 1860 10112
rect 1535 10081 1547 10084
rect 1489 10075 1547 10081
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 4540 10121 4568 10208
rect 9416 10180 9444 10208
rect 9324 10152 9444 10180
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4893 10115 4951 10121
rect 4893 10081 4905 10115
rect 4939 10112 4951 10115
rect 5534 10112 5540 10124
rect 4939 10084 5540 10112
rect 4939 10081 4951 10084
rect 4893 10075 4951 10081
rect 5534 10072 5540 10084
rect 5592 10112 5598 10124
rect 6822 10112 6828 10124
rect 5592 10084 6828 10112
rect 5592 10072 5598 10084
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7208 10084 7880 10112
rect 7208 10056 7236 10084
rect 7190 10004 7196 10056
rect 7248 10004 7254 10056
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7650 10044 7656 10056
rect 7515 10016 7656 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 7852 10053 7880 10084
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8110 10044 8116 10056
rect 8067 10016 8116 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 3142 9976 3148 9988
rect 2990 9948 3148 9976
rect 3142 9936 3148 9948
rect 3200 9976 3206 9988
rect 3786 9976 3792 9988
rect 3200 9948 3792 9976
rect 3200 9936 3206 9948
rect 3786 9936 3792 9948
rect 3844 9936 3850 9988
rect 7006 9976 7012 9988
rect 6394 9948 7012 9976
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 9324 9976 9352 10152
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 9508 10112 9536 10208
rect 9447 10084 9536 10112
rect 9677 10115 9735 10121
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10980 10112 11008 10208
rect 9723 10084 11008 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 11112 10084 11253 10112
rect 11112 10072 11118 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 12860 10084 13124 10112
rect 12860 10072 12866 10084
rect 13096 10056 13124 10084
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 13228 10084 13308 10112
rect 13228 10072 13234 10084
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 13280 10053 13308 10084
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10044 15439 10047
rect 15856 10044 15884 10208
rect 16500 10180 16528 10211
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 22738 10208 22744 10260
rect 22796 10248 22802 10260
rect 23477 10251 23535 10257
rect 23477 10248 23489 10251
rect 22796 10220 23489 10248
rect 22796 10208 22802 10220
rect 23477 10217 23489 10220
rect 23523 10217 23535 10251
rect 23477 10211 23535 10217
rect 16500 10152 18736 10180
rect 16482 10072 16488 10124
rect 16540 10112 16546 10124
rect 16540 10084 16896 10112
rect 16540 10072 16546 10084
rect 15427 10016 15884 10044
rect 16025 10047 16083 10053
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 16025 10013 16037 10047
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 7668 9948 9352 9976
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 3973 9911 4031 9917
rect 3973 9908 3985 9911
rect 3936 9880 3985 9908
rect 3936 9868 3942 9880
rect 3973 9877 3985 9880
rect 4019 9877 4031 9911
rect 3973 9871 4031 9877
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7668 9917 7696 9948
rect 10134 9936 10140 9988
rect 10192 9936 10198 9988
rect 11514 9936 11520 9988
rect 11572 9936 11578 9988
rect 12894 9976 12900 9988
rect 12742 9948 12900 9976
rect 12894 9936 12900 9948
rect 12952 9936 12958 9988
rect 14458 9936 14464 9988
rect 14516 9976 14522 9988
rect 16040 9976 16068 10007
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 16868 10053 16896 10084
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 18141 10115 18199 10121
rect 18141 10112 18153 10115
rect 17276 10084 18153 10112
rect 17276 10072 17282 10084
rect 18141 10081 18153 10084
rect 18187 10081 18199 10115
rect 18141 10075 18199 10081
rect 18708 10056 18736 10152
rect 18874 10140 18880 10192
rect 18932 10140 18938 10192
rect 19242 10140 19248 10192
rect 19300 10140 19306 10192
rect 19794 10140 19800 10192
rect 19852 10180 19858 10192
rect 19852 10152 20208 10180
rect 19852 10140 19858 10152
rect 19260 10112 19288 10140
rect 19260 10084 20024 10112
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 16172 10016 16221 10044
rect 16172 10004 16178 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 18046 10004 18052 10056
rect 18104 10044 18110 10056
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 18104 10016 18337 10044
rect 18104 10004 18110 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18601 10047 18659 10053
rect 18601 10013 18613 10047
rect 18647 10013 18659 10047
rect 18601 10007 18659 10013
rect 16298 9976 16304 9988
rect 14516 9948 16304 9976
rect 14516 9936 14522 9948
rect 16298 9936 16304 9948
rect 16356 9976 16362 9988
rect 16439 9979 16497 9985
rect 16439 9976 16451 9979
rect 16356 9948 16451 9976
rect 16356 9936 16362 9948
rect 16439 9945 16451 9948
rect 16485 9945 16497 9979
rect 18616 9976 18644 10007
rect 18690 10004 18696 10056
rect 18748 10004 18754 10056
rect 19610 10004 19616 10056
rect 19668 10044 19674 10056
rect 19996 10053 20024 10084
rect 20180 10053 20208 10152
rect 20898 10072 20904 10124
rect 20956 10072 20962 10124
rect 23750 10112 23756 10124
rect 22204 10084 23756 10112
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19668 10016 19809 10044
rect 19668 10004 19674 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 20165 10047 20223 10053
rect 20165 10013 20177 10047
rect 20211 10013 20223 10047
rect 20165 10007 20223 10013
rect 22204 9988 22232 10084
rect 23750 10072 23756 10084
rect 23808 10072 23814 10124
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 23164 10016 23213 10044
rect 23164 10004 23170 10016
rect 23201 10013 23213 10016
rect 23247 10013 23259 10047
rect 23201 10007 23259 10013
rect 24578 10004 24584 10056
rect 24636 10004 24642 10056
rect 24854 10025 24912 10031
rect 24854 9991 24866 10025
rect 24900 9991 24912 10025
rect 25498 10004 25504 10056
rect 25556 10004 25562 10056
rect 24854 9988 24912 9991
rect 16439 9939 16497 9945
rect 18156 9948 18644 9976
rect 18877 9979 18935 9985
rect 18156 9920 18184 9948
rect 18877 9945 18889 9979
rect 18923 9976 18935 9979
rect 19245 9979 19303 9985
rect 19245 9976 19257 9979
rect 18923 9948 19257 9976
rect 18923 9945 18935 9948
rect 18877 9939 18935 9945
rect 19245 9945 19257 9948
rect 19291 9945 19303 9979
rect 19245 9939 19303 9945
rect 21174 9936 21180 9988
rect 21232 9936 21238 9988
rect 22186 9936 22192 9988
rect 22244 9936 22250 9988
rect 22830 9936 22836 9988
rect 22888 9976 22894 9988
rect 22925 9979 22983 9985
rect 22925 9976 22937 9979
rect 22888 9948 22937 9976
rect 22888 9936 22894 9948
rect 22925 9945 22937 9948
rect 22971 9976 22983 9979
rect 23293 9979 23351 9985
rect 23293 9976 23305 9979
rect 22971 9948 23305 9976
rect 22971 9945 22983 9948
rect 22925 9939 22983 9945
rect 23293 9945 23305 9948
rect 23339 9945 23351 9979
rect 23293 9939 23351 9945
rect 24854 9936 24860 9988
rect 24912 9936 24918 9988
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 6972 9880 7297 9908
rect 6972 9868 6978 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 7653 9911 7711 9917
rect 7653 9877 7665 9911
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 7926 9868 7932 9920
rect 7984 9868 7990 9920
rect 11149 9911 11207 9917
rect 11149 9877 11161 9911
rect 11195 9908 11207 9911
rect 11698 9908 11704 9920
rect 11195 9880 11704 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 11698 9868 11704 9880
rect 11756 9908 11762 9920
rect 12342 9908 12348 9920
rect 11756 9880 12348 9908
rect 11756 9868 11762 9880
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12860 9880 13001 9908
rect 12860 9868 12866 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 13173 9911 13231 9917
rect 13173 9877 13185 9911
rect 13219 9908 13231 9911
rect 13354 9908 13360 9920
rect 13219 9880 13360 9908
rect 13219 9877 13231 9880
rect 13173 9871 13231 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 15197 9911 15255 9917
rect 15197 9877 15209 9911
rect 15243 9908 15255 9911
rect 15286 9908 15292 9920
rect 15243 9880 15292 9908
rect 15243 9877 15255 9880
rect 15197 9871 15255 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 18138 9868 18144 9920
rect 18196 9868 18202 9920
rect 20073 9911 20131 9917
rect 20073 9877 20085 9911
rect 20119 9908 20131 9911
rect 20438 9908 20444 9920
rect 20119 9880 20444 9908
rect 20119 9877 20131 9880
rect 20073 9871 20131 9877
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 23014 9868 23020 9920
rect 23072 9868 23078 9920
rect 23474 9868 23480 9920
rect 23532 9917 23538 9920
rect 23532 9911 23551 9917
rect 23539 9877 23551 9911
rect 23532 9871 23551 9877
rect 23532 9868 23538 9871
rect 23658 9868 23664 9920
rect 23716 9868 23722 9920
rect 24394 9868 24400 9920
rect 24452 9868 24458 9920
rect 24765 9911 24823 9917
rect 24765 9877 24777 9911
rect 24811 9908 24823 9911
rect 25038 9908 25044 9920
rect 24811 9880 25044 9908
rect 24811 9877 24823 9880
rect 24765 9871 24823 9877
rect 25038 9868 25044 9880
rect 25096 9868 25102 9920
rect 25314 9868 25320 9920
rect 25372 9868 25378 9920
rect 1104 9818 26656 9840
rect 1104 9766 7298 9818
rect 7350 9766 7362 9818
rect 7414 9766 7426 9818
rect 7478 9766 7490 9818
rect 7542 9766 7554 9818
rect 7606 9766 13646 9818
rect 13698 9766 13710 9818
rect 13762 9766 13774 9818
rect 13826 9766 13838 9818
rect 13890 9766 13902 9818
rect 13954 9766 19994 9818
rect 20046 9766 20058 9818
rect 20110 9766 20122 9818
rect 20174 9766 20186 9818
rect 20238 9766 20250 9818
rect 20302 9766 26342 9818
rect 26394 9766 26406 9818
rect 26458 9766 26470 9818
rect 26522 9766 26534 9818
rect 26586 9766 26598 9818
rect 26650 9766 26656 9818
rect 1104 9744 26656 9766
rect 5534 9704 5540 9716
rect 4172 9676 5540 9704
rect 4172 9636 4200 9676
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 7006 9704 7012 9716
rect 5644 9676 7012 9704
rect 5644 9636 5672 9676
rect 7006 9664 7012 9676
rect 7064 9704 7070 9716
rect 7558 9704 7564 9716
rect 7064 9676 7564 9704
rect 7064 9664 7070 9676
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 7650 9664 7656 9716
rect 7708 9704 7714 9716
rect 7834 9704 7840 9716
rect 7708 9676 7840 9704
rect 7708 9664 7714 9676
rect 7834 9664 7840 9676
rect 7892 9704 7898 9716
rect 8021 9707 8079 9713
rect 8021 9704 8033 9707
rect 7892 9676 8033 9704
rect 7892 9664 7898 9676
rect 8021 9673 8033 9676
rect 8067 9673 8079 9707
rect 8021 9667 8079 9673
rect 8110 9664 8116 9716
rect 8168 9664 8174 9716
rect 9398 9664 9404 9716
rect 9456 9664 9462 9716
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 13817 9707 13875 9713
rect 13817 9704 13829 9707
rect 13320 9676 13829 9704
rect 13320 9664 13326 9676
rect 13817 9673 13829 9676
rect 13863 9673 13875 9707
rect 21085 9707 21143 9713
rect 13817 9667 13875 9673
rect 18248 9676 19196 9704
rect 8128 9636 8156 9664
rect 9416 9636 9444 9664
rect 11054 9636 11060 9648
rect 3528 9608 4200 9636
rect 5014 9622 5672 9636
rect 5000 9608 5672 9622
rect 7576 9608 8248 9636
rect 9338 9608 9444 9636
rect 10060 9608 11060 9636
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 3528 9577 3556 9608
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 1912 9540 3525 9568
rect 1912 9528 1918 9540
rect 3513 9537 3525 9540
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 3878 9500 3884 9512
rect 3835 9472 3884 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 3878 9324 3884 9376
rect 3936 9364 3942 9376
rect 5000 9364 5028 9608
rect 5166 9528 5172 9580
rect 5224 9528 5230 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7576 9577 7604 9608
rect 7561 9571 7619 9577
rect 7561 9568 7573 9571
rect 7064 9540 7573 9568
rect 7064 9528 7070 9540
rect 7561 9537 7573 9540
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9537 8171 9571
rect 8220 9568 8248 9608
rect 10060 9577 10088 9608
rect 11054 9596 11060 9608
rect 11112 9636 11118 9648
rect 11149 9639 11207 9645
rect 11149 9636 11161 9639
rect 11112 9608 11161 9636
rect 11112 9596 11118 9608
rect 11149 9605 11161 9608
rect 11195 9636 11207 9639
rect 15749 9639 15807 9645
rect 11195 9608 11560 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 11532 9577 11560 9608
rect 15749 9605 15761 9639
rect 15795 9636 15807 9639
rect 18248 9636 18276 9676
rect 15795 9608 18276 9636
rect 15795 9605 15807 9608
rect 15749 9599 15807 9605
rect 18322 9596 18328 9648
rect 18380 9596 18386 9648
rect 19168 9636 19196 9676
rect 21085 9673 21097 9707
rect 21131 9704 21143 9707
rect 21174 9704 21180 9716
rect 21131 9676 21180 9704
rect 21131 9673 21143 9676
rect 21085 9667 21143 9673
rect 21174 9664 21180 9676
rect 21232 9664 21238 9716
rect 22738 9704 22744 9716
rect 22112 9676 22744 9704
rect 19168 9608 22048 9636
rect 10045 9571 10103 9577
rect 8220 9540 8800 9568
rect 8113 9531 8171 9537
rect 5184 9432 5212 9528
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 7248 9472 7389 9500
rect 7248 9460 7254 9472
rect 7377 9469 7389 9472
rect 7423 9469 7435 9503
rect 8128 9500 8156 9531
rect 8772 9512 8800 9540
rect 10045 9537 10057 9571
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 8202 9500 8208 9512
rect 8128 9472 8208 9500
rect 7377 9463 7435 9469
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 8754 9460 8760 9512
rect 8812 9460 8818 9512
rect 9674 9460 9680 9512
rect 9732 9460 9738 9512
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 5184 9404 5273 9432
rect 5261 9401 5273 9404
rect 5307 9401 5319 9435
rect 5261 9395 5319 9401
rect 8128 9404 8984 9432
rect 8128 9376 8156 9404
rect 3936 9336 5028 9364
rect 3936 9324 3942 9336
rect 7742 9324 7748 9376
rect 7800 9324 7806 9376
rect 8110 9324 8116 9376
rect 8168 9324 8174 9376
rect 8294 9373 8300 9376
rect 8251 9367 8300 9373
rect 8251 9333 8263 9367
rect 8297 9333 8300 9367
rect 8251 9327 8300 9333
rect 8294 9324 8300 9327
rect 8352 9324 8358 9376
rect 8956 9364 8984 9404
rect 10428 9364 10456 9531
rect 12894 9528 12900 9580
rect 12952 9528 12958 9580
rect 13876 9571 13934 9577
rect 13876 9568 13888 9571
rect 13280 9540 13888 9568
rect 11790 9460 11796 9512
rect 11848 9460 11854 9512
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 13280 9500 13308 9540
rect 13876 9537 13888 9540
rect 13922 9568 13934 9571
rect 15841 9571 15899 9577
rect 13922 9540 15332 9568
rect 13922 9537 13934 9540
rect 13876 9531 13934 9537
rect 12308 9472 13308 9500
rect 13357 9503 13415 9509
rect 12308 9460 12314 9472
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 13446 9500 13452 9512
rect 13403 9472 13452 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 15194 9460 15200 9512
rect 15252 9460 15258 9512
rect 15304 9500 15332 9540
rect 15841 9537 15853 9571
rect 15887 9568 15899 9571
rect 16022 9568 16028 9580
rect 15887 9540 16028 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 21008 9577 21036 9608
rect 22020 9580 22048 9608
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9537 21051 9571
rect 20993 9531 21051 9537
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 15304 9472 15945 9500
rect 15933 9469 15945 9472
rect 15979 9500 15991 9503
rect 16114 9500 16120 9512
rect 15979 9472 16120 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9469 17647 9503
rect 17589 9463 17647 9469
rect 17865 9503 17923 9509
rect 17865 9469 17877 9503
rect 17911 9500 17923 9503
rect 18414 9500 18420 9512
rect 17911 9472 18420 9500
rect 17911 9469 17923 9472
rect 17865 9463 17923 9469
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 11020 9404 11652 9432
rect 11020 9392 11026 9404
rect 11330 9364 11336 9376
rect 8956 9336 11336 9364
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 11624 9364 11652 9404
rect 13078 9392 13084 9444
rect 13136 9432 13142 9444
rect 13265 9435 13323 9441
rect 13265 9432 13277 9435
rect 13136 9404 13277 9432
rect 13136 9392 13142 9404
rect 13265 9401 13277 9404
rect 13311 9401 13323 9435
rect 13265 9395 13323 9401
rect 14001 9435 14059 9441
rect 14001 9401 14013 9435
rect 14047 9432 14059 9435
rect 14090 9432 14096 9444
rect 14047 9404 14096 9432
rect 14047 9401 14059 9404
rect 14001 9395 14059 9401
rect 14090 9392 14096 9404
rect 14148 9392 14154 9444
rect 15212 9432 15240 9460
rect 15381 9435 15439 9441
rect 15381 9432 15393 9435
rect 15212 9404 15393 9432
rect 15381 9401 15393 9404
rect 15427 9401 15439 9435
rect 15381 9395 15439 9401
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 11624 9336 13461 9364
rect 13449 9333 13461 9336
rect 13495 9364 13507 9367
rect 14182 9364 14188 9376
rect 13495 9336 14188 9364
rect 13495 9333 13507 9336
rect 13449 9327 13507 9333
rect 14182 9324 14188 9336
rect 14240 9364 14246 9376
rect 15286 9364 15292 9376
rect 14240 9336 15292 9364
rect 14240 9324 14246 9336
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 17604 9364 17632 9463
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 19610 9460 19616 9512
rect 19668 9460 19674 9512
rect 20530 9392 20536 9444
rect 20588 9432 20594 9444
rect 20824 9432 20852 9531
rect 21266 9528 21272 9580
rect 21324 9568 21330 9580
rect 21324 9540 21680 9568
rect 21324 9528 21330 9540
rect 20901 9503 20959 9509
rect 20901 9469 20913 9503
rect 20947 9500 20959 9503
rect 21545 9503 21603 9509
rect 21545 9500 21557 9503
rect 20947 9472 21557 9500
rect 20947 9469 20959 9472
rect 20901 9463 20959 9469
rect 21545 9469 21557 9472
rect 21591 9469 21603 9503
rect 21652 9500 21680 9540
rect 22002 9528 22008 9580
rect 22060 9528 22066 9580
rect 22112 9500 22140 9676
rect 22738 9664 22744 9676
rect 22796 9664 22802 9716
rect 23014 9704 23020 9716
rect 22848 9676 23020 9704
rect 22848 9645 22876 9676
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 24854 9664 24860 9716
rect 24912 9664 24918 9716
rect 25038 9664 25044 9716
rect 25096 9664 25102 9716
rect 25225 9707 25283 9713
rect 25225 9673 25237 9707
rect 25271 9704 25283 9707
rect 25498 9704 25504 9716
rect 25271 9676 25504 9704
rect 25271 9673 25283 9676
rect 25225 9667 25283 9673
rect 25498 9664 25504 9676
rect 25556 9664 25562 9716
rect 22833 9639 22891 9645
rect 22833 9605 22845 9639
rect 22879 9605 22891 9639
rect 22833 9599 22891 9605
rect 23566 9596 23572 9648
rect 23624 9596 23630 9648
rect 24872 9636 24900 9664
rect 24780 9608 24900 9636
rect 25056 9636 25084 9664
rect 25317 9639 25375 9645
rect 25317 9636 25329 9639
rect 25056 9608 25329 9636
rect 24780 9577 24808 9608
rect 25317 9605 25329 9608
rect 25363 9605 25375 9639
rect 25317 9599 25375 9605
rect 24765 9571 24823 9577
rect 24765 9568 24777 9571
rect 24228 9540 24777 9568
rect 21652 9472 22140 9500
rect 22189 9503 22247 9509
rect 21545 9463 21603 9469
rect 22189 9469 22201 9503
rect 22235 9469 22247 9503
rect 22189 9463 22247 9469
rect 22204 9432 22232 9463
rect 22554 9460 22560 9512
rect 22612 9460 22618 9512
rect 22830 9500 22836 9512
rect 22664 9472 22836 9500
rect 22664 9432 22692 9472
rect 22830 9460 22836 9472
rect 22888 9460 22894 9512
rect 20588 9404 22692 9432
rect 20588 9392 20594 9404
rect 17862 9364 17868 9376
rect 17604 9336 17868 9364
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 21453 9367 21511 9373
rect 21453 9333 21465 9367
rect 21499 9364 21511 9367
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 21499 9336 21833 9364
rect 21499 9333 21511 9336
rect 21453 9327 21511 9333
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 21821 9327 21879 9333
rect 22922 9324 22928 9376
rect 22980 9364 22986 9376
rect 24228 9364 24256 9540
rect 24765 9537 24777 9540
rect 24811 9537 24823 9571
rect 24765 9531 24823 9537
rect 24854 9528 24860 9580
rect 24912 9528 24918 9580
rect 24673 9503 24731 9509
rect 24673 9469 24685 9503
rect 24719 9469 24731 9503
rect 24673 9463 24731 9469
rect 22980 9336 24256 9364
rect 22980 9324 22986 9336
rect 24302 9324 24308 9376
rect 24360 9324 24366 9376
rect 24688 9364 24716 9463
rect 25866 9460 25872 9512
rect 25924 9460 25930 9512
rect 24946 9364 24952 9376
rect 24688 9336 24952 9364
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 1104 9274 26496 9296
rect 1104 9222 4124 9274
rect 4176 9222 4188 9274
rect 4240 9222 4252 9274
rect 4304 9222 4316 9274
rect 4368 9222 4380 9274
rect 4432 9222 10472 9274
rect 10524 9222 10536 9274
rect 10588 9222 10600 9274
rect 10652 9222 10664 9274
rect 10716 9222 10728 9274
rect 10780 9222 16820 9274
rect 16872 9222 16884 9274
rect 16936 9222 16948 9274
rect 17000 9222 17012 9274
rect 17064 9222 17076 9274
rect 17128 9222 23168 9274
rect 23220 9222 23232 9274
rect 23284 9222 23296 9274
rect 23348 9222 23360 9274
rect 23412 9222 23424 9274
rect 23476 9222 26496 9274
rect 1104 9200 26496 9222
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 5902 9160 5908 9172
rect 4019 9132 5908 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 8202 9160 8208 9172
rect 7208 9132 8208 9160
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 7006 9024 7012 9036
rect 4212 8996 4660 9024
rect 4212 8984 4218 8996
rect 3510 8916 3516 8968
rect 3568 8916 3574 8968
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 4120 8928 4445 8956
rect 4120 8916 4126 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4522 8916 4528 8968
rect 4580 8916 4586 8968
rect 4632 8965 4660 8996
rect 6104 8996 7012 9024
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 3941 8891 3999 8897
rect 3941 8888 3953 8891
rect 3712 8860 3953 8888
rect 3712 8832 3740 8860
rect 3941 8857 3953 8860
rect 3987 8857 3999 8891
rect 3941 8851 3999 8857
rect 4157 8891 4215 8897
rect 4157 8857 4169 8891
rect 4203 8888 4215 8891
rect 6104 8888 6132 8996
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7208 9033 7236 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 10137 9163 10195 9169
rect 10137 9160 10149 9163
rect 9732 9132 10149 9160
rect 9732 9120 9738 9132
rect 10137 9129 10149 9132
rect 10183 9129 10195 9163
rect 10137 9123 10195 9129
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9160 12495 9163
rect 12802 9160 12808 9172
rect 12483 9132 12808 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 15470 9120 15476 9172
rect 15528 9120 15534 9172
rect 18414 9120 18420 9172
rect 18472 9160 18478 9172
rect 18785 9163 18843 9169
rect 18785 9160 18797 9163
rect 18472 9132 18797 9160
rect 18472 9120 18478 9132
rect 18785 9129 18797 9132
rect 18831 9129 18843 9163
rect 18785 9123 18843 9129
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 22143 9163 22201 9169
rect 22143 9160 22155 9163
rect 22060 9132 22155 9160
rect 22060 9120 22066 9132
rect 22143 9129 22155 9132
rect 22189 9129 22201 9163
rect 22143 9123 22201 9129
rect 23014 9120 23020 9172
rect 23072 9160 23078 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 23072 9132 23305 9160
rect 23072 9120 23078 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 24854 9160 24860 9172
rect 23293 9123 23351 9129
rect 24044 9132 24860 9160
rect 8021 9095 8079 9101
rect 8021 9061 8033 9095
rect 8067 9092 8079 9095
rect 11422 9092 11428 9104
rect 8067 9064 10824 9092
rect 8067 9061 8079 9064
rect 8021 9055 8079 9061
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 8993 7251 9027
rect 8113 9027 8171 9033
rect 8113 9024 8125 9027
rect 7193 8987 7251 8993
rect 7484 8996 8125 9024
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 4203 8860 6132 8888
rect 4203 8857 4215 8860
rect 4157 8851 4215 8857
rect 6178 8848 6184 8900
rect 6236 8848 6242 8900
rect 6472 8888 6500 8919
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 6733 8959 6791 8965
rect 6733 8956 6745 8959
rect 6604 8928 6745 8956
rect 6604 8916 6610 8928
rect 6733 8925 6745 8928
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 7484 8965 7512 8996
rect 8113 8993 8125 8996
rect 8159 8993 8171 9027
rect 8113 8987 8171 8993
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 10796 9033 10824 9064
rect 11256 9064 11428 9092
rect 10781 9027 10839 9033
rect 8260 8996 9628 9024
rect 8260 8984 8266 8996
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 7834 8916 7840 8968
rect 7892 8916 7898 8968
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8956 8965 8984 8996
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 8076 8928 8677 8956
rect 8076 8916 8082 8928
rect 8665 8925 8677 8928
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9447 8928 9505 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9600 8956 9628 8996
rect 10781 8993 10793 9027
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 10962 8956 10968 8968
rect 9600 8928 10968 8956
rect 9493 8919 9551 8925
rect 6932 8888 6960 8916
rect 6472 8860 6960 8888
rect 7653 8891 7711 8897
rect 7653 8857 7665 8891
rect 7699 8857 7711 8891
rect 7653 8851 7711 8857
rect 7745 8891 7803 8897
rect 7745 8857 7757 8891
rect 7791 8888 7803 8891
rect 8294 8888 8300 8900
rect 7791 8860 8300 8888
rect 7791 8857 7803 8860
rect 7745 8851 7803 8857
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 2961 8823 3019 8829
rect 2961 8820 2973 8823
rect 2924 8792 2973 8820
rect 2924 8780 2930 8792
rect 2961 8789 2973 8792
rect 3007 8789 3019 8823
rect 2961 8783 3019 8789
rect 3694 8780 3700 8832
rect 3752 8780 3758 8832
rect 3786 8780 3792 8832
rect 3844 8780 3850 8832
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4706 8820 4712 8832
rect 4295 8792 4712 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 7668 8820 7696 8851
rect 8294 8848 8300 8860
rect 8352 8888 8358 8900
rect 9033 8891 9091 8897
rect 9033 8888 9045 8891
rect 8352 8860 9045 8888
rect 8352 8848 8358 8860
rect 9033 8857 9045 8860
rect 9079 8857 9091 8891
rect 9232 8888 9260 8919
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11054 8916 11060 8968
rect 11112 8916 11118 8968
rect 11256 8965 11284 9064
rect 11422 9052 11428 9064
rect 11480 9092 11486 9104
rect 13078 9092 13084 9104
rect 11480 9064 13084 9092
rect 11480 9052 11486 9064
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 15102 9092 15108 9104
rect 14108 9064 15108 9092
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11882 9024 11888 9036
rect 11388 8996 11888 9024
rect 11388 8984 11394 8996
rect 11882 8984 11888 8996
rect 11940 9024 11946 9036
rect 14108 9024 14136 9064
rect 15102 9052 15108 9064
rect 15160 9052 15166 9104
rect 23201 9095 23259 9101
rect 23201 9061 23213 9095
rect 23247 9092 23259 9095
rect 24044 9092 24072 9132
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 23247 9064 24072 9092
rect 23247 9061 23259 9064
rect 23201 9055 23259 9061
rect 11940 8996 14136 9024
rect 11940 8984 11946 8996
rect 14182 8984 14188 9036
rect 14240 8984 14246 9036
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 14332 8996 14381 9024
rect 14332 8984 14338 8996
rect 14369 8993 14381 8996
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 16114 8984 16120 9036
rect 16172 8984 16178 9036
rect 20530 9024 20536 9036
rect 17880 8996 20536 9024
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 11756 8928 12081 8956
rect 11756 8916 11762 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 13265 8959 13323 8965
rect 13265 8956 13277 8959
rect 12860 8928 13277 8956
rect 12860 8916 12866 8928
rect 13265 8925 13277 8928
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8956 15899 8959
rect 17880 8956 17908 8996
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 22649 9027 22707 9033
rect 22649 8993 22661 9027
rect 22695 9024 22707 9027
rect 23474 9024 23480 9036
rect 22695 8996 23480 9024
rect 22695 8993 22707 8996
rect 22649 8987 22707 8993
rect 23474 8984 23480 8996
rect 23532 9024 23538 9036
rect 23934 9024 23940 9036
rect 23532 8996 23940 9024
rect 23532 8984 23538 8996
rect 23934 8984 23940 8996
rect 23992 9024 23998 9036
rect 24302 9024 24308 9036
rect 23992 8996 24308 9024
rect 23992 8984 23998 8996
rect 24302 8984 24308 8996
rect 24360 8984 24366 9036
rect 24673 9027 24731 9033
rect 24673 8993 24685 9027
rect 24719 9024 24731 9027
rect 25314 9024 25320 9036
rect 24719 8996 25320 9024
rect 24719 8993 24731 8996
rect 24673 8987 24731 8993
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 15887 8928 17908 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18693 8959 18751 8965
rect 18693 8956 18705 8959
rect 18012 8928 18705 8956
rect 18012 8916 18018 8928
rect 18693 8925 18705 8928
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8956 18843 8959
rect 18874 8956 18880 8968
rect 18831 8928 18880 8956
rect 18831 8925 18843 8928
rect 18785 8919 18843 8925
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 18969 8959 19027 8965
rect 18969 8925 18981 8959
rect 19015 8925 19027 8959
rect 18969 8919 19027 8925
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8956 20407 8959
rect 20622 8956 20628 8968
rect 20395 8928 20628 8956
rect 20395 8925 20407 8928
rect 20349 8919 20407 8925
rect 10042 8888 10048 8900
rect 9232 8860 10048 8888
rect 9033 8851 9091 8857
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 12158 8888 12164 8900
rect 11440 8860 12164 8888
rect 6880 8792 7696 8820
rect 6880 8780 6886 8792
rect 10226 8780 10232 8832
rect 10284 8780 10290 8832
rect 11440 8829 11468 8860
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12621 8891 12679 8897
rect 12621 8857 12633 8891
rect 12667 8888 12679 8891
rect 13078 8888 13084 8900
rect 12667 8860 13084 8888
rect 12667 8857 12679 8860
rect 12621 8851 12679 8857
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 17862 8848 17868 8900
rect 17920 8848 17926 8900
rect 18984 8888 19012 8919
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 20714 8916 20720 8968
rect 20772 8916 20778 8968
rect 22830 8916 22836 8968
rect 22888 8956 22894 8968
rect 22925 8959 22983 8965
rect 22925 8956 22937 8959
rect 22888 8928 22937 8956
rect 22888 8916 22894 8928
rect 22925 8925 22937 8928
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 23017 8959 23075 8965
rect 23017 8925 23029 8959
rect 23063 8956 23075 8959
rect 23566 8956 23572 8968
rect 23063 8928 23572 8956
rect 23063 8925 23075 8928
rect 23017 8919 23075 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 23658 8916 23664 8968
rect 23716 8916 23722 8968
rect 23750 8916 23756 8968
rect 23808 8956 23814 8968
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 23808 8928 24409 8956
rect 23808 8916 23814 8928
rect 24397 8925 24409 8928
rect 24443 8925 24455 8959
rect 24397 8919 24455 8925
rect 18984 8860 20484 8888
rect 20456 8832 20484 8860
rect 21542 8848 21548 8900
rect 21600 8848 21606 8900
rect 23584 8888 23612 8916
rect 23842 8888 23848 8900
rect 22066 8860 23336 8888
rect 23584 8860 23848 8888
rect 11425 8823 11483 8829
rect 11425 8789 11437 8823
rect 11471 8789 11483 8823
rect 11425 8783 11483 8789
rect 11517 8823 11575 8829
rect 11517 8789 11529 8823
rect 11563 8820 11575 8823
rect 11606 8820 11612 8832
rect 11563 8792 11612 8820
rect 11563 8789 11575 8792
rect 11517 8783 11575 8789
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 12032 8792 12265 8820
rect 12032 8780 12038 8792
rect 12253 8789 12265 8792
rect 12299 8789 12311 8823
rect 12253 8783 12311 8789
rect 12421 8823 12479 8829
rect 12421 8789 12433 8823
rect 12467 8820 12479 8823
rect 12526 8820 12532 8832
rect 12467 8792 12532 8820
rect 12467 8789 12479 8792
rect 12421 8783 12479 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 12710 8780 12716 8832
rect 12768 8780 12774 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 14461 8823 14519 8829
rect 14461 8820 14473 8823
rect 12952 8792 14473 8820
rect 12952 8780 12958 8792
rect 14461 8789 14473 8792
rect 14507 8789 14519 8823
rect 14461 8783 14519 8789
rect 14826 8780 14832 8832
rect 14884 8780 14890 8832
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 17402 8820 17408 8832
rect 15988 8792 17408 8820
rect 15988 8780 15994 8792
rect 17402 8780 17408 8792
rect 17460 8780 17466 8832
rect 20438 8780 20444 8832
rect 20496 8820 20502 8832
rect 22066 8820 22094 8860
rect 20496 8792 22094 8820
rect 22833 8823 22891 8829
rect 20496 8780 20502 8792
rect 22833 8789 22845 8823
rect 22879 8820 22891 8823
rect 23198 8820 23204 8832
rect 22879 8792 23204 8820
rect 22879 8789 22891 8792
rect 22833 8783 22891 8789
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 23308 8820 23336 8860
rect 23842 8848 23848 8860
rect 23900 8848 23906 8900
rect 24026 8848 24032 8900
rect 24084 8888 24090 8900
rect 24670 8888 24676 8900
rect 24084 8860 24676 8888
rect 24084 8848 24090 8860
rect 24670 8848 24676 8860
rect 24728 8888 24734 8900
rect 24728 8860 25162 8888
rect 24728 8848 24734 8860
rect 23566 8820 23572 8832
rect 23308 8792 23572 8820
rect 23566 8780 23572 8792
rect 23624 8780 23630 8832
rect 23753 8823 23811 8829
rect 23753 8789 23765 8823
rect 23799 8820 23811 8823
rect 24302 8820 24308 8832
rect 23799 8792 24308 8820
rect 23799 8789 23811 8792
rect 23753 8783 23811 8789
rect 24302 8780 24308 8792
rect 24360 8780 24366 8832
rect 24946 8780 24952 8832
rect 25004 8820 25010 8832
rect 26145 8823 26203 8829
rect 26145 8820 26157 8823
rect 25004 8792 26157 8820
rect 25004 8780 25010 8792
rect 26145 8789 26157 8792
rect 26191 8789 26203 8823
rect 26145 8783 26203 8789
rect 1104 8730 26656 8752
rect 1104 8678 7298 8730
rect 7350 8678 7362 8730
rect 7414 8678 7426 8730
rect 7478 8678 7490 8730
rect 7542 8678 7554 8730
rect 7606 8678 13646 8730
rect 13698 8678 13710 8730
rect 13762 8678 13774 8730
rect 13826 8678 13838 8730
rect 13890 8678 13902 8730
rect 13954 8678 19994 8730
rect 20046 8678 20058 8730
rect 20110 8678 20122 8730
rect 20174 8678 20186 8730
rect 20238 8678 20250 8730
rect 20302 8678 26342 8730
rect 26394 8678 26406 8730
rect 26458 8678 26470 8730
rect 26522 8678 26534 8730
rect 26586 8678 26598 8730
rect 26650 8678 26656 8730
rect 1104 8656 26656 8678
rect 3878 8616 3884 8628
rect 3344 8588 3884 8616
rect 3344 8548 3372 8588
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 4341 8619 4399 8625
rect 4341 8585 4353 8619
rect 4387 8616 4399 8619
rect 4522 8616 4528 8628
rect 4387 8588 4528 8616
rect 4387 8585 4399 8588
rect 4341 8579 4399 8585
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8018 8616 8024 8628
rect 7975 8588 8024 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 9490 8576 9496 8628
rect 9548 8576 9554 8628
rect 10226 8576 10232 8628
rect 10284 8576 10290 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10928 8588 10977 8616
rect 10928 8576 10934 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 11480 8588 11744 8616
rect 11480 8576 11486 8588
rect 4062 8548 4068 8560
rect 4120 8557 4126 8560
rect 4120 8551 4149 8557
rect 2898 8520 3372 8548
rect 3436 8520 4068 8548
rect 3436 8492 3464 8520
rect 4062 8508 4068 8520
rect 4137 8517 4149 8551
rect 4120 8511 4149 8517
rect 5445 8551 5503 8557
rect 5445 8517 5457 8551
rect 5491 8548 5503 8551
rect 5534 8548 5540 8560
rect 5491 8520 5540 8548
rect 5491 8517 5503 8520
rect 5445 8511 5503 8517
rect 4120 8508 4126 8511
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8548 6239 8551
rect 7285 8551 7343 8557
rect 7285 8548 7297 8551
rect 6227 8520 7297 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 7285 8517 7297 8520
rect 7331 8548 7343 8551
rect 8110 8548 8116 8560
rect 7331 8520 8116 8548
rect 7331 8517 7343 8520
rect 7285 8511 7343 8517
rect 8110 8508 8116 8520
rect 8168 8508 8174 8560
rect 9398 8548 9404 8560
rect 8970 8520 9404 8548
rect 9398 8508 9404 8520
rect 9456 8508 9462 8560
rect 9508 8548 9536 8576
rect 9508 8520 9720 8548
rect 3418 8440 3424 8492
rect 3476 8440 3482 8492
rect 3510 8440 3516 8492
rect 3568 8440 3574 8492
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 3789 8483 3847 8489
rect 3789 8480 3801 8483
rect 3660 8452 3801 8480
rect 3660 8440 3666 8452
rect 3789 8449 3801 8452
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 1412 8276 1440 8375
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 3528 8344 3556 8440
rect 3896 8412 3924 8443
rect 3712 8384 3924 8412
rect 3712 8356 3740 8384
rect 3605 8347 3663 8353
rect 3605 8344 3617 8347
rect 3528 8316 3617 8344
rect 3605 8313 3617 8316
rect 3651 8313 3663 8347
rect 3605 8307 3663 8313
rect 3694 8304 3700 8356
rect 3752 8304 3758 8356
rect 3988 8344 4016 8443
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6822 8480 6828 8492
rect 5960 8452 6828 8480
rect 5960 8440 5966 8452
rect 6822 8440 6828 8452
rect 6880 8480 6886 8492
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 6880 8452 7573 8480
rect 6880 8440 6886 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8480 7895 8483
rect 7926 8480 7932 8492
rect 7883 8452 7932 8480
rect 7883 8449 7895 8452
rect 7837 8443 7895 8449
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 9692 8489 9720 8520
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4522 8412 4528 8424
rect 4295 8384 4528 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 4982 8372 4988 8424
rect 5040 8372 5046 8424
rect 6546 8372 6552 8424
rect 6604 8372 6610 8424
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8412 9459 8415
rect 10244 8412 10272 8576
rect 11606 8548 11612 8560
rect 10888 8520 11612 8548
rect 10888 8489 10916 8520
rect 11606 8508 11612 8520
rect 11664 8508 11670 8560
rect 11716 8548 11744 8588
rect 11790 8576 11796 8628
rect 11848 8616 11854 8628
rect 11977 8619 12035 8625
rect 11977 8616 11989 8619
rect 11848 8588 11989 8616
rect 11848 8576 11854 8588
rect 11977 8585 11989 8588
rect 12023 8585 12035 8619
rect 11977 8579 12035 8585
rect 12544 8588 12756 8616
rect 12544 8548 12572 8588
rect 12728 8560 12756 8588
rect 13262 8576 13268 8628
rect 13320 8576 13326 8628
rect 14918 8576 14924 8628
rect 14976 8576 14982 8628
rect 15378 8576 15384 8628
rect 15436 8576 15442 8628
rect 15930 8616 15936 8628
rect 15856 8588 15936 8616
rect 11716 8520 12204 8548
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8480 11207 8483
rect 11885 8483 11943 8489
rect 11195 8452 11652 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 9447 8384 10272 8412
rect 10781 8415 10839 8421
rect 9447 8381 9459 8384
rect 9401 8375 9459 8381
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11054 8412 11060 8424
rect 10827 8384 11060 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11054 8372 11060 8384
rect 11112 8412 11118 8424
rect 11333 8415 11391 8421
rect 11333 8412 11345 8415
rect 11112 8384 11345 8412
rect 11112 8372 11118 8384
rect 11333 8381 11345 8384
rect 11379 8381 11391 8415
rect 11333 8375 11391 8381
rect 11146 8344 11152 8356
rect 3896 8316 4016 8344
rect 9600 8316 11152 8344
rect 1854 8276 1860 8288
rect 1412 8248 1860 8276
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 3145 8279 3203 8285
rect 3145 8245 3157 8279
rect 3191 8276 3203 8279
rect 3326 8276 3332 8288
rect 3191 8248 3332 8276
rect 3191 8245 3203 8248
rect 3145 8239 3203 8245
rect 3326 8236 3332 8248
rect 3384 8276 3390 8288
rect 3896 8276 3924 8316
rect 3384 8248 3924 8276
rect 3384 8236 3390 8248
rect 7282 8236 7288 8288
rect 7340 8276 7346 8288
rect 7377 8279 7435 8285
rect 7377 8276 7389 8279
rect 7340 8248 7389 8276
rect 7340 8236 7346 8248
rect 7377 8245 7389 8248
rect 7423 8245 7435 8279
rect 7377 8239 7435 8245
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9600 8276 9628 8316
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 8812 8248 9628 8276
rect 11348 8276 11376 8375
rect 11514 8372 11520 8424
rect 11572 8372 11578 8424
rect 11624 8412 11652 8452
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12066 8480 12072 8492
rect 11931 8452 12072 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12176 8489 12204 8520
rect 12268 8520 12572 8548
rect 12268 8489 12296 8520
rect 12710 8508 12716 8560
rect 12768 8508 12774 8560
rect 15396 8548 15424 8576
rect 15856 8557 15884 8588
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 19981 8619 20039 8625
rect 19981 8585 19993 8619
rect 20027 8616 20039 8619
rect 20346 8616 20352 8628
rect 20027 8588 20352 8616
rect 20027 8585 20039 8588
rect 19981 8579 20039 8585
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 22554 8616 22560 8628
rect 20680 8588 22560 8616
rect 20680 8576 20686 8588
rect 22554 8576 22560 8588
rect 22612 8616 22618 8628
rect 23750 8616 23756 8628
rect 22612 8588 23756 8616
rect 22612 8576 22618 8588
rect 23750 8576 23756 8588
rect 23808 8576 23814 8628
rect 24026 8616 24032 8628
rect 23860 8588 24032 8616
rect 15841 8551 15899 8557
rect 15396 8520 15516 8548
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12434 8440 12440 8492
rect 12492 8440 12498 8492
rect 12621 8490 12679 8495
rect 12544 8489 12679 8490
rect 12544 8462 12633 8489
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11624 8384 11805 8412
rect 11793 8381 11805 8384
rect 11839 8412 11851 8415
rect 11974 8412 11980 8424
rect 11839 8384 11980 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12544 8412 12572 8462
rect 12621 8455 12633 8462
rect 12667 8455 12679 8489
rect 12621 8449 12679 8455
rect 12713 8473 12771 8479
rect 12713 8439 12725 8473
rect 12759 8439 12771 8473
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 15488 8489 15516 8520
rect 15841 8517 15853 8551
rect 15887 8517 15899 8551
rect 15841 8511 15899 8517
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8449 15255 8483
rect 15197 8443 15255 8449
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8449 15531 8483
rect 15856 8480 15884 8511
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 16080 8520 17264 8548
rect 16080 8508 16086 8520
rect 17236 8489 17264 8520
rect 20714 8508 20720 8560
rect 20772 8548 20778 8560
rect 20901 8551 20959 8557
rect 20901 8548 20913 8551
rect 20772 8520 20913 8548
rect 20772 8508 20778 8520
rect 20901 8517 20913 8520
rect 20947 8517 20959 8551
rect 20901 8511 20959 8517
rect 23474 8508 23480 8560
rect 23532 8548 23538 8560
rect 23569 8551 23627 8557
rect 23569 8548 23581 8551
rect 23532 8520 23581 8548
rect 23532 8508 23538 8520
rect 23569 8517 23581 8520
rect 23615 8517 23627 8551
rect 23860 8548 23888 8588
rect 24026 8576 24032 8588
rect 24084 8616 24090 8628
rect 25593 8619 25651 8625
rect 25593 8616 25605 8619
rect 24084 8588 25605 8616
rect 24084 8576 24090 8588
rect 25593 8585 25605 8588
rect 25639 8616 25651 8619
rect 25866 8616 25872 8628
rect 25639 8588 25872 8616
rect 25639 8585 25651 8588
rect 25593 8579 25651 8585
rect 25866 8576 25872 8588
rect 25924 8576 25930 8628
rect 23569 8511 23627 8517
rect 23676 8520 23888 8548
rect 24121 8551 24179 8557
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15856 8452 16129 8480
rect 15473 8443 15531 8449
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 16347 8452 16681 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 19981 8483 20039 8489
rect 19981 8449 19993 8483
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 12713 8433 12771 8439
rect 12084 8384 12572 8412
rect 11532 8344 11560 8372
rect 11885 8347 11943 8353
rect 11885 8344 11897 8347
rect 11532 8316 11897 8344
rect 11885 8313 11897 8316
rect 11931 8313 11943 8347
rect 11885 8307 11943 8313
rect 12084 8276 12112 8384
rect 12728 8356 12756 8433
rect 12250 8304 12256 8356
rect 12308 8344 12314 8356
rect 12345 8347 12403 8353
rect 12345 8344 12357 8347
rect 12308 8316 12357 8344
rect 12308 8304 12314 8316
rect 12345 8313 12357 8316
rect 12391 8313 12403 8347
rect 12345 8307 12403 8313
rect 12710 8304 12716 8356
rect 12768 8304 12774 8356
rect 15212 8344 15240 8443
rect 15396 8412 15424 8443
rect 17770 8412 17776 8424
rect 15396 8384 17776 8412
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 19702 8372 19708 8424
rect 19760 8372 19766 8424
rect 19996 8412 20024 8443
rect 20346 8440 20352 8492
rect 20404 8440 20410 8492
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 20993 8483 21051 8489
rect 20993 8449 21005 8483
rect 21039 8480 21051 8483
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21039 8452 21833 8480
rect 21039 8449 21051 8452
rect 20993 8443 21051 8449
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22925 8483 22983 8489
rect 22925 8449 22937 8483
rect 22971 8449 22983 8483
rect 22925 8443 22983 8449
rect 20824 8412 20852 8443
rect 21266 8412 21272 8424
rect 19996 8384 21272 8412
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 22370 8372 22376 8424
rect 22428 8372 22434 8424
rect 22940 8412 22968 8443
rect 23014 8440 23020 8492
rect 23072 8480 23078 8492
rect 23109 8483 23167 8489
rect 23109 8480 23121 8483
rect 23072 8452 23121 8480
rect 23072 8440 23078 8452
rect 23109 8449 23121 8452
rect 23155 8449 23167 8483
rect 23109 8443 23167 8449
rect 23198 8440 23204 8492
rect 23256 8480 23262 8492
rect 23676 8480 23704 8520
rect 24121 8517 24133 8551
rect 24167 8548 24179 8551
rect 24394 8548 24400 8560
rect 24167 8520 24400 8548
rect 24167 8517 24179 8520
rect 24121 8511 24179 8517
rect 24394 8508 24400 8520
rect 24452 8508 24458 8560
rect 24670 8508 24676 8560
rect 24728 8508 24734 8560
rect 23256 8452 23704 8480
rect 23256 8440 23262 8452
rect 23566 8412 23572 8424
rect 22940 8384 23572 8412
rect 23566 8372 23572 8384
rect 23624 8372 23630 8424
rect 23750 8372 23756 8424
rect 23808 8412 23814 8424
rect 23845 8415 23903 8421
rect 23845 8412 23857 8415
rect 23808 8384 23857 8412
rect 23808 8372 23814 8384
rect 23845 8381 23857 8384
rect 23891 8381 23903 8415
rect 24578 8412 24584 8424
rect 23845 8375 23903 8381
rect 23952 8384 24584 8412
rect 16114 8344 16120 8356
rect 15212 8316 16120 8344
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 19886 8304 19892 8356
rect 19944 8304 19950 8356
rect 20533 8347 20591 8353
rect 20533 8313 20545 8347
rect 20579 8344 20591 8347
rect 20806 8344 20812 8356
rect 20579 8316 20812 8344
rect 20579 8313 20591 8316
rect 20533 8307 20591 8313
rect 20806 8304 20812 8316
rect 20864 8304 20870 8356
rect 22922 8304 22928 8356
rect 22980 8344 22986 8356
rect 23017 8347 23075 8353
rect 23017 8344 23029 8347
rect 22980 8316 23029 8344
rect 22980 8304 22986 8316
rect 23017 8313 23029 8316
rect 23063 8313 23075 8347
rect 23952 8344 23980 8384
rect 24578 8372 24584 8384
rect 24636 8372 24642 8424
rect 24854 8372 24860 8424
rect 24912 8412 24918 8424
rect 24912 8384 25820 8412
rect 24912 8372 24918 8384
rect 25792 8356 25820 8384
rect 23017 8307 23075 8313
rect 23768 8316 23980 8344
rect 11348 8248 12112 8276
rect 8812 8236 8818 8248
rect 12802 8236 12808 8288
rect 12860 8236 12866 8288
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15657 8279 15715 8285
rect 15657 8276 15669 8279
rect 15344 8248 15669 8276
rect 15344 8236 15350 8248
rect 15657 8245 15669 8248
rect 15703 8245 15715 8279
rect 15657 8239 15715 8245
rect 16206 8236 16212 8288
rect 16264 8236 16270 8288
rect 16390 8236 16396 8288
rect 16448 8276 16454 8288
rect 18322 8276 18328 8288
rect 16448 8248 18328 8276
rect 16448 8236 16454 8248
rect 18322 8236 18328 8248
rect 18380 8236 18386 8288
rect 23569 8279 23627 8285
rect 23569 8245 23581 8279
rect 23615 8276 23627 8279
rect 23658 8276 23664 8288
rect 23615 8248 23664 8276
rect 23615 8245 23627 8248
rect 23569 8239 23627 8245
rect 23658 8236 23664 8248
rect 23716 8236 23722 8288
rect 23768 8285 23796 8316
rect 25774 8304 25780 8356
rect 25832 8304 25838 8356
rect 23753 8279 23811 8285
rect 23753 8245 23765 8279
rect 23799 8245 23811 8279
rect 23753 8239 23811 8245
rect 1104 8186 26496 8208
rect 1104 8134 4124 8186
rect 4176 8134 4188 8186
rect 4240 8134 4252 8186
rect 4304 8134 4316 8186
rect 4368 8134 4380 8186
rect 4432 8134 10472 8186
rect 10524 8134 10536 8186
rect 10588 8134 10600 8186
rect 10652 8134 10664 8186
rect 10716 8134 10728 8186
rect 10780 8134 16820 8186
rect 16872 8134 16884 8186
rect 16936 8134 16948 8186
rect 17000 8134 17012 8186
rect 17064 8134 17076 8186
rect 17128 8134 23168 8186
rect 23220 8134 23232 8186
rect 23284 8134 23296 8186
rect 23348 8134 23360 8186
rect 23412 8134 23424 8186
rect 23476 8134 26496 8186
rect 1104 8112 26496 8134
rect 3970 8032 3976 8084
rect 4028 8032 4034 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 13998 8072 14004 8084
rect 4120 8044 14004 8072
rect 4120 8032 4126 8044
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 16206 8072 16212 8084
rect 15396 8044 16212 8072
rect 4522 7964 4528 8016
rect 4580 7964 4586 8016
rect 10042 7964 10048 8016
rect 10100 7964 10106 8016
rect 12158 7964 12164 8016
rect 12216 8004 12222 8016
rect 12216 7976 13032 8004
rect 12216 7964 12222 7976
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2866 7936 2872 7948
rect 2179 7908 2872 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4540 7936 4568 7964
rect 4111 7908 4568 7936
rect 4801 7939 4859 7945
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 5442 7936 5448 7948
rect 4847 7908 5448 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 6733 7939 6791 7945
rect 6733 7936 6745 7939
rect 6604 7908 6745 7936
rect 6604 7896 6610 7908
rect 6733 7905 6745 7908
rect 6779 7936 6791 7939
rect 7098 7936 7104 7948
rect 6779 7908 7104 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8754 7936 8760 7948
rect 8352 7908 8760 7936
rect 8352 7896 8358 7908
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7936 10747 7939
rect 10870 7936 10876 7948
rect 10735 7908 10876 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 10870 7896 10876 7908
rect 10928 7936 10934 7948
rect 10928 7908 12940 7936
rect 10928 7896 10934 7908
rect 1854 7828 1860 7880
rect 1912 7828 1918 7880
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 2774 7760 2780 7812
rect 2832 7760 2838 7812
rect 3804 7800 3832 7831
rect 3970 7828 3976 7880
rect 4028 7828 4034 7880
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4540 7800 4568 7828
rect 3804 7772 4568 7800
rect 4632 7744 4660 7831
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 12032 7840 12633 7868
rect 12032 7828 12038 7840
rect 12621 7837 12633 7840
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 6914 7800 6920 7812
rect 6210 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 7009 7803 7067 7809
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 7282 7800 7288 7812
rect 7055 7772 7288 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 7282 7760 7288 7772
rect 7340 7760 7346 7812
rect 7650 7760 7656 7812
rect 7708 7760 7714 7812
rect 11149 7803 11207 7809
rect 11149 7769 11161 7803
rect 11195 7800 11207 7803
rect 11514 7800 11520 7812
rect 11195 7772 11520 7800
rect 11195 7769 11207 7772
rect 11149 7763 11207 7769
rect 11514 7760 11520 7772
rect 11572 7760 11578 7812
rect 12912 7800 12940 7908
rect 13004 7877 13032 7976
rect 13170 7964 13176 8016
rect 13228 8004 13234 8016
rect 14829 8007 14887 8013
rect 14829 8004 14841 8007
rect 13228 7976 14841 8004
rect 13228 7964 13234 7976
rect 13446 7896 13452 7948
rect 13504 7896 13510 7948
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13464 7800 13492 7896
rect 12912 7772 13492 7800
rect 14568 7800 14596 7976
rect 14829 7973 14841 7976
rect 14875 7973 14887 8007
rect 14829 7967 14887 7973
rect 15194 7936 15200 7948
rect 14660 7908 15200 7936
rect 14660 7877 14688 7908
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 15059 7840 15240 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 15105 7803 15163 7809
rect 15105 7800 15117 7803
rect 14568 7772 15117 7800
rect 15105 7769 15117 7772
rect 15151 7769 15163 7803
rect 15212 7800 15240 7840
rect 15286 7828 15292 7880
rect 15344 7828 15350 7880
rect 15396 7877 15424 8044
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 23014 8032 23020 8084
rect 23072 8072 23078 8084
rect 23293 8075 23351 8081
rect 23293 8072 23305 8075
rect 23072 8044 23305 8072
rect 23072 8032 23078 8044
rect 23293 8041 23305 8044
rect 23339 8041 23351 8075
rect 23293 8035 23351 8041
rect 23566 8032 23572 8084
rect 23624 8032 23630 8084
rect 19518 7964 19524 8016
rect 19576 8004 19582 8016
rect 19576 7976 20760 8004
rect 19576 7964 19582 7976
rect 15473 7939 15531 7945
rect 15473 7905 15485 7939
rect 15519 7936 15531 7939
rect 19886 7936 19892 7948
rect 15519 7908 17356 7936
rect 15519 7905 15531 7908
rect 15473 7899 15531 7905
rect 17328 7880 17356 7908
rect 19444 7908 19892 7936
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7837 15439 7871
rect 15381 7831 15439 7837
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18874 7868 18880 7880
rect 18831 7840 18880 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19444 7877 19472 7908
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 20622 7896 20628 7948
rect 20680 7896 20686 7948
rect 20732 7936 20760 7976
rect 22554 7936 22560 7948
rect 20732 7908 22560 7936
rect 22554 7896 22560 7908
rect 22612 7896 22618 7948
rect 24029 7939 24087 7945
rect 24029 7936 24041 7939
rect 23400 7908 24041 7936
rect 23400 7880 23428 7908
rect 24029 7905 24041 7908
rect 24075 7905 24087 7939
rect 24029 7899 24087 7905
rect 18969 7871 19027 7877
rect 18969 7837 18981 7871
rect 19015 7837 19027 7871
rect 18969 7831 19027 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 19794 7868 19800 7880
rect 19659 7840 19800 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 15654 7800 15660 7812
rect 15212 7772 15660 7800
rect 15105 7763 15163 7769
rect 15654 7760 15660 7772
rect 15712 7760 15718 7812
rect 15749 7803 15807 7809
rect 15749 7769 15761 7803
rect 15795 7769 15807 7803
rect 18690 7800 18696 7812
rect 16974 7772 18696 7800
rect 15749 7763 15807 7769
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 4614 7732 4620 7744
rect 3651 7704 4620 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 6595 7735 6653 7741
rect 6595 7701 6607 7735
rect 6641 7732 6653 7735
rect 7190 7732 7196 7744
rect 6641 7704 7196 7732
rect 6641 7701 6653 7704
rect 6595 7695 6653 7701
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 12066 7692 12072 7744
rect 12124 7692 12130 7744
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 12805 7735 12863 7741
rect 12805 7732 12817 7735
rect 12308 7704 12817 7732
rect 12308 7692 12314 7704
rect 12805 7701 12817 7704
rect 12851 7701 12863 7735
rect 12805 7695 12863 7701
rect 14550 7692 14556 7744
rect 14608 7692 14614 7744
rect 15203 7735 15261 7741
rect 15203 7701 15215 7735
rect 15249 7732 15261 7735
rect 15764 7732 15792 7763
rect 15249 7704 15792 7732
rect 15249 7701 15261 7704
rect 15203 7695 15261 7701
rect 16482 7692 16488 7744
rect 16540 7732 16546 7744
rect 17052 7732 17080 7772
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 18984 7800 19012 7831
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 23014 7828 23020 7880
rect 23072 7828 23078 7880
rect 23201 7871 23259 7877
rect 23201 7837 23213 7871
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 18984 7772 20760 7800
rect 20732 7744 20760 7772
rect 20806 7760 20812 7812
rect 20864 7800 20870 7812
rect 20901 7803 20959 7809
rect 20901 7800 20913 7803
rect 20864 7772 20913 7800
rect 20864 7760 20870 7772
rect 20901 7769 20913 7772
rect 20947 7769 20959 7803
rect 20901 7763 20959 7769
rect 21174 7760 21180 7812
rect 21232 7800 21238 7812
rect 23216 7800 23244 7831
rect 23382 7828 23388 7880
rect 23440 7828 23446 7880
rect 23753 7871 23811 7877
rect 23753 7837 23765 7871
rect 23799 7837 23811 7871
rect 23753 7831 23811 7837
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7837 23903 7871
rect 23845 7831 23903 7837
rect 21232 7772 21390 7800
rect 22388 7772 23244 7800
rect 21232 7760 21238 7772
rect 16540 7704 17080 7732
rect 17221 7735 17279 7741
rect 16540 7692 16546 7704
rect 17221 7701 17233 7735
rect 17267 7732 17279 7735
rect 17402 7732 17408 7744
rect 17267 7704 17408 7732
rect 17267 7701 17279 7704
rect 17221 7695 17279 7701
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 17678 7692 17684 7744
rect 17736 7732 17742 7744
rect 18877 7735 18935 7741
rect 18877 7732 18889 7735
rect 17736 7704 18889 7732
rect 17736 7692 17742 7704
rect 18877 7701 18889 7704
rect 18923 7701 18935 7735
rect 18877 7695 18935 7701
rect 19245 7735 19303 7741
rect 19245 7701 19257 7735
rect 19291 7732 19303 7735
rect 19334 7732 19340 7744
rect 19291 7704 19340 7732
rect 19291 7701 19303 7704
rect 19245 7695 19303 7701
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 20714 7692 20720 7744
rect 20772 7692 20778 7744
rect 21284 7732 21312 7772
rect 22388 7744 22416 7772
rect 22186 7732 22192 7744
rect 21284 7704 22192 7732
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22370 7692 22376 7744
rect 22428 7692 22434 7744
rect 22462 7692 22468 7744
rect 22520 7692 22526 7744
rect 23768 7732 23796 7831
rect 23860 7800 23888 7831
rect 23934 7828 23940 7880
rect 23992 7828 23998 7880
rect 24026 7800 24032 7812
rect 23860 7772 24032 7800
rect 24026 7760 24032 7772
rect 24084 7760 24090 7812
rect 23842 7732 23848 7744
rect 23768 7704 23848 7732
rect 23842 7692 23848 7704
rect 23900 7732 23906 7744
rect 24210 7732 24216 7744
rect 23900 7704 24216 7732
rect 23900 7692 23906 7704
rect 24210 7692 24216 7704
rect 24268 7692 24274 7744
rect 1104 7642 26656 7664
rect 1104 7590 7298 7642
rect 7350 7590 7362 7642
rect 7414 7590 7426 7642
rect 7478 7590 7490 7642
rect 7542 7590 7554 7642
rect 7606 7590 13646 7642
rect 13698 7590 13710 7642
rect 13762 7590 13774 7642
rect 13826 7590 13838 7642
rect 13890 7590 13902 7642
rect 13954 7590 19994 7642
rect 20046 7590 20058 7642
rect 20110 7590 20122 7642
rect 20174 7590 20186 7642
rect 20238 7590 20250 7642
rect 20302 7590 26342 7642
rect 26394 7590 26406 7642
rect 26458 7590 26470 7642
rect 26522 7590 26534 7642
rect 26586 7590 26598 7642
rect 26650 7590 26656 7642
rect 1104 7568 26656 7590
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 1728 7500 2145 7528
rect 1728 7488 1734 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 2133 7491 2191 7497
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3786 7528 3792 7540
rect 3099 7500 3792 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 7098 7528 7104 7540
rect 4172 7500 7104 7528
rect 3878 7420 3884 7472
rect 3936 7420 3942 7472
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 3145 7395 3203 7401
rect 2363 7364 2728 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2700 7265 2728 7364
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 3510 7392 3516 7404
rect 3191 7364 3516 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 4172 7401 4200 7500
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 10597 7531 10655 7537
rect 10597 7528 10609 7531
rect 9732 7500 10609 7528
rect 9732 7488 9738 7500
rect 10597 7497 10609 7500
rect 10643 7497 10655 7531
rect 10597 7491 10655 7497
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 12066 7528 12072 7540
rect 12023 7500 12072 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 12802 7528 12808 7540
rect 12636 7500 12808 7528
rect 4433 7463 4491 7469
rect 4433 7429 4445 7463
rect 4479 7460 4491 7463
rect 4706 7460 4712 7472
rect 4479 7432 4712 7460
rect 4479 7429 4491 7432
rect 4433 7423 4491 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 6914 7460 6920 7472
rect 5658 7432 6920 7460
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 9692 7460 9720 7488
rect 9614 7432 9720 7460
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 12636 7460 12664 7500
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 14550 7528 14556 7540
rect 14016 7500 14556 7528
rect 9824 7432 10548 7460
rect 9824 7420 9830 7432
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 5902 7352 5908 7404
rect 5960 7392 5966 7404
rect 10520 7401 10548 7432
rect 12084 7432 12664 7460
rect 12084 7401 12112 7432
rect 12710 7420 12716 7472
rect 12768 7420 12774 7472
rect 14016 7460 14044 7500
rect 14550 7488 14556 7500
rect 14608 7528 14614 7540
rect 14608 7500 15792 7528
rect 14608 7488 14614 7500
rect 15764 7460 15792 7500
rect 16022 7488 16028 7540
rect 16080 7537 16086 7540
rect 16080 7531 16129 7537
rect 16080 7497 16083 7531
rect 16117 7497 16129 7531
rect 16080 7491 16129 7497
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 19518 7528 19524 7540
rect 17635 7500 19524 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 16080 7488 16086 7491
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 19613 7531 19671 7537
rect 19613 7497 19625 7531
rect 19659 7528 19671 7531
rect 19886 7528 19892 7540
rect 19659 7500 19892 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 20346 7488 20352 7540
rect 20404 7488 20410 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 20717 7531 20775 7537
rect 20717 7528 20729 7531
rect 20588 7500 20729 7528
rect 20588 7488 20594 7500
rect 20717 7497 20729 7500
rect 20763 7497 20775 7531
rect 20717 7491 20775 7497
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 21266 7528 21272 7540
rect 20864 7500 21272 7528
rect 20864 7488 20870 7500
rect 21266 7488 21272 7500
rect 21324 7528 21330 7540
rect 23293 7531 23351 7537
rect 21324 7500 22094 7528
rect 21324 7488 21330 7500
rect 16482 7460 16488 7472
rect 13938 7432 14044 7460
rect 15686 7432 16488 7460
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 18690 7420 18696 7472
rect 18748 7420 18754 7472
rect 20073 7463 20131 7469
rect 20073 7429 20085 7463
rect 20119 7460 20131 7463
rect 20548 7460 20576 7488
rect 20119 7432 20576 7460
rect 20119 7429 20131 7432
rect 20073 7423 20131 7429
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5960 7364 6009 7392
rect 5960 7352 5966 7364
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6181 7395 6239 7401
rect 6181 7361 6193 7395
rect 6227 7392 6239 7395
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6227 7364 7389 7392
rect 6227 7361 6239 7364
rect 6181 7355 6239 7361
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 4890 7324 4896 7336
rect 3384 7296 4896 7324
rect 3384 7284 3390 7296
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5224 7296 6101 7324
rect 5224 7284 5230 7296
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 2685 7259 2743 7265
rect 2685 7225 2697 7259
rect 2731 7225 2743 7259
rect 2685 7219 2743 7225
rect 7944 7200 7972 7287
rect 10042 7284 10048 7336
rect 10100 7284 10106 7336
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7293 10379 7327
rect 10520 7324 10548 7355
rect 16114 7352 16120 7404
rect 16172 7392 16178 7404
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 16172 7364 17233 7392
rect 16172 7352 16178 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 19889 7395 19947 7401
rect 19889 7392 19901 7395
rect 17221 7355 17279 7361
rect 19812 7364 19901 7392
rect 10520 7296 12204 7324
rect 10321 7287 10379 7293
rect 10336 7256 10364 7287
rect 11514 7256 11520 7268
rect 10336 7228 11520 7256
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3605 7191 3663 7197
rect 3605 7188 3617 7191
rect 2832 7160 3617 7188
rect 2832 7148 2838 7160
rect 3605 7157 3617 7160
rect 3651 7157 3663 7191
rect 3605 7151 3663 7157
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5040 7160 5917 7188
rect 5040 7148 5046 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 5905 7151 5963 7157
rect 7926 7148 7932 7200
rect 7984 7188 7990 7200
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 7984 7160 8585 7188
rect 7984 7148 7990 7160
rect 8573 7157 8585 7160
rect 8619 7188 8631 7191
rect 9490 7188 9496 7200
rect 8619 7160 9496 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 11606 7148 11612 7200
rect 11664 7148 11670 7200
rect 12176 7188 12204 7296
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 12492 7296 14289 7324
rect 12492 7284 12498 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7324 14703 7327
rect 16022 7324 16028 7336
rect 14691 7296 16028 7324
rect 14691 7293 14703 7296
rect 14645 7287 14703 7293
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 17310 7284 17316 7336
rect 17368 7324 17374 7336
rect 17862 7324 17868 7336
rect 17368 7296 17868 7324
rect 17368 7284 17374 7296
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 18141 7327 18199 7333
rect 18141 7293 18153 7327
rect 18187 7324 18199 7327
rect 19705 7327 19763 7333
rect 19705 7324 19717 7327
rect 18187 7296 19717 7324
rect 18187 7293 18199 7296
rect 18141 7287 18199 7293
rect 19705 7293 19717 7296
rect 19751 7293 19763 7327
rect 19705 7287 19763 7293
rect 17770 7216 17776 7268
rect 17828 7216 17834 7268
rect 12894 7188 12900 7200
rect 12176 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 14182 7148 14188 7200
rect 14240 7148 14246 7200
rect 17586 7148 17592 7200
rect 17644 7148 17650 7200
rect 18874 7148 18880 7200
rect 18932 7188 18938 7200
rect 19812 7188 19840 7364
rect 19889 7361 19901 7364
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 20165 7395 20223 7401
rect 20165 7361 20177 7395
rect 20211 7361 20223 7395
rect 21177 7395 21235 7401
rect 21177 7392 21189 7395
rect 20165 7355 20223 7361
rect 20916 7364 21189 7392
rect 20180 7256 20208 7355
rect 20806 7256 20812 7268
rect 20180 7228 20812 7256
rect 20806 7216 20812 7228
rect 20864 7216 20870 7268
rect 20916 7188 20944 7364
rect 21177 7361 21189 7364
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21818 7392 21824 7404
rect 21407 7364 21824 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21818 7352 21824 7364
rect 21876 7352 21882 7404
rect 22066 7392 22094 7500
rect 23293 7497 23305 7531
rect 23339 7528 23351 7531
rect 23382 7528 23388 7540
rect 23339 7500 23388 7528
rect 23339 7497 23351 7500
rect 23293 7491 23351 7497
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 24210 7488 24216 7540
rect 24268 7488 24274 7540
rect 24302 7488 24308 7540
rect 24360 7528 24366 7540
rect 24578 7528 24584 7540
rect 24360 7500 24584 7528
rect 24360 7488 24366 7500
rect 24578 7488 24584 7500
rect 24636 7488 24642 7540
rect 23400 7460 23428 7488
rect 24121 7463 24179 7469
rect 24121 7460 24133 7463
rect 22940 7432 23704 7460
rect 22646 7392 22652 7404
rect 22066 7364 22652 7392
rect 22646 7352 22652 7364
rect 22704 7392 22710 7404
rect 22940 7401 22968 7432
rect 22925 7395 22983 7401
rect 22704 7364 22876 7392
rect 22704 7352 22710 7364
rect 20993 7327 21051 7333
rect 20993 7293 21005 7327
rect 21039 7324 21051 7327
rect 22370 7324 22376 7336
rect 21039 7296 22376 7324
rect 21039 7293 21051 7296
rect 20993 7287 21051 7293
rect 22370 7284 22376 7296
rect 22428 7324 22434 7336
rect 22741 7327 22799 7333
rect 22741 7324 22753 7327
rect 22428 7296 22753 7324
rect 22428 7284 22434 7296
rect 22741 7293 22753 7296
rect 22787 7293 22799 7327
rect 22848 7324 22876 7364
rect 22925 7361 22937 7395
rect 22971 7361 22983 7395
rect 22925 7355 22983 7361
rect 23014 7352 23020 7404
rect 23072 7392 23078 7404
rect 23676 7401 23704 7432
rect 23768 7432 24133 7460
rect 23201 7395 23259 7401
rect 23201 7392 23213 7395
rect 23072 7364 23213 7392
rect 23072 7352 23078 7364
rect 23201 7361 23213 7364
rect 23247 7361 23259 7395
rect 23201 7355 23259 7361
rect 23385 7395 23443 7401
rect 23385 7361 23397 7395
rect 23431 7361 23443 7395
rect 23385 7355 23443 7361
rect 23661 7395 23719 7401
rect 23661 7361 23673 7395
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 23400 7324 23428 7355
rect 22848 7296 23428 7324
rect 22741 7287 22799 7293
rect 22278 7216 22284 7268
rect 22336 7256 22342 7268
rect 23109 7259 23167 7265
rect 23109 7256 23121 7259
rect 22336 7228 23121 7256
rect 22336 7216 22342 7228
rect 23109 7225 23121 7228
rect 23155 7256 23167 7259
rect 23768 7256 23796 7432
rect 24121 7429 24133 7432
rect 24167 7429 24179 7463
rect 24228 7460 24256 7488
rect 24397 7463 24455 7469
rect 24397 7460 24409 7463
rect 24228 7432 24409 7460
rect 24121 7423 24179 7429
rect 24397 7429 24409 7432
rect 24443 7429 24455 7463
rect 24397 7423 24455 7429
rect 23842 7352 23848 7404
rect 23900 7352 23906 7404
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7392 23995 7395
rect 23983 7364 24072 7392
rect 23983 7361 23995 7364
rect 23937 7355 23995 7361
rect 23155 7228 23796 7256
rect 23155 7225 23167 7228
rect 23109 7219 23167 7225
rect 18932 7160 20944 7188
rect 18932 7148 18938 7160
rect 21542 7148 21548 7200
rect 21600 7148 21606 7200
rect 23845 7191 23903 7197
rect 23845 7157 23857 7191
rect 23891 7188 23903 7191
rect 24044 7188 24072 7364
rect 24486 7352 24492 7404
rect 24544 7392 24550 7404
rect 24581 7395 24639 7401
rect 24581 7392 24593 7395
rect 24544 7364 24593 7392
rect 24544 7352 24550 7364
rect 24581 7361 24593 7364
rect 24627 7361 24639 7395
rect 24581 7355 24639 7361
rect 24765 7395 24823 7401
rect 24765 7361 24777 7395
rect 24811 7392 24823 7395
rect 25038 7392 25044 7404
rect 24811 7364 25044 7392
rect 24811 7361 24823 7364
rect 24765 7355 24823 7361
rect 25038 7352 25044 7364
rect 25096 7352 25102 7404
rect 25222 7352 25228 7404
rect 25280 7352 25286 7404
rect 24394 7188 24400 7200
rect 23891 7160 24400 7188
rect 23891 7157 23903 7160
rect 23845 7151 23903 7157
rect 24394 7148 24400 7160
rect 24452 7148 24458 7200
rect 24854 7148 24860 7200
rect 24912 7148 24918 7200
rect 24946 7148 24952 7200
rect 25004 7188 25010 7200
rect 25041 7191 25099 7197
rect 25041 7188 25053 7191
rect 25004 7160 25053 7188
rect 25004 7148 25010 7160
rect 25041 7157 25053 7160
rect 25087 7157 25099 7191
rect 25041 7151 25099 7157
rect 1104 7098 26496 7120
rect 1104 7046 4124 7098
rect 4176 7046 4188 7098
rect 4240 7046 4252 7098
rect 4304 7046 4316 7098
rect 4368 7046 4380 7098
rect 4432 7046 10472 7098
rect 10524 7046 10536 7098
rect 10588 7046 10600 7098
rect 10652 7046 10664 7098
rect 10716 7046 10728 7098
rect 10780 7046 16820 7098
rect 16872 7046 16884 7098
rect 16936 7046 16948 7098
rect 17000 7046 17012 7098
rect 17064 7046 17076 7098
rect 17128 7046 23168 7098
rect 23220 7046 23232 7098
rect 23284 7046 23296 7098
rect 23348 7046 23360 7098
rect 23412 7046 23424 7098
rect 23476 7046 26496 7098
rect 1104 7024 26496 7046
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 10492 6987 10550 6993
rect 4396 6956 5028 6984
rect 4396 6944 4402 6956
rect 3786 6876 3792 6928
rect 3844 6876 3850 6928
rect 4709 6919 4767 6925
rect 4709 6885 4721 6919
rect 4755 6885 4767 6919
rect 4709 6879 4767 6885
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3418 6848 3424 6860
rect 3283 6820 3424 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 4724 6848 4752 6879
rect 3568 6820 4752 6848
rect 3568 6808 3574 6820
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 4706 6789 4712 6792
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 3200 6752 4353 6780
rect 3200 6740 3206 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4544 6783 4602 6789
rect 4544 6782 4556 6783
rect 4341 6743 4399 6749
rect 4519 6749 4556 6782
rect 4590 6749 4602 6783
rect 4519 6743 4602 6749
rect 4676 6783 4712 6789
rect 4676 6749 4688 6783
rect 4676 6743 4712 6749
rect 3421 6715 3479 6721
rect 3421 6681 3433 6715
rect 3467 6681 3479 6715
rect 3421 6675 3479 6681
rect 3436 6644 3464 6675
rect 3602 6672 3608 6724
rect 3660 6712 3666 6724
rect 3878 6712 3884 6724
rect 3660 6684 3884 6712
rect 3660 6672 3666 6684
rect 3878 6672 3884 6684
rect 3936 6672 3942 6724
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 4519 6712 4547 6743
rect 4706 6740 4712 6743
rect 4764 6740 4770 6792
rect 5000 6789 5028 6956
rect 10492 6953 10504 6987
rect 10538 6984 10550 6987
rect 11146 6984 11152 6996
rect 10538 6956 11152 6984
rect 10538 6953 10550 6956
rect 10492 6947 10550 6953
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 11974 6944 11980 6996
rect 12032 6944 12038 6996
rect 16022 6944 16028 6996
rect 16080 6984 16086 6996
rect 16117 6987 16175 6993
rect 16117 6984 16129 6987
rect 16080 6956 16129 6984
rect 16080 6944 16086 6956
rect 16117 6953 16129 6956
rect 16163 6953 16175 6987
rect 16117 6947 16175 6953
rect 17586 6944 17592 6996
rect 17644 6984 17650 6996
rect 23293 6987 23351 6993
rect 17644 6956 22094 6984
rect 17644 6944 17650 6956
rect 8021 6919 8079 6925
rect 8021 6885 8033 6919
rect 8067 6885 8079 6919
rect 8021 6879 8079 6885
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 7926 6848 7932 6860
rect 5767 6820 7932 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8036 6848 8064 6879
rect 15194 6876 15200 6928
rect 15252 6916 15258 6928
rect 15657 6919 15715 6925
rect 15657 6916 15669 6919
rect 15252 6888 15669 6916
rect 15252 6876 15258 6888
rect 15657 6885 15669 6888
rect 15703 6916 15715 6919
rect 16390 6916 16396 6928
rect 15703 6888 16396 6916
rect 15703 6885 15715 6888
rect 15657 6879 15715 6885
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 22066 6916 22094 6956
rect 23293 6953 23305 6987
rect 23339 6984 23351 6987
rect 23566 6984 23572 6996
rect 23339 6956 23572 6984
rect 23339 6953 23351 6956
rect 23293 6947 23351 6953
rect 23566 6944 23572 6956
rect 23624 6984 23630 6996
rect 23753 6987 23811 6993
rect 23624 6956 23704 6984
rect 23624 6944 23630 6956
rect 23477 6919 23535 6925
rect 23477 6916 23489 6919
rect 22066 6888 23489 6916
rect 23477 6885 23489 6888
rect 23523 6885 23535 6919
rect 23676 6916 23704 6956
rect 23753 6953 23765 6987
rect 23799 6984 23811 6987
rect 23934 6984 23940 6996
rect 23799 6956 23940 6984
rect 23799 6953 23811 6956
rect 23753 6947 23811 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 24026 6944 24032 6996
rect 24084 6944 24090 6996
rect 25038 6944 25044 6996
rect 25096 6984 25102 6996
rect 26050 6984 26056 6996
rect 25096 6956 26056 6984
rect 25096 6944 25102 6956
rect 26050 6944 26056 6956
rect 26108 6984 26114 6996
rect 26145 6987 26203 6993
rect 26145 6984 26157 6987
rect 26108 6956 26157 6984
rect 26108 6944 26114 6956
rect 26145 6953 26157 6956
rect 26191 6953 26203 6987
rect 26145 6947 26203 6953
rect 23845 6919 23903 6925
rect 23845 6916 23857 6919
rect 23676 6888 23857 6916
rect 23477 6879 23535 6885
rect 23845 6885 23857 6888
rect 23891 6916 23903 6919
rect 24044 6916 24072 6944
rect 23891 6888 24072 6916
rect 23891 6885 23903 6888
rect 23845 6879 23903 6885
rect 8036 6820 9076 6848
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5353 6783 5411 6789
rect 5353 6780 5365 6783
rect 5031 6752 5365 6780
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 5353 6749 5365 6752
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 7883 6752 8156 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 5552 6712 5580 6743
rect 5994 6712 6000 6724
rect 4028 6684 6000 6712
rect 4028 6672 4034 6684
rect 5994 6672 6000 6684
rect 6052 6672 6058 6724
rect 4062 6644 4068 6656
rect 3436 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6644 4126 6656
rect 4338 6644 4344 6656
rect 4120 6616 4344 6644
rect 4120 6604 4126 6616
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 8128 6644 8156 6752
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 9048 6780 9076 6820
rect 9490 6808 9496 6860
rect 9548 6808 9554 6860
rect 10226 6808 10232 6860
rect 10284 6848 10290 6860
rect 11514 6848 11520 6860
rect 10284 6820 11520 6848
rect 10284 6808 10290 6820
rect 11514 6808 11520 6820
rect 11572 6848 11578 6860
rect 12069 6851 12127 6857
rect 12069 6848 12081 6851
rect 11572 6820 12081 6848
rect 11572 6808 11578 6820
rect 12069 6817 12081 6820
rect 12115 6848 12127 6851
rect 12434 6848 12440 6860
rect 12115 6820 12440 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 14182 6808 14188 6860
rect 14240 6848 14246 6860
rect 14642 6848 14648 6860
rect 14240 6820 14648 6848
rect 14240 6808 14246 6820
rect 14642 6808 14648 6820
rect 14700 6848 14706 6860
rect 14921 6851 14979 6857
rect 14921 6848 14933 6851
rect 14700 6820 14933 6848
rect 14700 6808 14706 6820
rect 14921 6817 14933 6820
rect 14967 6817 14979 6851
rect 19061 6851 19119 6857
rect 14921 6811 14979 6817
rect 15488 6820 16252 6848
rect 10042 6780 10048 6792
rect 9048 6752 10048 6780
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 15488 6780 15516 6820
rect 16224 6789 16252 6820
rect 19061 6817 19073 6851
rect 19107 6848 19119 6851
rect 19702 6848 19708 6860
rect 19107 6820 19708 6848
rect 19107 6817 19119 6820
rect 19061 6811 19119 6817
rect 19702 6808 19708 6820
rect 19760 6848 19766 6860
rect 19981 6851 20039 6857
rect 19981 6848 19993 6851
rect 19760 6820 19993 6848
rect 19760 6808 19766 6820
rect 19981 6817 19993 6820
rect 20027 6848 20039 6851
rect 20165 6851 20223 6857
rect 20165 6848 20177 6851
rect 20027 6820 20177 6848
rect 20027 6817 20039 6820
rect 19981 6811 20039 6817
rect 20165 6817 20177 6820
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 21545 6851 21603 6857
rect 21545 6817 21557 6851
rect 21591 6848 21603 6851
rect 22097 6851 22155 6857
rect 22097 6848 22109 6851
rect 21591 6820 22109 6848
rect 21591 6817 21603 6820
rect 21545 6811 21603 6817
rect 22097 6817 22109 6820
rect 22143 6817 22155 6851
rect 22097 6811 22155 6817
rect 23109 6851 23167 6857
rect 23109 6817 23121 6851
rect 23155 6848 23167 6851
rect 23937 6851 23995 6857
rect 23155 6820 23888 6848
rect 23155 6817 23167 6820
rect 23109 6811 23167 6817
rect 23860 6792 23888 6820
rect 23937 6817 23949 6851
rect 23983 6848 23995 6851
rect 24762 6848 24768 6860
rect 23983 6820 24768 6848
rect 23983 6817 23995 6820
rect 23937 6811 23995 6817
rect 24762 6808 24768 6820
rect 24820 6808 24826 6860
rect 14599 6752 15516 6780
rect 15565 6783 15623 6789
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 15565 6749 15577 6783
rect 15611 6780 15623 6783
rect 16025 6783 16083 6789
rect 16025 6780 16037 6783
rect 15611 6752 16037 6780
rect 15611 6749 15623 6752
rect 15565 6743 15623 6749
rect 16025 6749 16037 6752
rect 16071 6749 16083 6783
rect 16025 6743 16083 6749
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16574 6780 16580 6792
rect 16255 6752 16580 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 17310 6740 17316 6792
rect 17368 6740 17374 6792
rect 18690 6740 18696 6792
rect 18748 6740 18754 6792
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 21637 6783 21695 6789
rect 21637 6780 21649 6783
rect 19392 6752 21649 6780
rect 19392 6740 19398 6752
rect 21637 6749 21649 6752
rect 21683 6749 21695 6783
rect 21637 6743 21695 6749
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6749 21971 6783
rect 21913 6743 21971 6749
rect 23385 6783 23443 6789
rect 23385 6749 23397 6783
rect 23431 6780 23443 6783
rect 23474 6780 23480 6792
rect 23431 6752 23480 6780
rect 23431 6749 23443 6752
rect 23385 6743 23443 6749
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 9309 6715 9367 6721
rect 9309 6712 9321 6715
rect 8803 6684 9321 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 9309 6681 9321 6684
rect 9355 6681 9367 6715
rect 9309 6675 9367 6681
rect 9692 6684 10994 6712
rect 9692 6656 9720 6684
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8128 6616 8953 6644
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9088 6616 9413 6644
rect 9088 6604 9094 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 10888 6644 10916 6684
rect 12342 6672 12348 6724
rect 12400 6672 12406 6724
rect 12894 6672 12900 6724
rect 12952 6672 12958 6724
rect 15838 6672 15844 6724
rect 15896 6672 15902 6724
rect 17589 6715 17647 6721
rect 17589 6681 17601 6715
rect 17635 6712 17647 6715
rect 17678 6712 17684 6724
rect 17635 6684 17684 6712
rect 17635 6681 17647 6684
rect 17589 6675 17647 6681
rect 17678 6672 17684 6684
rect 17736 6672 17742 6724
rect 19794 6672 19800 6724
rect 19852 6712 19858 6724
rect 20901 6715 20959 6721
rect 20901 6712 20913 6715
rect 19852 6684 20913 6712
rect 19852 6672 19858 6684
rect 20901 6681 20913 6684
rect 20947 6681 20959 6715
rect 21928 6712 21956 6743
rect 23474 6740 23480 6752
rect 23532 6740 23538 6792
rect 23750 6740 23756 6792
rect 23808 6740 23814 6792
rect 23842 6740 23848 6792
rect 23900 6740 23906 6792
rect 24213 6783 24271 6789
rect 24213 6749 24225 6783
rect 24259 6780 24271 6783
rect 24302 6780 24308 6792
rect 24259 6752 24308 6780
rect 24259 6749 24271 6752
rect 24213 6743 24271 6749
rect 24302 6740 24308 6752
rect 24360 6740 24366 6792
rect 24397 6783 24455 6789
rect 24397 6749 24409 6783
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 20901 6675 20959 6681
rect 21652 6684 21956 6712
rect 23768 6712 23796 6740
rect 24412 6712 24440 6743
rect 23768 6684 24440 6712
rect 11790 6644 11796 6656
rect 10888 6616 11796 6644
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 13817 6647 13875 6653
rect 13817 6613 13829 6647
rect 13863 6644 13875 6647
rect 13998 6644 14004 6656
rect 13863 6616 14004 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 14458 6604 14464 6656
rect 14516 6604 14522 6656
rect 19426 6604 19432 6656
rect 19484 6604 19490 6656
rect 20809 6647 20867 6653
rect 20809 6613 20821 6647
rect 20855 6644 20867 6647
rect 21652 6644 21680 6684
rect 24670 6672 24676 6724
rect 24728 6672 24734 6724
rect 25682 6672 25688 6724
rect 25740 6672 25746 6724
rect 20855 6616 21680 6644
rect 20855 6613 20867 6616
rect 20809 6607 20867 6613
rect 21726 6604 21732 6656
rect 21784 6604 21790 6656
rect 22830 6604 22836 6656
rect 22888 6604 22894 6656
rect 23658 6604 23664 6656
rect 23716 6644 23722 6656
rect 24121 6647 24179 6653
rect 24121 6644 24133 6647
rect 23716 6616 24133 6644
rect 23716 6604 23722 6616
rect 24121 6613 24133 6616
rect 24167 6613 24179 6647
rect 24121 6607 24179 6613
rect 1104 6554 26656 6576
rect 1104 6502 7298 6554
rect 7350 6502 7362 6554
rect 7414 6502 7426 6554
rect 7478 6502 7490 6554
rect 7542 6502 7554 6554
rect 7606 6502 13646 6554
rect 13698 6502 13710 6554
rect 13762 6502 13774 6554
rect 13826 6502 13838 6554
rect 13890 6502 13902 6554
rect 13954 6502 19994 6554
rect 20046 6502 20058 6554
rect 20110 6502 20122 6554
rect 20174 6502 20186 6554
rect 20238 6502 20250 6554
rect 20302 6502 26342 6554
rect 26394 6502 26406 6554
rect 26458 6502 26470 6554
rect 26522 6502 26534 6554
rect 26586 6502 26598 6554
rect 26650 6502 26656 6554
rect 1104 6480 26656 6502
rect 3142 6400 3148 6452
rect 3200 6400 3206 6452
rect 3510 6400 3516 6452
rect 3568 6400 3574 6452
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 3786 6440 3792 6452
rect 3651 6412 3792 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 3936 6412 4169 6440
rect 3936 6400 3942 6412
rect 4157 6409 4169 6412
rect 4203 6409 4215 6443
rect 4157 6403 4215 6409
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 4798 6440 4804 6452
rect 4387 6412 4804 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 3528 6372 3556 6400
rect 3528 6344 3740 6372
rect 2774 6264 2780 6316
rect 2832 6264 2838 6316
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3602 6304 3608 6316
rect 3467 6276 3608 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3712 6313 3740 6344
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6273 3755 6307
rect 3988 6304 4016 6332
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3988 6276 4077 6304
rect 3697 6267 3755 6273
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4356 6304 4384 6403
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6409 5963 6443
rect 5905 6403 5963 6409
rect 4295 6276 4384 6304
rect 4479 6341 4537 6347
rect 4479 6307 4491 6341
rect 4525 6338 4537 6341
rect 4525 6307 4547 6338
rect 4614 6332 4620 6384
rect 4672 6332 4678 6384
rect 4709 6375 4767 6381
rect 4709 6341 4721 6375
rect 4755 6372 4767 6375
rect 4890 6372 4896 6384
rect 4755 6344 4896 6372
rect 4755 6341 4767 6344
rect 4709 6335 4767 6341
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 4982 6332 4988 6384
rect 5040 6332 5046 6384
rect 5920 6372 5948 6403
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 8110 6440 8116 6452
rect 6472 6412 8116 6440
rect 5920 6344 6224 6372
rect 4479 6301 4547 6307
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4519 6248 4547 6301
rect 4632 6304 4660 6332
rect 4801 6307 4859 6313
rect 4801 6304 4813 6307
rect 4632 6276 4813 6304
rect 1394 6196 1400 6248
rect 1452 6196 1458 6248
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 1719 6208 3249 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 4519 6236 4528 6248
rect 3237 6199 3295 6205
rect 3712 6208 4528 6236
rect 3712 6180 3740 6208
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 3694 6128 3700 6180
rect 3752 6128 3758 6180
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4632 6100 4660 6276
rect 4801 6273 4813 6276
rect 4847 6273 4859 6307
rect 4801 6267 4859 6273
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 5626 6304 5632 6316
rect 5491 6276 5632 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 6196 6313 6224 6344
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6227 6276 6377 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6236 5227 6239
rect 5534 6236 5540 6248
rect 5215 6208 5540 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 6012 6236 6040 6267
rect 6472 6236 6500 6412
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8260 6412 8861 6440
rect 8260 6400 8266 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 10689 6443 10747 6449
rect 10689 6409 10701 6443
rect 10735 6440 10747 6443
rect 10870 6440 10876 6452
rect 10735 6412 10876 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 11146 6400 11152 6452
rect 11204 6400 11210 6452
rect 11606 6400 11612 6452
rect 11664 6400 11670 6452
rect 11790 6400 11796 6452
rect 11848 6400 11854 6452
rect 13998 6400 14004 6452
rect 14056 6400 14062 6452
rect 14458 6400 14464 6452
rect 14516 6440 14522 6452
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14516 6412 14841 6440
rect 14516 6400 14522 6412
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 18874 6400 18880 6452
rect 18932 6400 18938 6452
rect 19334 6400 19340 6452
rect 19392 6400 19398 6452
rect 19610 6440 19616 6452
rect 19444 6412 19616 6440
rect 9674 6372 9680 6384
rect 8680 6344 9680 6372
rect 6012 6208 6500 6236
rect 4798 6128 4804 6180
rect 4856 6168 4862 6180
rect 5350 6168 5356 6180
rect 4856 6140 5356 6168
rect 4856 6128 4862 6140
rect 5350 6128 5356 6140
rect 5408 6168 5414 6180
rect 6012 6168 6040 6208
rect 7098 6196 7104 6248
rect 7156 6196 7162 6248
rect 7377 6239 7435 6245
rect 7377 6205 7389 6239
rect 7423 6236 7435 6239
rect 7926 6236 7932 6248
rect 7423 6208 7932 6236
rect 7423 6205 7435 6208
rect 7377 6199 7435 6205
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 8496 6236 8524 6290
rect 8680 6236 8708 6344
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 11624 6372 11652 6400
rect 11348 6344 11652 6372
rect 11808 6372 11836 6400
rect 11808 6344 12282 6372
rect 11348 6313 11376 6344
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 11514 6264 11520 6316
rect 11572 6264 11578 6316
rect 14016 6304 14044 6400
rect 19352 6313 19380 6400
rect 19444 6313 19472 6412
rect 19610 6400 19616 6412
rect 19668 6440 19674 6452
rect 20622 6440 20628 6452
rect 19668 6412 20628 6440
rect 19668 6400 19674 6412
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 21177 6443 21235 6449
rect 21177 6409 21189 6443
rect 21223 6409 21235 6443
rect 21177 6403 21235 6409
rect 19705 6375 19763 6381
rect 19705 6341 19717 6375
rect 19751 6372 19763 6375
rect 19794 6372 19800 6384
rect 19751 6344 19800 6372
rect 19751 6341 19763 6344
rect 19705 6335 19763 6341
rect 19794 6332 19800 6344
rect 19852 6332 19858 6384
rect 21192 6372 21220 6403
rect 21726 6400 21732 6452
rect 21784 6400 21790 6452
rect 21818 6400 21824 6452
rect 21876 6400 21882 6452
rect 22554 6400 22560 6452
rect 22612 6400 22618 6452
rect 22830 6400 22836 6452
rect 22888 6400 22894 6452
rect 23842 6400 23848 6452
rect 23900 6400 23906 6452
rect 24213 6443 24271 6449
rect 24213 6409 24225 6443
rect 24259 6440 24271 6443
rect 24670 6440 24676 6452
rect 24259 6412 24676 6440
rect 24259 6409 24271 6412
rect 24213 6403 24271 6409
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 21361 6375 21419 6381
rect 21361 6372 21373 6375
rect 21192 6344 21373 6372
rect 21361 6341 21373 6344
rect 21407 6372 21419 6375
rect 21744 6372 21772 6400
rect 21407 6344 21772 6372
rect 22848 6372 22876 6400
rect 22848 6344 23060 6372
rect 21407 6341 21419 6344
rect 21361 6335 21419 6341
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 14016 6276 14197 6304
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6273 19487 6307
rect 21174 6304 21180 6316
rect 20838 6276 21180 6304
rect 19429 6267 19487 6273
rect 21174 6264 21180 6276
rect 21232 6264 21238 6316
rect 21545 6307 21603 6313
rect 21545 6273 21557 6307
rect 21591 6273 21603 6307
rect 21545 6267 21603 6273
rect 21637 6307 21695 6313
rect 21637 6273 21649 6307
rect 21683 6304 21695 6307
rect 22186 6304 22192 6316
rect 21683 6276 22192 6304
rect 21683 6273 21695 6276
rect 21637 6267 21695 6273
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8496 6208 8708 6236
rect 8772 6208 8953 6236
rect 5408 6140 6040 6168
rect 5408 6128 5414 6140
rect 4571 6072 4660 6100
rect 5721 6103 5779 6109
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 5810 6100 5816 6112
rect 5767 6072 5816 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 5902 6060 5908 6112
rect 5960 6100 5966 6112
rect 6546 6100 6552 6112
rect 5960 6072 6552 6100
rect 5960 6060 5966 6072
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 7116 6100 7144 6196
rect 8588 6112 8616 6208
rect 8772 6112 8800 6208
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 9214 6196 9220 6248
rect 9272 6196 9278 6248
rect 11790 6196 11796 6248
rect 11848 6196 11854 6248
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13280 6208 13921 6236
rect 8110 6100 8116 6112
rect 7116 6072 8116 6100
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 10226 6100 10232 6112
rect 8812 6072 10232 6100
rect 8812 6060 8818 6072
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 13280 6109 13308 6208
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6236 16267 6239
rect 17402 6236 17408 6248
rect 16255 6208 17408 6236
rect 16255 6205 16267 6208
rect 16209 6199 16267 6205
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 19426 6128 19432 6180
rect 19484 6128 19490 6180
rect 13265 6103 13323 6109
rect 13265 6100 13277 6103
rect 12860 6072 13277 6100
rect 12860 6060 12866 6072
rect 13265 6069 13277 6072
rect 13311 6069 13323 6103
rect 13265 6063 13323 6069
rect 13354 6060 13360 6112
rect 13412 6060 13418 6112
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 15252 6072 15577 6100
rect 15252 6060 15258 6072
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 15565 6063 15623 6069
rect 19245 6103 19303 6109
rect 19245 6069 19257 6103
rect 19291 6100 19303 6103
rect 19444 6100 19472 6128
rect 19291 6072 19472 6100
rect 21560 6100 21588 6267
rect 22186 6264 22192 6276
rect 22244 6264 22250 6316
rect 22741 6307 22799 6313
rect 22741 6273 22753 6307
rect 22787 6273 22799 6307
rect 22741 6267 22799 6273
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 22373 6239 22431 6245
rect 22373 6236 22385 6239
rect 21784 6208 22385 6236
rect 21784 6196 21790 6208
rect 22373 6205 22385 6208
rect 22419 6205 22431 6239
rect 22373 6199 22431 6205
rect 21637 6171 21695 6177
rect 21637 6137 21649 6171
rect 21683 6168 21695 6171
rect 22756 6168 22784 6267
rect 22830 6264 22836 6316
rect 22888 6264 22894 6316
rect 23032 6313 23060 6344
rect 23017 6307 23075 6313
rect 23017 6273 23029 6307
rect 23063 6273 23075 6307
rect 23017 6267 23075 6273
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6273 23167 6307
rect 23109 6267 23167 6273
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6304 23535 6307
rect 23566 6304 23572 6316
rect 23523 6276 23572 6304
rect 23523 6273 23535 6276
rect 23477 6267 23535 6273
rect 22922 6236 22928 6248
rect 21683 6140 22784 6168
rect 22857 6208 22928 6236
rect 21683 6137 21695 6140
rect 21637 6131 21695 6137
rect 21726 6100 21732 6112
rect 21560 6072 21732 6100
rect 19291 6069 19303 6072
rect 19245 6063 19303 6069
rect 21726 6060 21732 6072
rect 21784 6060 21790 6112
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 22857 6100 22885 6208
rect 22922 6196 22928 6208
rect 22980 6196 22986 6248
rect 23124 6236 23152 6267
rect 23566 6264 23572 6276
rect 23624 6264 23630 6316
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6304 23811 6307
rect 23860 6304 23888 6400
rect 24302 6332 24308 6384
rect 24360 6332 24366 6384
rect 24578 6332 24584 6384
rect 24636 6332 24642 6384
rect 25501 6375 25559 6381
rect 25501 6372 25513 6375
rect 24780 6344 25513 6372
rect 23799 6276 23888 6304
rect 23799 6273 23811 6276
rect 23753 6267 23811 6273
rect 23032 6208 23152 6236
rect 24320 6236 24348 6332
rect 24394 6264 24400 6316
rect 24452 6264 24458 6316
rect 24486 6264 24492 6316
rect 24544 6264 24550 6316
rect 24780 6313 24808 6344
rect 25501 6341 25513 6344
rect 25547 6341 25559 6375
rect 25501 6335 25559 6341
rect 24765 6307 24823 6313
rect 24765 6273 24777 6307
rect 24811 6273 24823 6307
rect 24765 6267 24823 6273
rect 25225 6307 25283 6313
rect 25225 6273 25237 6307
rect 25271 6273 25283 6307
rect 25225 6267 25283 6273
rect 24857 6239 24915 6245
rect 24857 6236 24869 6239
rect 24320 6208 24869 6236
rect 23032 6180 23060 6208
rect 24857 6205 24869 6208
rect 24903 6205 24915 6239
rect 24857 6199 24915 6205
rect 25130 6196 25136 6248
rect 25188 6196 25194 6248
rect 23014 6128 23020 6180
rect 23072 6128 23078 6180
rect 25240 6168 25268 6267
rect 26050 6264 26056 6316
rect 26108 6264 26114 6316
rect 23492 6140 25268 6168
rect 23492 6112 23520 6140
rect 22612 6072 22885 6100
rect 22612 6060 22618 6072
rect 22922 6060 22928 6112
rect 22980 6100 22986 6112
rect 23201 6103 23259 6109
rect 23201 6100 23213 6103
rect 22980 6072 23213 6100
rect 22980 6060 22986 6072
rect 23201 6069 23213 6072
rect 23247 6069 23259 6103
rect 23201 6063 23259 6069
rect 23474 6060 23480 6112
rect 23532 6060 23538 6112
rect 1104 6010 26496 6032
rect 1104 5958 4124 6010
rect 4176 5958 4188 6010
rect 4240 5958 4252 6010
rect 4304 5958 4316 6010
rect 4368 5958 4380 6010
rect 4432 5958 10472 6010
rect 10524 5958 10536 6010
rect 10588 5958 10600 6010
rect 10652 5958 10664 6010
rect 10716 5958 10728 6010
rect 10780 5958 16820 6010
rect 16872 5958 16884 6010
rect 16936 5958 16948 6010
rect 17000 5958 17012 6010
rect 17064 5958 17076 6010
rect 17128 5958 23168 6010
rect 23220 5958 23232 6010
rect 23284 5958 23296 6010
rect 23348 5958 23360 6010
rect 23412 5958 23424 6010
rect 23476 5958 26496 6010
rect 1104 5936 26496 5958
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3200 5868 3433 5896
rect 3200 5856 3206 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 3421 5859 3479 5865
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3660 5868 3801 5896
rect 3660 5856 3666 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4430 5896 4436 5908
rect 4019 5868 4436 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4430 5856 4436 5868
rect 4488 5896 4494 5908
rect 4798 5896 4804 5908
rect 4488 5868 4804 5896
rect 4488 5856 4494 5868
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5445 5899 5503 5905
rect 5445 5896 5457 5899
rect 4948 5868 5457 5896
rect 4948 5856 4954 5868
rect 5445 5865 5457 5868
rect 5491 5865 5503 5899
rect 5445 5859 5503 5865
rect 5534 5856 5540 5908
rect 5592 5856 5598 5908
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5684 5868 5825 5896
rect 5684 5856 5690 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 5813 5859 5871 5865
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 8662 5896 8668 5908
rect 6604 5868 8668 5896
rect 6604 5856 6610 5868
rect 8662 5856 8668 5868
rect 8720 5896 8726 5908
rect 9030 5896 9036 5908
rect 8720 5868 9036 5896
rect 8720 5856 8726 5868
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9214 5856 9220 5908
rect 9272 5896 9278 5908
rect 9861 5899 9919 5905
rect 9861 5896 9873 5899
rect 9272 5868 9873 5896
rect 9272 5856 9278 5868
rect 9861 5865 9873 5868
rect 9907 5865 9919 5899
rect 9861 5859 9919 5865
rect 11609 5899 11667 5905
rect 11609 5865 11621 5899
rect 11655 5896 11667 5899
rect 11790 5896 11796 5908
rect 11655 5868 11796 5896
rect 11655 5865 11667 5868
rect 11609 5859 11667 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 13354 5896 13360 5908
rect 12406 5868 13360 5896
rect 3160 5701 3188 5856
rect 3344 5732 4200 5760
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3234 5584 3240 5636
rect 3292 5584 3298 5636
rect 3053 5559 3111 5565
rect 3053 5525 3065 5559
rect 3099 5556 3111 5559
rect 3344 5556 3372 5732
rect 3878 5652 3884 5704
rect 3936 5652 3942 5704
rect 4172 5692 4200 5732
rect 4798 5692 4804 5704
rect 4172 5664 4804 5692
rect 3453 5627 3511 5633
rect 3453 5593 3465 5627
rect 3499 5624 3511 5627
rect 3896 5624 3924 5652
rect 4172 5633 4200 5664
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5074 5652 5080 5704
rect 5132 5652 5138 5704
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5661 5503 5695
rect 5552 5692 5580 5856
rect 6089 5763 6147 5769
rect 6089 5729 6101 5763
rect 6135 5729 6147 5763
rect 6089 5723 6147 5729
rect 5629 5695 5687 5701
rect 5629 5692 5641 5695
rect 5552 5664 5641 5692
rect 5445 5655 5503 5661
rect 5629 5661 5641 5664
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 3499 5596 3924 5624
rect 4157 5627 4215 5633
rect 3499 5593 3511 5596
rect 3453 5587 3511 5593
rect 4157 5593 4169 5627
rect 4203 5593 4215 5627
rect 5460 5624 5488 5655
rect 6104 5624 6132 5723
rect 6914 5720 6920 5772
rect 6972 5720 6978 5772
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8168 5732 8401 5760
rect 8168 5720 8174 5732
rect 8389 5729 8401 5732
rect 8435 5729 8447 5763
rect 9048 5760 9076 5856
rect 9048 5732 9904 5760
rect 8389 5723 8447 5729
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 6932 5692 6960 5720
rect 6227 5664 6684 5692
rect 6932 5664 7038 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 4157 5587 4215 5593
rect 4264 5596 6132 5624
rect 3099 5528 3372 5556
rect 3099 5525 3111 5528
rect 3053 5519 3111 5525
rect 3602 5516 3608 5568
rect 3660 5516 3666 5568
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3947 5559 4005 5565
rect 3947 5556 3959 5559
rect 3752 5528 3959 5556
rect 3752 5516 3758 5528
rect 3947 5525 3959 5528
rect 3993 5525 4005 5559
rect 3947 5519 4005 5525
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4264 5556 4292 5596
rect 6454 5584 6460 5636
rect 6512 5584 6518 5636
rect 4120 5528 4292 5556
rect 5261 5559 5319 5565
rect 4120 5516 4126 5528
rect 5261 5525 5273 5559
rect 5307 5556 5319 5559
rect 6472 5556 6500 5584
rect 6656 5565 6684 5664
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9674 5652 9680 5704
rect 9732 5652 9738 5704
rect 9876 5701 9904 5732
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5692 9919 5695
rect 10318 5692 10324 5704
rect 9907 5664 10324 5692
rect 9907 5661 9919 5664
rect 9861 5655 9919 5661
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5692 11483 5695
rect 11885 5695 11943 5701
rect 11885 5692 11897 5695
rect 11471 5664 11897 5692
rect 11471 5661 11483 5664
rect 11425 5655 11483 5661
rect 11885 5661 11897 5664
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5692 12127 5695
rect 12406 5692 12434 5868
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 14090 5856 14096 5908
rect 14148 5856 14154 5908
rect 21726 5856 21732 5908
rect 21784 5856 21790 5908
rect 22738 5856 22744 5908
rect 22796 5856 22802 5908
rect 22830 5856 22836 5908
rect 22888 5856 22894 5908
rect 22922 5856 22928 5908
rect 22980 5856 22986 5908
rect 24949 5899 25007 5905
rect 24949 5865 24961 5899
rect 24995 5896 25007 5899
rect 25222 5896 25228 5908
rect 24995 5868 25228 5896
rect 24995 5865 25007 5868
rect 24949 5859 25007 5865
rect 25222 5856 25228 5868
rect 25280 5856 25286 5908
rect 12710 5788 12716 5840
rect 12768 5828 12774 5840
rect 13449 5831 13507 5837
rect 13449 5828 13461 5831
rect 12768 5800 13461 5828
rect 12768 5788 12774 5800
rect 13449 5797 13461 5800
rect 13495 5797 13507 5831
rect 13449 5791 13507 5797
rect 12115 5664 12434 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 13078 5652 13084 5704
rect 13136 5652 13142 5704
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5692 13691 5695
rect 14108 5692 14136 5856
rect 14642 5788 14648 5840
rect 14700 5788 14706 5840
rect 21361 5831 21419 5837
rect 21361 5797 21373 5831
rect 21407 5828 21419 5831
rect 21634 5828 21640 5840
rect 21407 5800 21640 5828
rect 21407 5797 21419 5800
rect 21361 5791 21419 5797
rect 16574 5720 16580 5772
rect 16632 5760 16638 5772
rect 16632 5732 17540 5760
rect 16632 5720 16638 5732
rect 17512 5704 17540 5732
rect 19610 5720 19616 5772
rect 19668 5720 19674 5772
rect 13679 5664 14136 5692
rect 14185 5695 14243 5701
rect 13679 5661 13691 5664
rect 13633 5655 13691 5661
rect 14185 5661 14197 5695
rect 14231 5661 14243 5695
rect 14185 5655 14243 5661
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5692 17279 5695
rect 17310 5692 17316 5704
rect 17267 5664 17316 5692
rect 17267 5661 17279 5664
rect 17221 5655 17279 5661
rect 8113 5627 8171 5633
rect 8113 5593 8125 5627
rect 8159 5624 8171 5627
rect 8941 5627 8999 5633
rect 8941 5624 8953 5627
rect 8159 5596 8953 5624
rect 8159 5593 8171 5596
rect 8113 5587 8171 5593
rect 8941 5593 8953 5596
rect 8987 5593 8999 5627
rect 8941 5587 8999 5593
rect 12253 5627 12311 5633
rect 12253 5593 12265 5627
rect 12299 5624 12311 5627
rect 12342 5624 12348 5636
rect 12299 5596 12348 5624
rect 12299 5593 12311 5596
rect 12253 5587 12311 5593
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 13096 5624 13124 5652
rect 14200 5624 14228 5655
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 17402 5652 17408 5704
rect 17460 5652 17466 5704
rect 17494 5652 17500 5704
rect 17552 5652 17558 5704
rect 21468 5701 21496 5800
rect 21634 5788 21640 5800
rect 21692 5788 21698 5840
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 13096 5596 15716 5624
rect 5307 5528 6500 5556
rect 6641 5559 6699 5565
rect 5307 5525 5319 5528
rect 5261 5519 5319 5525
rect 6641 5525 6653 5559
rect 6687 5556 6699 5559
rect 7098 5556 7104 5568
rect 6687 5528 7104 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 13170 5516 13176 5568
rect 13228 5556 13234 5568
rect 14369 5559 14427 5565
rect 14369 5556 14381 5559
rect 13228 5528 14381 5556
rect 13228 5516 13234 5528
rect 14369 5525 14381 5528
rect 14415 5556 14427 5559
rect 14458 5556 14464 5568
rect 14415 5528 14464 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 14458 5516 14464 5528
rect 14516 5556 14522 5568
rect 15286 5556 15292 5568
rect 14516 5528 15292 5556
rect 14516 5516 14522 5528
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 15473 5559 15531 5565
rect 15473 5525 15485 5559
rect 15519 5556 15531 5559
rect 15562 5556 15568 5568
rect 15519 5528 15568 5556
rect 15519 5525 15531 5528
rect 15473 5519 15531 5525
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 15688 5556 15716 5596
rect 16482 5584 16488 5636
rect 16540 5584 16546 5636
rect 16942 5584 16948 5636
rect 17000 5584 17006 5636
rect 19886 5584 19892 5636
rect 19944 5584 19950 5636
rect 21174 5624 21180 5636
rect 21114 5596 21180 5624
rect 21174 5584 21180 5596
rect 21232 5624 21238 5636
rect 21744 5624 21772 5856
rect 21913 5831 21971 5837
rect 21913 5797 21925 5831
rect 21959 5828 21971 5831
rect 22848 5828 22876 5856
rect 21959 5800 22876 5828
rect 21959 5797 21971 5800
rect 21913 5791 21971 5797
rect 22940 5760 22968 5856
rect 23109 5831 23167 5837
rect 23109 5797 23121 5831
rect 23155 5797 23167 5831
rect 23109 5791 23167 5797
rect 22756 5732 22968 5760
rect 22756 5701 22784 5732
rect 22741 5695 22799 5701
rect 22741 5661 22753 5695
rect 22787 5661 22799 5695
rect 22741 5655 22799 5661
rect 22925 5695 22983 5701
rect 22925 5661 22937 5695
rect 22971 5692 22983 5695
rect 23014 5692 23020 5704
rect 22971 5664 23020 5692
rect 22971 5661 22983 5664
rect 22925 5655 22983 5661
rect 22830 5624 22836 5636
rect 21232 5596 21404 5624
rect 21744 5596 22836 5624
rect 21232 5584 21238 5596
rect 17681 5559 17739 5565
rect 17681 5556 17693 5559
rect 15688 5528 17693 5556
rect 17681 5525 17693 5528
rect 17727 5556 17739 5559
rect 17862 5556 17868 5568
rect 17727 5528 17868 5556
rect 17727 5525 17739 5528
rect 17681 5519 17739 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 21376 5556 21404 5596
rect 22830 5584 22836 5596
rect 22888 5584 22894 5636
rect 22940 5624 22968 5655
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 23124 5692 23152 5791
rect 24765 5763 24823 5769
rect 24765 5729 24777 5763
rect 24811 5760 24823 5763
rect 24946 5760 24952 5772
rect 24811 5732 24952 5760
rect 24811 5729 24823 5732
rect 24765 5723 24823 5729
rect 24946 5720 24952 5732
rect 25004 5720 25010 5772
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 23124 5664 23213 5692
rect 23201 5661 23213 5664
rect 23247 5661 23259 5695
rect 23201 5655 23259 5661
rect 25038 5652 25044 5704
rect 25096 5652 25102 5704
rect 22940 5596 24532 5624
rect 21910 5556 21916 5568
rect 21376 5528 21916 5556
rect 21910 5516 21916 5528
rect 21968 5516 21974 5568
rect 22646 5516 22652 5568
rect 22704 5556 22710 5568
rect 23198 5556 23204 5568
rect 22704 5528 23204 5556
rect 22704 5516 22710 5528
rect 23198 5516 23204 5528
rect 23256 5556 23262 5568
rect 24504 5565 24532 5596
rect 23385 5559 23443 5565
rect 23385 5556 23397 5559
rect 23256 5528 23397 5556
rect 23256 5516 23262 5528
rect 23385 5525 23397 5528
rect 23431 5525 23443 5559
rect 23385 5519 23443 5525
rect 24489 5559 24547 5565
rect 24489 5525 24501 5559
rect 24535 5525 24547 5559
rect 24489 5519 24547 5525
rect 1104 5466 26656 5488
rect 1104 5414 7298 5466
rect 7350 5414 7362 5466
rect 7414 5414 7426 5466
rect 7478 5414 7490 5466
rect 7542 5414 7554 5466
rect 7606 5414 13646 5466
rect 13698 5414 13710 5466
rect 13762 5414 13774 5466
rect 13826 5414 13838 5466
rect 13890 5414 13902 5466
rect 13954 5414 19994 5466
rect 20046 5414 20058 5466
rect 20110 5414 20122 5466
rect 20174 5414 20186 5466
rect 20238 5414 20250 5466
rect 20302 5414 26342 5466
rect 26394 5414 26406 5466
rect 26458 5414 26470 5466
rect 26522 5414 26534 5466
rect 26586 5414 26598 5466
rect 26650 5414 26656 5466
rect 1104 5392 26656 5414
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5321 3203 5355
rect 3145 5315 3203 5321
rect 3160 5284 3188 5315
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 4341 5355 4399 5361
rect 4341 5352 4353 5355
rect 3568 5324 4353 5352
rect 3568 5312 3574 5324
rect 4341 5321 4353 5324
rect 4387 5321 4399 5355
rect 4341 5315 4399 5321
rect 4890 5312 4896 5364
rect 4948 5312 4954 5364
rect 5629 5355 5687 5361
rect 5629 5321 5641 5355
rect 5675 5352 5687 5355
rect 5718 5352 5724 5364
rect 5675 5324 5724 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 8297 5355 8355 5361
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 9490 5352 9496 5364
rect 8343 5324 9496 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 9674 5312 9680 5364
rect 9732 5312 9738 5364
rect 14921 5355 14979 5361
rect 14921 5321 14933 5355
rect 14967 5352 14979 5355
rect 15102 5352 15108 5364
rect 14967 5324 15108 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 16574 5352 16580 5364
rect 15488 5324 16580 5352
rect 3234 5284 3240 5296
rect 3160 5256 3240 5284
rect 3234 5244 3240 5256
rect 3292 5284 3298 5296
rect 3973 5287 4031 5293
rect 3973 5284 3985 5287
rect 3292 5256 3985 5284
rect 3292 5244 3298 5256
rect 3973 5253 3985 5256
rect 4019 5284 4031 5287
rect 4062 5284 4068 5296
rect 4019 5256 4068 5284
rect 4019 5253 4031 5256
rect 3973 5247 4031 5253
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 2806 5188 2912 5216
rect 2884 5160 2912 5188
rect 3602 5176 3608 5228
rect 3660 5176 3666 5228
rect 3694 5176 3700 5228
rect 3752 5176 3758 5228
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 4908 5216 4936 5312
rect 8386 5284 8392 5296
rect 8128 5256 8392 5284
rect 5077 5219 5135 5225
rect 5077 5216 5089 5219
rect 4908 5188 5089 5216
rect 4249 5179 4307 5185
rect 5077 5185 5089 5188
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 1719 5120 2774 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 2746 5080 2774 5120
rect 2866 5108 2872 5160
rect 2924 5108 2930 5160
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 3712 5148 3740 5176
rect 3559 5120 3740 5148
rect 3881 5151 3939 5157
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 3970 5148 3976 5160
rect 3927 5120 3976 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 2746 5052 3341 5080
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 4264 5080 4292 5179
rect 7098 5176 7104 5228
rect 7156 5176 7162 5228
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8128 5225 8156 5256
rect 8386 5244 8392 5256
rect 8444 5284 8450 5296
rect 9692 5284 9720 5312
rect 8444 5256 9720 5284
rect 8444 5244 8450 5256
rect 11974 5244 11980 5296
rect 12032 5284 12038 5296
rect 12345 5287 12403 5293
rect 12345 5284 12357 5287
rect 12032 5256 12357 5284
rect 12032 5244 12038 5256
rect 12345 5253 12357 5256
rect 12391 5253 12403 5287
rect 12345 5247 12403 5253
rect 12636 5256 13492 5284
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9674 5216 9680 5228
rect 8803 5188 9680 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 12636 5225 12664 5256
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 12621 5219 12679 5225
rect 12621 5185 12633 5219
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5216 12771 5219
rect 12802 5216 12808 5228
rect 12759 5188 12808 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 5166 5108 5172 5160
rect 5224 5148 5230 5160
rect 5353 5151 5411 5157
rect 5353 5148 5365 5151
rect 5224 5120 5365 5148
rect 5224 5108 5230 5120
rect 5353 5117 5365 5120
rect 5399 5117 5411 5151
rect 5353 5111 5411 5117
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5148 7803 5151
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 7791 5120 7849 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 7837 5117 7849 5120
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 3329 5043 3387 5049
rect 3896 5052 4292 5080
rect 3896 5024 3924 5052
rect 4706 5040 4712 5092
rect 4764 5080 4770 5092
rect 5920 5080 5948 5108
rect 4764 5052 5948 5080
rect 7944 5080 7972 5176
rect 12544 5148 12572 5179
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 13004 5157 13032 5256
rect 13464 5225 13492 5256
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5216 13507 5219
rect 13633 5219 13691 5225
rect 13495 5188 13584 5216
rect 13495 5185 13507 5188
rect 13449 5179 13507 5185
rect 12989 5151 13047 5157
rect 12544 5120 12664 5148
rect 8573 5083 8631 5089
rect 8573 5080 8585 5083
rect 7944 5052 8585 5080
rect 4764 5040 4770 5052
rect 8573 5049 8585 5052
rect 8619 5049 8631 5083
rect 12636 5080 12664 5120
rect 12989 5117 13001 5151
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 13372 5080 13400 5179
rect 13556 5092 13584 5188
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13446 5080 13452 5092
rect 12636 5052 13452 5080
rect 8573 5043 8631 5049
rect 13004 5024 13032 5052
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 13538 5040 13544 5092
rect 13596 5040 13602 5092
rect 13648 5080 13676 5179
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 14424 5188 15117 5216
rect 14424 5176 14430 5188
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 15212 5148 15240 5179
rect 15378 5176 15384 5228
rect 15436 5176 15442 5228
rect 15488 5225 15516 5324
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 16669 5355 16727 5361
rect 16669 5321 16681 5355
rect 16715 5352 16727 5355
rect 16942 5352 16948 5364
rect 16715 5324 16948 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 19886 5312 19892 5364
rect 19944 5352 19950 5364
rect 19981 5355 20039 5361
rect 19981 5352 19993 5355
rect 19944 5324 19993 5352
rect 19944 5312 19950 5324
rect 19981 5321 19993 5324
rect 20027 5321 20039 5355
rect 19981 5315 20039 5321
rect 21542 5312 21548 5364
rect 21600 5312 21606 5364
rect 22557 5355 22615 5361
rect 22557 5352 22569 5355
rect 22112 5324 22569 5352
rect 16390 5284 16396 5296
rect 15764 5256 16396 5284
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 15562 5176 15568 5228
rect 15620 5176 15626 5228
rect 15764 5225 15792 5256
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 16485 5287 16543 5293
rect 16485 5253 16497 5287
rect 16531 5284 16543 5287
rect 17037 5287 17095 5293
rect 17037 5284 17049 5287
rect 16531 5256 17049 5284
rect 16531 5253 16543 5256
rect 16485 5247 16543 5253
rect 17037 5253 17049 5256
rect 17083 5253 17095 5287
rect 17037 5247 17095 5253
rect 17586 5244 17592 5296
rect 17644 5244 17650 5296
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 15838 5176 15844 5228
rect 15896 5216 15902 5228
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 15896 5188 16865 5216
rect 15896 5176 15902 5188
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 17218 5216 17224 5228
rect 17175 5188 17224 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 18690 5176 18696 5228
rect 18748 5176 18754 5228
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5216 20223 5219
rect 21560 5216 21588 5312
rect 22112 5293 22140 5324
rect 22557 5321 22569 5324
rect 22603 5352 22615 5355
rect 22738 5352 22744 5364
rect 22603 5324 22744 5352
rect 22603 5321 22615 5324
rect 22557 5315 22615 5321
rect 22738 5312 22744 5324
rect 22796 5312 22802 5364
rect 23198 5312 23204 5364
rect 23256 5312 23262 5364
rect 23566 5312 23572 5364
rect 23624 5352 23630 5364
rect 24305 5355 24363 5361
rect 24305 5352 24317 5355
rect 23624 5324 24317 5352
rect 23624 5312 23630 5324
rect 24305 5321 24317 5324
rect 24351 5321 24363 5355
rect 25130 5352 25136 5364
rect 24305 5315 24363 5321
rect 24412 5324 25136 5352
rect 22097 5287 22155 5293
rect 22097 5253 22109 5287
rect 22143 5253 22155 5287
rect 22097 5247 22155 5253
rect 22189 5287 22247 5293
rect 22189 5253 22201 5287
rect 22235 5284 22247 5287
rect 22462 5284 22468 5296
rect 22235 5256 22468 5284
rect 22235 5253 22247 5256
rect 22189 5247 22247 5253
rect 22462 5244 22468 5256
rect 22520 5244 22526 5296
rect 22646 5244 22652 5296
rect 22704 5284 22710 5296
rect 22704 5256 23060 5284
rect 22704 5244 22710 5256
rect 20211 5188 21588 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 22002 5176 22008 5228
rect 22060 5176 22066 5228
rect 22278 5176 22284 5228
rect 22336 5225 22342 5228
rect 22336 5219 22365 5225
rect 22353 5185 22365 5219
rect 22336 5179 22365 5185
rect 22336 5176 22342 5179
rect 22738 5176 22744 5228
rect 22796 5176 22802 5228
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 23032 5225 23060 5256
rect 23216 5225 23244 5312
rect 24210 5244 24216 5296
rect 24268 5284 24274 5296
rect 24412 5284 24440 5324
rect 25130 5312 25136 5324
rect 25188 5352 25194 5364
rect 25406 5352 25412 5364
rect 25188 5324 25412 5352
rect 25188 5312 25194 5324
rect 25406 5312 25412 5324
rect 25464 5312 25470 5364
rect 24268 5256 24440 5284
rect 24489 5287 24547 5293
rect 24268 5244 24274 5256
rect 24489 5253 24501 5287
rect 24535 5284 24547 5287
rect 25222 5284 25228 5296
rect 24535 5256 25228 5284
rect 24535 5253 24547 5256
rect 24489 5247 24547 5253
rect 25222 5244 25228 5256
rect 25280 5244 25286 5296
rect 23017 5219 23075 5225
rect 23017 5185 23029 5219
rect 23063 5185 23075 5219
rect 23017 5179 23075 5185
rect 23201 5219 23259 5225
rect 23201 5185 23213 5219
rect 23247 5185 23259 5219
rect 23201 5179 23259 5185
rect 23658 5176 23664 5228
rect 23716 5216 23722 5228
rect 24121 5219 24179 5225
rect 24121 5216 24133 5219
rect 23716 5188 24133 5216
rect 23716 5176 23722 5188
rect 24121 5185 24133 5188
rect 24167 5185 24179 5219
rect 24121 5179 24179 5185
rect 15580 5148 15608 5176
rect 15933 5151 15991 5157
rect 15933 5148 15945 5151
rect 15212 5120 15945 5148
rect 15933 5117 15945 5120
rect 15979 5148 15991 5151
rect 16390 5148 16396 5160
rect 15979 5120 16396 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 17310 5108 17316 5160
rect 17368 5108 17374 5160
rect 18138 5148 18144 5160
rect 17420 5120 18144 5148
rect 14642 5080 14648 5092
rect 13648 5052 14648 5080
rect 3878 4972 3884 5024
rect 3936 4972 3942 5024
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 5169 5015 5227 5021
rect 5169 5012 5181 5015
rect 4856 4984 5181 5012
rect 4856 4972 4862 4984
rect 5169 4981 5181 4984
rect 5215 5012 5227 5015
rect 5534 5012 5540 5024
rect 5215 4984 5540 5012
rect 5215 4981 5227 4984
rect 5169 4975 5227 4981
rect 5534 4972 5540 4984
rect 5592 5012 5598 5024
rect 5902 5012 5908 5024
rect 5592 4984 5908 5012
rect 5592 4972 5598 4984
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 12618 4972 12624 5024
rect 12676 4972 12682 5024
rect 12986 4972 12992 5024
rect 13044 4972 13050 5024
rect 13262 4972 13268 5024
rect 13320 4972 13326 5024
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 13648 5012 13676 5052
rect 14642 5040 14648 5052
rect 14700 5040 14706 5092
rect 15102 5040 15108 5092
rect 15160 5080 15166 5092
rect 15286 5080 15292 5092
rect 15160 5052 15292 5080
rect 15160 5040 15166 5052
rect 15286 5040 15292 5052
rect 15344 5080 15350 5092
rect 17420 5080 17448 5120
rect 18138 5108 18144 5120
rect 18196 5108 18202 5160
rect 22186 5108 22192 5160
rect 22244 5148 22250 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22244 5120 22477 5148
rect 22244 5108 22250 5120
rect 22465 5117 22477 5120
rect 22511 5148 22523 5151
rect 22756 5148 22784 5176
rect 24228 5148 24256 5244
rect 22511 5120 24256 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 15344 5052 17448 5080
rect 15344 5040 15350 5052
rect 13412 4984 13676 5012
rect 13817 5015 13875 5021
rect 13412 4972 13418 4984
rect 13817 4981 13829 5015
rect 13863 5012 13875 5015
rect 14182 5012 14188 5024
rect 13863 4984 14188 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 15657 5015 15715 5021
rect 15657 4981 15669 5015
rect 15703 5012 15715 5015
rect 16114 5012 16120 5024
rect 15703 4984 16120 5012
rect 15703 4981 15715 4984
rect 15657 4975 15715 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 17678 4972 17684 5024
rect 17736 5012 17742 5024
rect 18230 5012 18236 5024
rect 17736 4984 18236 5012
rect 17736 4972 17742 4984
rect 18230 4972 18236 4984
rect 18288 5012 18294 5024
rect 19061 5015 19119 5021
rect 19061 5012 19073 5015
rect 18288 4984 19073 5012
rect 18288 4972 18294 4984
rect 19061 4981 19073 4984
rect 19107 5012 19119 5015
rect 19242 5012 19248 5024
rect 19107 4984 19248 5012
rect 19107 4981 19119 4984
rect 19061 4975 19119 4981
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 21266 4972 21272 5024
rect 21324 5012 21330 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 21324 4984 21833 5012
rect 21324 4972 21330 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 21821 4975 21879 4981
rect 23385 5015 23443 5021
rect 23385 4981 23397 5015
rect 23431 5012 23443 5015
rect 23842 5012 23848 5024
rect 23431 4984 23848 5012
rect 23431 4981 23443 4984
rect 23385 4975 23443 4981
rect 23842 4972 23848 4984
rect 23900 4972 23906 5024
rect 23934 4972 23940 5024
rect 23992 4972 23998 5024
rect 26145 5015 26203 5021
rect 26145 4981 26157 5015
rect 26191 5012 26203 5015
rect 26510 5012 26516 5024
rect 26191 4984 26516 5012
rect 26191 4981 26203 4984
rect 26145 4975 26203 4981
rect 26510 4972 26516 4984
rect 26568 4972 26574 5024
rect 1104 4922 26496 4944
rect 1104 4870 4124 4922
rect 4176 4870 4188 4922
rect 4240 4870 4252 4922
rect 4304 4870 4316 4922
rect 4368 4870 4380 4922
rect 4432 4870 10472 4922
rect 10524 4870 10536 4922
rect 10588 4870 10600 4922
rect 10652 4870 10664 4922
rect 10716 4870 10728 4922
rect 10780 4870 16820 4922
rect 16872 4870 16884 4922
rect 16936 4870 16948 4922
rect 17000 4870 17012 4922
rect 17064 4870 17076 4922
rect 17128 4870 23168 4922
rect 23220 4870 23232 4922
rect 23284 4870 23296 4922
rect 23348 4870 23360 4922
rect 23412 4870 23424 4922
rect 23476 4870 26496 4922
rect 1104 4848 26496 4870
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 3602 4808 3608 4820
rect 2823 4780 3608 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 3694 4768 3700 4820
rect 3752 4768 3758 4820
rect 4433 4811 4491 4817
rect 4433 4777 4445 4811
rect 4479 4808 4491 4811
rect 4798 4808 4804 4820
rect 4479 4780 4804 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 5074 4808 5080 4820
rect 4939 4780 5080 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 5629 4811 5687 4817
rect 5629 4777 5641 4811
rect 5675 4808 5687 4811
rect 5810 4808 5816 4820
rect 5675 4780 5816 4808
rect 5675 4777 5687 4780
rect 5629 4771 5687 4777
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 9674 4768 9680 4820
rect 9732 4768 9738 4820
rect 10042 4768 10048 4820
rect 10100 4768 10106 4820
rect 12618 4768 12624 4820
rect 12676 4768 12682 4820
rect 13262 4768 13268 4820
rect 13320 4768 13326 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 14366 4808 14372 4820
rect 13679 4780 14372 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 14737 4811 14795 4817
rect 14737 4777 14749 4811
rect 14783 4808 14795 4811
rect 15378 4808 15384 4820
rect 14783 4780 15384 4808
rect 14783 4777 14795 4780
rect 14737 4771 14795 4777
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 15657 4811 15715 4817
rect 15657 4777 15669 4811
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 3234 4740 3240 4752
rect 2792 4712 3240 4740
rect 2792 4672 2820 4712
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 3329 4743 3387 4749
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 3712 4740 3740 4768
rect 3375 4712 3740 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 4706 4700 4712 4752
rect 4764 4700 4770 4752
rect 4816 4740 4844 4768
rect 8202 4740 8208 4752
rect 4816 4712 5948 4740
rect 2608 4644 2820 4672
rect 2608 4613 2636 4644
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4573 2651 4607
rect 2593 4567 2651 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2792 4604 2820 4644
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 3050 4672 3056 4684
rect 2915 4644 3056 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 3050 4632 3056 4644
rect 3108 4672 3114 4684
rect 3786 4672 3792 4684
rect 3108 4644 3792 4672
rect 3108 4632 3114 4644
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 4724 4672 4752 4700
rect 3988 4644 4752 4672
rect 5000 4644 5764 4672
rect 3988 4613 4016 4644
rect 2961 4607 3019 4613
rect 2961 4604 2973 4607
rect 2792 4576 2973 4604
rect 2685 4567 2743 4573
rect 2961 4573 2973 4576
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4522 4604 4528 4616
rect 4203 4576 4528 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 2700 4536 2728 4567
rect 3160 4536 3188 4567
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 3878 4536 3884 4548
rect 2700 4508 3884 4536
rect 3878 4496 3884 4508
rect 3936 4536 3942 4548
rect 4617 4539 4675 4545
rect 3936 4508 4292 4536
rect 3936 4496 3942 4508
rect 4264 4477 4292 4508
rect 4617 4505 4629 4539
rect 4663 4536 4675 4539
rect 4706 4536 4712 4548
rect 4663 4508 4712 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 4706 4496 4712 4508
rect 4764 4536 4770 4548
rect 5000 4536 5028 4644
rect 5276 4613 5304 4644
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 4764 4508 5028 4536
rect 4764 4496 4770 4508
rect 4430 4477 4436 4480
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4437 4307 4471
rect 4249 4431 4307 4437
rect 4417 4471 4436 4477
rect 4417 4437 4429 4471
rect 4417 4431 4436 4437
rect 4430 4428 4436 4431
rect 4488 4428 4494 4480
rect 5092 4468 5120 4567
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 5166 4496 5172 4548
rect 5224 4496 5230 4548
rect 5399 4539 5457 4545
rect 5399 4505 5411 4539
rect 5445 4536 5457 4539
rect 5626 4536 5632 4548
rect 5445 4508 5632 4536
rect 5445 4505 5457 4508
rect 5399 4499 5457 4505
rect 5626 4496 5632 4508
rect 5684 4496 5690 4548
rect 5736 4536 5764 4644
rect 5920 4606 5948 4712
rect 7116 4712 8208 4740
rect 5994 4606 6000 4616
rect 5920 4578 6000 4606
rect 5994 4564 6000 4578
rect 6052 4564 6058 4616
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 7116 4604 7144 4712
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 7561 4675 7619 4681
rect 7561 4672 7573 4675
rect 7248 4644 7573 4672
rect 7248 4632 7254 4644
rect 7561 4641 7573 4644
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4672 7711 4675
rect 8386 4672 8392 4684
rect 7699 4644 8392 4672
rect 7699 4641 7711 4644
rect 7653 4635 7711 4641
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8662 4632 8668 4684
rect 8720 4632 8726 4684
rect 8864 4644 10088 4672
rect 8864 4616 8892 4644
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 7116 4576 7297 4604
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8481 4607 8539 4613
rect 8481 4604 8493 4607
rect 7883 4576 8493 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 8481 4573 8493 4576
rect 8527 4604 8539 4607
rect 8846 4604 8852 4616
rect 8527 4576 8852 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 5813 4539 5871 4545
rect 5813 4536 5825 4539
rect 5736 4508 5825 4536
rect 5813 4505 5825 4508
rect 5859 4536 5871 4539
rect 6656 4536 6684 4564
rect 5859 4508 6684 4536
rect 7193 4539 7251 4545
rect 5859 4505 5871 4508
rect 5813 4499 5871 4505
rect 7193 4505 7205 4539
rect 7239 4536 7251 4539
rect 7760 4536 7788 4567
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 8938 4564 8944 4616
rect 8996 4564 9002 4616
rect 10060 4613 10088 4644
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9048 4576 9873 4604
rect 7239 4508 7788 4536
rect 7239 4505 7251 4508
rect 7193 4499 7251 4505
rect 8202 4496 8208 4548
rect 8260 4536 8266 4548
rect 8389 4539 8447 4545
rect 8389 4536 8401 4539
rect 8260 4508 8401 4536
rect 8260 4496 8266 4508
rect 8389 4505 8401 4508
rect 8435 4536 8447 4539
rect 9048 4536 9076 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 12636 4604 12664 4768
rect 13170 4740 13176 4752
rect 12820 4712 13176 4740
rect 12820 4681 12848 4712
rect 13170 4700 13176 4712
rect 13228 4700 13234 4752
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4641 12863 4675
rect 12805 4635 12863 4641
rect 12986 4632 12992 4684
rect 13044 4632 13050 4684
rect 13280 4613 13308 4768
rect 13446 4700 13452 4752
rect 13504 4740 13510 4752
rect 15470 4740 15476 4752
rect 13504 4712 13952 4740
rect 13504 4700 13510 4712
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 12636 4576 13185 4604
rect 10045 4567 10103 4573
rect 13173 4573 13185 4576
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4573 13323 4607
rect 13265 4567 13323 4573
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 13924 4613 13952 4712
rect 14108 4712 15476 4740
rect 13725 4607 13783 4613
rect 13725 4604 13737 4607
rect 13596 4576 13737 4604
rect 13596 4564 13602 4576
rect 13725 4573 13737 4576
rect 13771 4573 13783 4607
rect 13725 4567 13783 4573
rect 13909 4607 13967 4613
rect 13909 4573 13921 4607
rect 13955 4604 13967 4607
rect 13998 4604 14004 4616
rect 13955 4576 14004 4604
rect 13955 4573 13967 4576
rect 13909 4567 13967 4573
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 14108 4613 14136 4712
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 15672 4672 15700 4771
rect 15746 4768 15752 4820
rect 15804 4768 15810 4820
rect 15838 4768 15844 4820
rect 15896 4768 15902 4820
rect 16114 4768 16120 4820
rect 16172 4808 16178 4820
rect 16758 4808 16764 4820
rect 16172 4780 16764 4808
rect 16172 4768 16178 4780
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 17218 4768 17224 4820
rect 17276 4768 17282 4820
rect 17405 4811 17463 4817
rect 17405 4777 17417 4811
rect 17451 4808 17463 4811
rect 17586 4808 17592 4820
rect 17451 4780 17592 4808
rect 17451 4777 17463 4780
rect 17405 4771 17463 4777
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 22002 4768 22008 4820
rect 22060 4808 22066 4820
rect 22833 4811 22891 4817
rect 22833 4808 22845 4811
rect 22060 4780 22845 4808
rect 22060 4768 22066 4780
rect 22833 4777 22845 4780
rect 22879 4777 22891 4811
rect 22833 4771 22891 4777
rect 23150 4780 23704 4808
rect 15764 4740 15792 4768
rect 16301 4743 16359 4749
rect 16301 4740 16313 4743
rect 15764 4712 16313 4740
rect 16301 4709 16313 4712
rect 16347 4709 16359 4743
rect 17236 4740 17264 4768
rect 17773 4743 17831 4749
rect 17773 4740 17785 4743
rect 17236 4712 17785 4740
rect 16301 4703 16359 4709
rect 17773 4709 17785 4712
rect 17819 4740 17831 4743
rect 17957 4743 18015 4749
rect 17957 4740 17969 4743
rect 17819 4712 17969 4740
rect 17819 4709 17831 4712
rect 17773 4703 17831 4709
rect 17957 4709 17969 4712
rect 18003 4709 18015 4743
rect 17957 4703 18015 4709
rect 16945 4675 17003 4681
rect 16945 4672 16957 4675
rect 14200 4644 14503 4672
rect 14093 4607 14151 4613
rect 14093 4573 14105 4607
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 8435 4508 9076 4536
rect 9585 4539 9643 4545
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 9585 4505 9597 4539
rect 9631 4536 9643 4539
rect 10318 4536 10324 4548
rect 9631 4508 10324 4536
rect 9631 4505 9643 4508
rect 9585 4499 9643 4505
rect 10318 4496 10324 4508
rect 10376 4496 10382 4548
rect 12713 4539 12771 4545
rect 12713 4505 12725 4539
rect 12759 4536 12771 4539
rect 12986 4536 12992 4548
rect 12759 4508 12992 4536
rect 12759 4505 12771 4508
rect 12713 4499 12771 4505
rect 12986 4496 12992 4508
rect 13044 4536 13050 4548
rect 13354 4536 13360 4548
rect 13044 4508 13360 4536
rect 13044 4496 13050 4508
rect 13354 4496 13360 4508
rect 13412 4496 13418 4548
rect 13464 4536 13492 4564
rect 14200 4536 14228 4644
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 14475 4613 14503 4644
rect 14660 4644 15240 4672
rect 15672 4644 16957 4672
rect 14660 4616 14688 4644
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 14475 4607 14539 4613
rect 14475 4576 14493 4607
rect 14369 4567 14427 4573
rect 14481 4573 14493 4576
rect 14527 4573 14539 4607
rect 14481 4567 14539 4573
rect 13464 4508 14228 4536
rect 14384 4536 14412 4567
rect 14642 4564 14648 4616
rect 14700 4564 14706 4616
rect 14918 4564 14924 4616
rect 14976 4604 14982 4616
rect 15212 4613 15240 4644
rect 16945 4641 16957 4644
rect 16991 4672 17003 4675
rect 17313 4675 17371 4681
rect 16991 4644 17264 4672
rect 16991 4641 17003 4644
rect 16945 4635 17003 4641
rect 15105 4607 15163 4613
rect 15105 4604 15117 4607
rect 14976 4576 15117 4604
rect 14976 4564 14982 4576
rect 15105 4573 15117 4576
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4604 15255 4607
rect 15286 4604 15292 4616
rect 15243 4576 15292 4604
rect 15243 4573 15255 4576
rect 15197 4567 15255 4573
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 15427 4576 15945 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 14734 4536 14740 4548
rect 14384 4508 14740 4536
rect 14734 4496 14740 4508
rect 14792 4496 14798 4548
rect 14829 4539 14887 4545
rect 14829 4505 14841 4539
rect 14875 4536 14887 4539
rect 14875 4508 15424 4536
rect 14875 4505 14887 4508
rect 14829 4499 14887 4505
rect 5534 4468 5540 4480
rect 5092 4440 5540 4468
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 5776 4440 6101 4468
rect 5776 4428 5782 4440
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 7377 4471 7435 4477
rect 7377 4437 7389 4471
rect 7423 4468 7435 4471
rect 7650 4468 7656 4480
rect 7423 4440 7656 4468
rect 7423 4437 7435 4440
rect 7377 4431 7435 4437
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 8294 4468 8300 4480
rect 8067 4440 8300 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 11790 4428 11796 4480
rect 11848 4468 11854 4480
rect 12345 4471 12403 4477
rect 12345 4468 12357 4471
rect 11848 4440 12357 4468
rect 11848 4428 11854 4440
rect 12345 4437 12357 4440
rect 12391 4437 12403 4471
rect 12345 4431 12403 4437
rect 13078 4428 13084 4480
rect 13136 4468 13142 4480
rect 13725 4471 13783 4477
rect 13725 4468 13737 4471
rect 13136 4440 13737 4468
rect 13136 4428 13142 4440
rect 13725 4437 13737 4440
rect 13771 4468 13783 4471
rect 13998 4468 14004 4480
rect 13771 4440 14004 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 14090 4428 14096 4480
rect 14148 4468 14154 4480
rect 15010 4468 15016 4480
rect 14148 4440 15016 4468
rect 14148 4428 14154 4440
rect 15010 4428 15016 4440
rect 15068 4428 15074 4480
rect 15396 4468 15424 4508
rect 15470 4496 15476 4548
rect 15528 4536 15534 4548
rect 15948 4536 15976 4567
rect 16022 4564 16028 4616
rect 16080 4564 16086 4616
rect 16390 4564 16396 4616
rect 16448 4564 16454 4616
rect 16482 4564 16488 4616
rect 16540 4604 16546 4616
rect 16853 4607 16911 4613
rect 16853 4604 16865 4607
rect 16540 4576 16865 4604
rect 16540 4564 16546 4576
rect 16853 4573 16865 4576
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 17037 4607 17095 4613
rect 17037 4573 17049 4607
rect 17083 4573 17095 4607
rect 17037 4567 17095 4573
rect 16114 4536 16120 4548
rect 15528 4508 15884 4536
rect 15948 4508 16120 4536
rect 15528 4496 15534 4508
rect 15856 4480 15884 4508
rect 16114 4496 16120 4508
rect 16172 4496 16178 4548
rect 16301 4539 16359 4545
rect 16301 4505 16313 4539
rect 16347 4536 16359 4539
rect 16666 4536 16672 4548
rect 16347 4508 16672 4536
rect 16347 4505 16359 4508
rect 16301 4499 16359 4505
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 15654 4468 15660 4480
rect 15712 4477 15718 4480
rect 15712 4471 15736 4477
rect 15396 4440 15660 4468
rect 15654 4428 15660 4440
rect 15724 4437 15736 4471
rect 15712 4431 15736 4437
rect 15712 4428 15718 4431
rect 15838 4428 15844 4480
rect 15896 4468 15902 4480
rect 16485 4471 16543 4477
rect 16485 4468 16497 4471
rect 15896 4440 16497 4468
rect 15896 4428 15902 4440
rect 16485 4437 16497 4440
rect 16531 4437 16543 4471
rect 16868 4468 16896 4567
rect 17052 4536 17080 4567
rect 17126 4564 17132 4616
rect 17184 4564 17190 4616
rect 17236 4604 17264 4644
rect 17313 4641 17325 4675
rect 17359 4672 17371 4675
rect 17865 4675 17923 4681
rect 17359 4644 17632 4672
rect 17359 4641 17371 4644
rect 17313 4635 17371 4641
rect 17402 4604 17408 4616
rect 17236 4576 17408 4604
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 17494 4564 17500 4616
rect 17552 4564 17558 4616
rect 17604 4613 17632 4644
rect 17865 4641 17877 4675
rect 17911 4672 17923 4675
rect 17911 4644 19012 4672
rect 17911 4641 17923 4644
rect 17865 4635 17923 4641
rect 18984 4616 19012 4644
rect 19352 4644 19564 4672
rect 19352 4616 19380 4644
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 18138 4564 18144 4616
rect 18196 4564 18202 4616
rect 18414 4564 18420 4616
rect 18472 4604 18478 4616
rect 18472 4576 18828 4604
rect 18472 4564 18478 4576
rect 17218 4536 17224 4548
rect 17052 4508 17224 4536
rect 17218 4496 17224 4508
rect 17276 4536 17282 4548
rect 17512 4536 17540 4564
rect 17276 4508 17540 4536
rect 18156 4536 18184 4564
rect 18156 4508 18460 4536
rect 17276 4496 17282 4508
rect 17586 4468 17592 4480
rect 16868 4440 17592 4468
rect 16485 4431 16543 4437
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18325 4471 18383 4477
rect 18325 4468 18337 4471
rect 17920 4440 18337 4468
rect 17920 4428 17926 4440
rect 18325 4437 18337 4440
rect 18371 4437 18383 4471
rect 18432 4468 18460 4508
rect 18506 4496 18512 4548
rect 18564 4496 18570 4548
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4505 18751 4539
rect 18800 4536 18828 4576
rect 18966 4564 18972 4616
rect 19024 4564 19030 4616
rect 19334 4564 19340 4616
rect 19392 4564 19398 4616
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 19536 4613 19564 4644
rect 20622 4632 20628 4684
rect 20680 4632 20686 4684
rect 22649 4675 22707 4681
rect 22649 4641 22661 4675
rect 22695 4672 22707 4675
rect 22695 4644 22968 4672
rect 22695 4641 22707 4644
rect 22649 4635 22707 4641
rect 22940 4616 22968 4644
rect 19521 4607 19579 4613
rect 19521 4573 19533 4607
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19794 4564 19800 4616
rect 19852 4564 19858 4616
rect 22738 4564 22744 4616
rect 22796 4606 22802 4616
rect 22796 4578 22839 4606
rect 22796 4564 22802 4578
rect 22922 4564 22928 4616
rect 22980 4604 22986 4616
rect 23150 4604 23178 4780
rect 23566 4700 23572 4752
rect 23624 4700 23630 4752
rect 23584 4672 23612 4700
rect 23492 4644 23612 4672
rect 22980 4576 23178 4604
rect 23293 4607 23351 4613
rect 22980 4564 22986 4576
rect 23293 4573 23305 4607
rect 23339 4598 23351 4607
rect 23492 4604 23520 4644
rect 23400 4598 23520 4604
rect 23339 4576 23520 4598
rect 23569 4607 23627 4613
rect 23339 4573 23428 4576
rect 23293 4570 23428 4573
rect 23569 4573 23581 4607
rect 23615 4604 23627 4607
rect 23676 4604 23704 4780
rect 25222 4632 25228 4684
rect 25280 4632 25286 4684
rect 23615 4576 23704 4604
rect 23615 4573 23627 4576
rect 23293 4567 23351 4570
rect 23569 4567 23627 4573
rect 19889 4539 19947 4545
rect 19889 4536 19901 4539
rect 18800 4508 19901 4536
rect 18693 4499 18751 4505
rect 19889 4505 19901 4508
rect 19935 4505 19947 4539
rect 19889 4499 19947 4505
rect 18708 4468 18736 4499
rect 20898 4496 20904 4548
rect 20956 4496 20962 4548
rect 21910 4496 21916 4548
rect 21968 4496 21974 4548
rect 23584 4536 23612 4567
rect 23934 4564 23940 4616
rect 23992 4604 23998 4616
rect 24486 4604 24492 4616
rect 23992 4576 24492 4604
rect 23992 4564 23998 4576
rect 24486 4564 24492 4576
rect 24544 4604 24550 4616
rect 25317 4607 25375 4613
rect 25317 4604 25329 4607
rect 24544 4576 25329 4604
rect 24544 4564 24550 4576
rect 25317 4573 25329 4576
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 23658 4536 23664 4548
rect 23584 4508 23664 4536
rect 23658 4496 23664 4508
rect 23716 4496 23722 4548
rect 24210 4496 24216 4548
rect 24268 4496 24274 4548
rect 18432 4440 18736 4468
rect 18325 4431 18383 4437
rect 18874 4428 18880 4480
rect 18932 4428 18938 4480
rect 18966 4428 18972 4480
rect 19024 4468 19030 4480
rect 19337 4471 19395 4477
rect 19337 4468 19349 4471
rect 19024 4440 19349 4468
rect 19024 4428 19030 4440
rect 19337 4437 19349 4440
rect 19383 4437 19395 4471
rect 19337 4431 19395 4437
rect 19610 4428 19616 4480
rect 19668 4428 19674 4480
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 22922 4468 22928 4480
rect 22336 4440 22928 4468
rect 22336 4428 22342 4440
rect 22922 4428 22928 4440
rect 22980 4428 22986 4480
rect 23014 4428 23020 4480
rect 23072 4468 23078 4480
rect 23109 4471 23167 4477
rect 23109 4468 23121 4471
rect 23072 4440 23121 4468
rect 23072 4428 23078 4440
rect 23109 4437 23121 4440
rect 23155 4437 23167 4471
rect 23109 4431 23167 4437
rect 23290 4428 23296 4480
rect 23348 4468 23354 4480
rect 23477 4471 23535 4477
rect 23477 4468 23489 4471
rect 23348 4440 23489 4468
rect 23348 4428 23354 4440
rect 23477 4437 23489 4440
rect 23523 4468 23535 4471
rect 24228 4468 24256 4496
rect 23523 4440 24256 4468
rect 23523 4437 23535 4440
rect 23477 4431 23535 4437
rect 24578 4428 24584 4480
rect 24636 4428 24642 4480
rect 24854 4428 24860 4480
rect 24912 4468 24918 4480
rect 25409 4471 25467 4477
rect 25409 4468 25421 4471
rect 24912 4440 25421 4468
rect 24912 4428 24918 4440
rect 25409 4437 25421 4440
rect 25455 4437 25467 4471
rect 25409 4431 25467 4437
rect 1104 4378 26656 4400
rect 1104 4326 7298 4378
rect 7350 4326 7362 4378
rect 7414 4326 7426 4378
rect 7478 4326 7490 4378
rect 7542 4326 7554 4378
rect 7606 4326 13646 4378
rect 13698 4326 13710 4378
rect 13762 4326 13774 4378
rect 13826 4326 13838 4378
rect 13890 4326 13902 4378
rect 13954 4326 19994 4378
rect 20046 4326 20058 4378
rect 20110 4326 20122 4378
rect 20174 4326 20186 4378
rect 20238 4326 20250 4378
rect 20302 4326 26342 4378
rect 26394 4326 26406 4378
rect 26458 4326 26470 4378
rect 26522 4326 26534 4378
rect 26586 4326 26598 4378
rect 26650 4326 26656 4378
rect 1104 4304 26656 4326
rect 3050 4224 3056 4276
rect 3108 4224 3114 4276
rect 5442 4264 5448 4276
rect 4014 4236 5448 4264
rect 4014 4208 4042 4236
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5721 4267 5779 4273
rect 5721 4264 5733 4267
rect 5592 4236 5733 4264
rect 5592 4224 5598 4236
rect 5721 4233 5733 4236
rect 5767 4233 5779 4267
rect 5721 4227 5779 4233
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6089 4267 6147 4273
rect 6089 4264 6101 4267
rect 6052 4236 6101 4264
rect 6052 4224 6058 4236
rect 6089 4233 6101 4236
rect 6135 4233 6147 4267
rect 6089 4227 6147 4233
rect 3970 4196 3976 4208
rect 4028 4205 4042 4208
rect 4028 4199 4057 4205
rect 3160 4168 3976 4196
rect 3160 4137 3188 4168
rect 3970 4156 3976 4168
rect 4045 4165 4057 4199
rect 4028 4159 4057 4165
rect 5261 4199 5319 4205
rect 5261 4165 5273 4199
rect 5307 4196 5319 4199
rect 5810 4196 5816 4208
rect 5307 4168 5816 4196
rect 5307 4165 5319 4168
rect 5261 4159 5319 4165
rect 4028 4156 4034 4159
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 6104 4196 6132 4227
rect 6362 4224 6368 4276
rect 6420 4224 6426 4276
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 7469 4267 7527 4273
rect 7469 4264 7481 4267
rect 7248 4236 7481 4264
rect 7248 4224 7254 4236
rect 7469 4233 7481 4236
rect 7515 4233 7527 4267
rect 7469 4227 7527 4233
rect 8297 4267 8355 4273
rect 8297 4233 8309 4267
rect 8343 4264 8355 4267
rect 8938 4264 8944 4276
rect 8343 4236 8944 4264
rect 8343 4233 8355 4236
rect 8297 4227 8355 4233
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10226 4264 10232 4276
rect 10100 4236 10232 4264
rect 10100 4224 10106 4236
rect 10226 4224 10232 4236
rect 10284 4264 10290 4276
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 10284 4236 10517 4264
rect 10284 4224 10290 4236
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 10505 4227 10563 4233
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 13596 4236 13676 4264
rect 13596 4224 13602 4236
rect 6104 4168 6408 4196
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3510 4088 3516 4140
rect 3568 4128 3574 4140
rect 3568 4118 3648 4128
rect 3698 4121 3756 4127
rect 3698 4118 3710 4121
rect 3568 4100 3710 4118
rect 3568 4088 3574 4100
rect 3620 4090 3710 4100
rect 3698 4087 3710 4090
rect 3744 4087 3756 4121
rect 3786 4088 3792 4140
rect 3844 4088 3850 4140
rect 3878 4088 3884 4140
rect 3936 4088 3942 4140
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 5350 4088 5356 4140
rect 5408 4088 5414 4140
rect 5442 4088 5448 4140
rect 5500 4137 5506 4140
rect 5500 4131 5529 4137
rect 5517 4097 5529 4131
rect 5500 4091 5529 4097
rect 5500 4088 5506 4091
rect 5902 4088 5908 4140
rect 5960 4088 5966 4140
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 6104 4100 6193 4128
rect 3698 4081 3756 4087
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4029 3295 4063
rect 3237 4023 3295 4029
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4203 4032 4261 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 5074 4060 5080 4072
rect 4847 4032 5080 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 3252 3992 3280 4023
rect 3326 3992 3332 4004
rect 3252 3964 3332 3992
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 2682 3884 2688 3936
rect 2740 3884 2746 3936
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 3513 3927 3571 3933
rect 3513 3924 3525 3927
rect 3292 3896 3525 3924
rect 3292 3884 3298 3896
rect 3513 3893 3525 3896
rect 3559 3893 3571 3927
rect 3513 3887 3571 3893
rect 4430 3884 4436 3936
rect 4488 3924 4494 3936
rect 4614 3924 4620 3936
rect 4488 3896 4620 3924
rect 4488 3884 4494 3896
rect 4614 3884 4620 3896
rect 4672 3924 4678 3936
rect 4816 3924 4844 4023
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 5718 4060 5724 4072
rect 5675 4032 5724 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 4672 3896 4844 3924
rect 4672 3884 4678 3896
rect 4982 3884 4988 3936
rect 5040 3884 5046 3936
rect 5092 3924 5120 4020
rect 6104 4004 6132 4100
rect 6181 4097 6193 4100
rect 6227 4097 6239 4131
rect 6181 4091 6239 4097
rect 6380 4069 6408 4168
rect 6638 4156 6644 4208
rect 6696 4156 6702 4208
rect 9769 4199 9827 4205
rect 9769 4165 9781 4199
rect 9815 4196 9827 4199
rect 9815 4168 10088 4196
rect 9815 4165 9827 4168
rect 9769 4159 9827 4165
rect 6640 4153 6698 4156
rect 6640 4119 6652 4153
rect 6686 4119 6698 4153
rect 6640 4113 6698 4119
rect 7650 4088 7656 4140
rect 7708 4088 7714 4140
rect 10060 4128 10088 4168
rect 13170 4156 13176 4208
rect 13228 4196 13234 4208
rect 13648 4196 13676 4236
rect 13924 4236 14503 4264
rect 13924 4208 13952 4236
rect 13228 4168 13676 4196
rect 13228 4156 13234 4168
rect 6365 4063 6423 4069
rect 6365 4029 6377 4063
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 6086 3952 6092 4004
rect 6144 3992 6150 4004
rect 6840 3992 6868 4023
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 8680 4060 8708 4114
rect 10060 4100 10272 4128
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 8628 4032 8708 4060
rect 8772 4032 10057 4060
rect 8628 4020 8634 4032
rect 6144 3964 6868 3992
rect 6144 3952 6150 3964
rect 8772 3936 8800 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10244 4060 10272 4100
rect 10318 4088 10324 4140
rect 10376 4088 10382 4140
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10468 4100 10609 4128
rect 10468 4088 10474 4100
rect 10597 4097 10609 4100
rect 10643 4128 10655 4131
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10643 4100 10701 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10689 4097 10701 4100
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 11440 4100 12190 4128
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 10244 4032 10793 4060
rect 10045 4023 10103 4029
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 10060 3992 10088 4023
rect 10060 3964 10364 3992
rect 10336 3936 10364 3964
rect 11440 3936 11468 4100
rect 11517 4063 11575 4069
rect 11517 4029 11529 4063
rect 11563 4060 11575 4063
rect 13170 4060 13176 4072
rect 11563 4032 13176 4060
rect 11563 4029 11575 4032
rect 11517 4023 11575 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13541 4063 13599 4069
rect 13311 4032 13492 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 5092 3896 6561 3924
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 7984 3896 8217 3924
rect 7984 3884 7990 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8205 3887 8263 3893
rect 8754 3884 8760 3936
rect 8812 3884 8818 3936
rect 10134 3884 10140 3936
rect 10192 3884 10198 3936
rect 10318 3884 10324 3936
rect 10376 3884 10382 3936
rect 11422 3884 11428 3936
rect 11480 3884 11486 3936
rect 13464 3924 13492 4032
rect 13541 4029 13553 4063
rect 13587 4029 13599 4063
rect 13648 4060 13676 4168
rect 13906 4156 13912 4208
rect 13964 4156 13970 4208
rect 13998 4156 14004 4208
rect 14056 4156 14062 4208
rect 14366 4205 14372 4208
rect 14343 4199 14372 4205
rect 14343 4165 14355 4199
rect 14343 4159 14372 4165
rect 14366 4156 14372 4159
rect 14424 4156 14430 4208
rect 14475 4205 14503 4236
rect 14568 4236 14780 4264
rect 14568 4205 14596 4236
rect 14461 4199 14519 4205
rect 14461 4165 14473 4199
rect 14507 4165 14519 4199
rect 14461 4159 14519 4165
rect 14553 4199 14611 4205
rect 14553 4165 14565 4199
rect 14599 4165 14611 4199
rect 14553 4159 14611 4165
rect 14016 4128 14044 4156
rect 14645 4131 14703 4137
rect 14016 4126 14504 4128
rect 14645 4126 14657 4131
rect 14016 4100 14657 4126
rect 14476 4098 14657 4100
rect 14645 4097 14657 4098
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 13648 4032 14197 4060
rect 13541 4023 13599 4029
rect 14185 4029 14197 4032
rect 14231 4060 14243 4063
rect 14366 4060 14372 4072
rect 14231 4032 14372 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 13556 3992 13584 4023
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14752 4060 14780 4236
rect 15654 4224 15660 4276
rect 15712 4224 15718 4276
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 17313 4267 17371 4273
rect 17313 4264 17325 4267
rect 16632 4236 17325 4264
rect 16632 4224 16638 4236
rect 17313 4233 17325 4236
rect 17359 4233 17371 4267
rect 18598 4264 18604 4276
rect 17313 4227 17371 4233
rect 18064 4236 18604 4264
rect 15010 4088 15016 4140
rect 15068 4128 15074 4140
rect 15672 4128 15700 4224
rect 17773 4199 17831 4205
rect 17773 4196 17785 4199
rect 16960 4168 17785 4196
rect 16301 4131 16359 4137
rect 16301 4128 16313 4131
rect 15068 4100 15608 4128
rect 15672 4100 16313 4128
rect 15068 4088 15074 4100
rect 14476 4032 14780 4060
rect 14829 4063 14887 4069
rect 14476 4004 14504 4032
rect 14829 4029 14841 4063
rect 14875 4060 14887 4063
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 14875 4032 15485 4060
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15580 4060 15608 4100
rect 16301 4097 16313 4100
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16666 4088 16672 4140
rect 16724 4088 16730 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 16960 4137 16988 4168
rect 17773 4165 17785 4168
rect 17819 4165 17831 4199
rect 17773 4159 17831 4165
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16816 4100 16865 4128
rect 16816 4088 16822 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15580 4032 15853 4060
rect 15473 4023 15531 4029
rect 15841 4029 15853 4032
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 15930 4020 15936 4072
rect 15988 4020 15994 4072
rect 16022 4020 16028 4072
rect 16080 4020 16086 4072
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 16960 4060 16988 4091
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 17460 4100 17509 4128
rect 17460 4088 17466 4100
rect 17497 4097 17509 4100
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 17586 4088 17592 4140
rect 17644 4088 17650 4140
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 18064 4137 18092 4236
rect 18598 4224 18604 4236
rect 18656 4224 18662 4276
rect 19242 4224 19248 4276
rect 19300 4264 19306 4276
rect 19705 4267 19763 4273
rect 19705 4264 19717 4267
rect 19300 4236 19717 4264
rect 19300 4224 19306 4236
rect 19705 4233 19717 4236
rect 19751 4233 19763 4267
rect 19705 4227 19763 4233
rect 19794 4224 19800 4276
rect 19852 4224 19858 4276
rect 22278 4224 22284 4276
rect 22336 4224 22342 4276
rect 23842 4264 23848 4276
rect 22848 4236 23848 4264
rect 19812 4196 19840 4224
rect 19889 4199 19947 4205
rect 19889 4196 19901 4199
rect 18156 4168 19901 4196
rect 18156 4140 18184 4168
rect 19889 4165 19901 4168
rect 19935 4165 19947 4199
rect 19889 4159 19947 4165
rect 22189 4199 22247 4205
rect 22189 4165 22201 4199
rect 22235 4196 22247 4199
rect 22848 4196 22876 4236
rect 23842 4224 23848 4236
rect 23900 4224 23906 4276
rect 25314 4224 25320 4276
rect 25372 4264 25378 4276
rect 25501 4267 25559 4273
rect 25501 4264 25513 4267
rect 25372 4236 25513 4264
rect 25372 4224 25378 4236
rect 25501 4233 25513 4236
rect 25547 4233 25559 4267
rect 25501 4227 25559 4233
rect 22925 4199 22983 4205
rect 22925 4196 22937 4199
rect 22235 4168 22937 4196
rect 22235 4165 22247 4168
rect 22189 4159 22247 4165
rect 22925 4165 22937 4168
rect 22971 4165 22983 4199
rect 22925 4159 22983 4165
rect 23014 4156 23020 4208
rect 23072 4156 23078 4208
rect 23290 4156 23296 4208
rect 23348 4196 23354 4208
rect 23477 4199 23535 4205
rect 23477 4196 23489 4199
rect 23348 4168 23489 4196
rect 23348 4156 23354 4168
rect 23477 4165 23489 4168
rect 23523 4165 23535 4199
rect 23477 4159 23535 4165
rect 23566 4156 23572 4208
rect 23624 4196 23630 4208
rect 24302 4196 24308 4208
rect 23624 4168 24308 4196
rect 23624 4156 23630 4168
rect 24302 4156 24308 4168
rect 24360 4156 24366 4208
rect 25682 4196 25688 4208
rect 25254 4168 25688 4196
rect 25682 4156 25688 4168
rect 25740 4156 25746 4208
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 17920 4100 18061 4128
rect 17920 4088 17926 4100
rect 18049 4097 18061 4100
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 18138 4088 18144 4140
rect 18196 4088 18202 4140
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4128 18383 4131
rect 19610 4128 19616 4140
rect 18371 4100 19616 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 19797 4131 19855 4137
rect 19797 4097 19809 4131
rect 19843 4097 19855 4131
rect 19797 4091 19855 4097
rect 16172 4032 16988 4060
rect 16172 4020 16178 4032
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 18156 4060 18184 4088
rect 17184 4032 18184 4060
rect 18233 4063 18291 4069
rect 17184 4020 17190 4032
rect 18233 4029 18245 4063
rect 18279 4060 18291 4063
rect 18966 4060 18972 4072
rect 18279 4032 18972 4060
rect 18279 4029 18291 4032
rect 18233 4023 18291 4029
rect 18966 4020 18972 4032
rect 19024 4020 19030 4072
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 19392 4032 19533 4060
rect 19392 4020 19398 4032
rect 19521 4029 19533 4032
rect 19567 4029 19579 4063
rect 19521 4023 19579 4029
rect 13814 3992 13820 4004
rect 13556 3964 13820 3992
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 14458 3952 14464 4004
rect 14516 3952 14522 4004
rect 14921 3995 14979 4001
rect 14921 3992 14933 3995
rect 14568 3964 14933 3992
rect 14568 3924 14596 3964
rect 14921 3961 14933 3964
rect 14967 3961 14979 3995
rect 14921 3955 14979 3961
rect 15286 3952 15292 4004
rect 15344 3992 15350 4004
rect 16040 3992 16068 4020
rect 15344 3964 16712 3992
rect 15344 3952 15350 3964
rect 13464 3896 14596 3924
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16684 3933 16712 3964
rect 17218 3952 17224 4004
rect 17276 3952 17282 4004
rect 18141 3995 18199 4001
rect 18141 3961 18153 3995
rect 18187 3992 18199 3995
rect 18414 3992 18420 4004
rect 18187 3964 18420 3992
rect 18187 3961 18199 3964
rect 18141 3955 18199 3961
rect 18414 3952 18420 3964
rect 18472 3952 18478 4004
rect 18598 3952 18604 4004
rect 18656 3992 18662 4004
rect 19812 3992 19840 4091
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 20349 4131 20407 4137
rect 20349 4128 20361 4131
rect 20036 4100 20361 4128
rect 20036 4088 20042 4100
rect 20349 4097 20361 4100
rect 20395 4097 20407 4131
rect 23135 4131 23193 4137
rect 23135 4128 23147 4131
rect 20349 4091 20407 4097
rect 22850 4121 22908 4127
rect 22850 4087 22862 4121
rect 22896 4118 22908 4121
rect 22896 4090 22968 4118
rect 22896 4087 22908 4090
rect 22850 4081 22908 4087
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22511 4032 22784 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 18656 3964 19840 3992
rect 18656 3952 18662 3964
rect 16393 3927 16451 3933
rect 16393 3924 16405 3927
rect 16172 3896 16405 3924
rect 16172 3884 16178 3896
rect 16393 3893 16405 3896
rect 16439 3893 16451 3927
rect 16393 3887 16451 3893
rect 16669 3927 16727 3933
rect 16669 3893 16681 3927
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 17129 3927 17187 3933
rect 17129 3893 17141 3927
rect 17175 3924 17187 3927
rect 17236 3924 17264 3952
rect 17175 3896 17264 3924
rect 17175 3893 17187 3896
rect 17129 3887 17187 3893
rect 17770 3884 17776 3936
rect 17828 3884 17834 3936
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 18506 3924 18512 3936
rect 18012 3896 18512 3924
rect 18012 3884 18018 3896
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 18782 3884 18788 3936
rect 18840 3884 18846 3936
rect 20070 3884 20076 3936
rect 20128 3884 20134 3936
rect 20165 3927 20223 3933
rect 20165 3893 20177 3927
rect 20211 3924 20223 3927
rect 20346 3924 20352 3936
rect 20211 3896 20352 3924
rect 20211 3893 20223 3896
rect 20165 3887 20223 3893
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 21818 3884 21824 3936
rect 21876 3884 21882 3936
rect 22646 3884 22652 3936
rect 22704 3884 22710 3936
rect 22756 3924 22784 4032
rect 22940 3992 22968 4090
rect 23032 4100 23147 4128
rect 23032 4072 23060 4100
rect 23135 4097 23147 4100
rect 23181 4097 23193 4131
rect 23135 4091 23193 4097
rect 23382 4088 23388 4140
rect 23440 4088 23446 4140
rect 23658 4088 23664 4140
rect 23716 4088 23722 4140
rect 23750 4088 23756 4140
rect 23808 4088 23814 4140
rect 23014 4020 23020 4072
rect 23072 4020 23078 4072
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4060 23351 4063
rect 23566 4060 23572 4072
rect 23339 4032 23572 4060
rect 23339 4029 23351 4032
rect 23293 4023 23351 4029
rect 23566 4020 23572 4032
rect 23624 4020 23630 4072
rect 23385 3995 23443 4001
rect 23385 3992 23397 3995
rect 22940 3964 23397 3992
rect 23385 3961 23397 3964
rect 23431 3961 23443 3995
rect 23385 3955 23443 3961
rect 23676 3924 23704 4088
rect 24026 4020 24032 4072
rect 24084 4020 24090 4072
rect 25222 3924 25228 3936
rect 22756 3896 25228 3924
rect 25222 3884 25228 3896
rect 25280 3884 25286 3936
rect 1104 3834 26496 3856
rect 1104 3782 4124 3834
rect 4176 3782 4188 3834
rect 4240 3782 4252 3834
rect 4304 3782 4316 3834
rect 4368 3782 4380 3834
rect 4432 3782 10472 3834
rect 10524 3782 10536 3834
rect 10588 3782 10600 3834
rect 10652 3782 10664 3834
rect 10716 3782 10728 3834
rect 10780 3782 16820 3834
rect 16872 3782 16884 3834
rect 16936 3782 16948 3834
rect 17000 3782 17012 3834
rect 17064 3782 17076 3834
rect 17128 3782 23168 3834
rect 23220 3782 23232 3834
rect 23284 3782 23296 3834
rect 23348 3782 23360 3834
rect 23412 3782 23424 3834
rect 23476 3782 26496 3834
rect 1104 3760 26496 3782
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 3326 3720 3332 3732
rect 3283 3692 3332 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 3786 3680 3792 3732
rect 3844 3720 3850 3732
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 3844 3692 4169 3720
rect 3844 3680 3850 3692
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 4798 3720 4804 3732
rect 4157 3683 4215 3689
rect 4632 3692 4804 3720
rect 3344 3584 3372 3680
rect 4632 3584 4660 3692
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 4982 3729 4988 3732
rect 4972 3723 4988 3729
rect 4972 3689 4984 3723
rect 4972 3683 4988 3689
rect 4982 3680 4988 3683
rect 5040 3680 5046 3732
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 6362 3720 6368 3732
rect 5684 3692 6368 3720
rect 5684 3680 5690 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 6457 3723 6515 3729
rect 6457 3689 6469 3723
rect 6503 3720 6515 3723
rect 6638 3720 6644 3732
rect 6503 3692 6644 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 8757 3723 8815 3729
rect 8757 3689 8769 3723
rect 8803 3720 8815 3723
rect 8846 3720 8852 3732
rect 8803 3692 8852 3720
rect 8803 3689 8815 3692
rect 8757 3683 8815 3689
rect 8846 3680 8852 3692
rect 8904 3680 8910 3732
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 15930 3720 15936 3732
rect 14976 3692 15936 3720
rect 14976 3680 14982 3692
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 16264 3692 16313 3720
rect 16264 3680 16270 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16301 3683 16359 3689
rect 7006 3584 7012 3596
rect 3344 3556 4660 3584
rect 4632 3528 4660 3556
rect 4724 3556 7012 3584
rect 1394 3476 1400 3528
rect 1452 3516 1458 3528
rect 1489 3519 1547 3525
rect 1489 3516 1501 3519
rect 1452 3488 1501 3516
rect 1452 3476 1458 3488
rect 1489 3485 1501 3488
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 1504 3380 1532 3479
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4062 3516 4068 3528
rect 2924 3488 4068 3516
rect 2924 3476 2930 3488
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4522 3516 4528 3528
rect 4387 3488 4528 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 4614 3476 4620 3528
rect 4672 3476 4678 3528
rect 4724 3525 4752 3556
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 8864 3584 8892 3680
rect 13909 3655 13967 3661
rect 11992 3624 13860 3652
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8864 3556 9137 3584
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 10318 3544 10324 3596
rect 10376 3584 10382 3596
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 10376 3556 10701 3584
rect 10376 3544 10382 3556
rect 10689 3553 10701 3556
rect 10735 3584 10747 3587
rect 11514 3584 11520 3596
rect 10735 3556 11520 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 11514 3544 11520 3556
rect 11572 3584 11578 3596
rect 11992 3584 12020 3624
rect 13832 3596 13860 3624
rect 13909 3621 13921 3655
rect 13955 3652 13967 3655
rect 14274 3652 14280 3664
rect 13955 3624 14280 3652
rect 13955 3621 13967 3624
rect 13909 3615 13967 3621
rect 14274 3612 14280 3624
rect 14332 3612 14338 3664
rect 11572 3556 12020 3584
rect 12713 3587 12771 3593
rect 11572 3544 11578 3556
rect 12713 3553 12725 3587
rect 12759 3584 12771 3587
rect 12759 3556 13400 3584
rect 12759 3553 12771 3556
rect 12713 3547 12771 3553
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 9140 3488 10180 3516
rect 1762 3408 1768 3460
rect 1820 3408 1826 3460
rect 4724 3448 4752 3479
rect 6914 3448 6920 3460
rect 3160 3420 4752 3448
rect 6210 3420 6920 3448
rect 2774 3380 2780 3392
rect 1504 3352 2780 3380
rect 2774 3340 2780 3352
rect 2832 3380 2838 3392
rect 3160 3380 3188 3420
rect 6288 3392 6316 3420
rect 6914 3408 6920 3420
rect 6972 3408 6978 3460
rect 7285 3451 7343 3457
rect 7285 3417 7297 3451
rect 7331 3417 7343 3451
rect 8570 3448 8576 3460
rect 8510 3420 8576 3448
rect 7285 3411 7343 3417
rect 2832 3352 3188 3380
rect 4525 3383 4583 3389
rect 2832 3340 2838 3352
rect 4525 3349 4537 3383
rect 4571 3380 4583 3383
rect 4706 3380 4712 3392
rect 4571 3352 4712 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 6270 3340 6276 3392
rect 6328 3340 6334 3392
rect 7300 3380 7328 3411
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 8202 3380 8208 3392
rect 7300 3352 8208 3380
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 8588 3380 8616 3408
rect 9140 3380 9168 3488
rect 9214 3408 9220 3460
rect 9272 3448 9278 3460
rect 9861 3451 9919 3457
rect 9861 3448 9873 3451
rect 9272 3420 9873 3448
rect 9272 3408 9278 3420
rect 9861 3417 9873 3420
rect 9907 3417 9919 3451
rect 9861 3411 9919 3417
rect 9490 3380 9496 3392
rect 8588 3352 9496 3380
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 9766 3340 9772 3392
rect 9824 3340 9830 3392
rect 10152 3380 10180 3488
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10284 3488 10425 3516
rect 10284 3476 10290 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 13078 3476 13084 3528
rect 13136 3516 13142 3528
rect 13173 3519 13231 3525
rect 13173 3516 13185 3519
rect 13136 3488 13185 3516
rect 13136 3476 13142 3488
rect 13173 3485 13185 3488
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 13262 3476 13268 3528
rect 13320 3476 13326 3528
rect 13372 3516 13400 3556
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 13872 3556 14565 3584
rect 13872 3544 13878 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 14826 3544 14832 3596
rect 14884 3584 14890 3596
rect 16316 3584 16344 3683
rect 17770 3680 17776 3732
rect 17828 3720 17834 3732
rect 17828 3692 19012 3720
rect 17828 3680 17834 3692
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 14884 3556 16252 3584
rect 16316 3556 16957 3584
rect 14884 3544 14890 3556
rect 16224 3516 16252 3556
rect 16945 3553 16957 3556
rect 16991 3553 17003 3587
rect 16945 3547 17003 3553
rect 17310 3544 17316 3596
rect 17368 3544 17374 3596
rect 18874 3544 18880 3596
rect 18932 3544 18938 3596
rect 18984 3584 19012 3692
rect 19978 3680 19984 3732
rect 20036 3680 20042 3732
rect 20070 3680 20076 3732
rect 20128 3680 20134 3732
rect 22738 3680 22744 3732
rect 22796 3680 22802 3732
rect 23566 3680 23572 3732
rect 23624 3680 23630 3732
rect 24026 3680 24032 3732
rect 24084 3720 24090 3732
rect 24213 3723 24271 3729
rect 24213 3720 24225 3723
rect 24084 3692 24225 3720
rect 24084 3680 24090 3692
rect 24213 3689 24225 3692
rect 24259 3689 24271 3723
rect 24213 3683 24271 3689
rect 24302 3680 24308 3732
rect 24360 3720 24366 3732
rect 24360 3692 24992 3720
rect 24360 3680 24366 3692
rect 19337 3587 19395 3593
rect 19337 3584 19349 3587
rect 18984 3556 19349 3584
rect 19337 3553 19349 3556
rect 19383 3553 19395 3587
rect 19337 3547 19395 3553
rect 17126 3516 17132 3528
rect 13372 3488 14136 3516
rect 16224 3488 17132 3516
rect 10962 3408 10968 3460
rect 11020 3408 11026 3460
rect 11422 3448 11428 3460
rect 11072 3420 11428 3448
rect 11072 3380 11100 3420
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 12989 3451 13047 3457
rect 12989 3417 13001 3451
rect 13035 3417 13047 3451
rect 13280 3448 13308 3476
rect 14108 3460 14136 3488
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 18690 3476 18696 3528
rect 18748 3476 18754 3528
rect 18892 3516 18920 3544
rect 19150 3516 19156 3528
rect 18892 3488 19156 3516
rect 19150 3476 19156 3488
rect 19208 3516 19214 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19208 3488 19533 3516
rect 19208 3476 19214 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 20088 3516 20116 3680
rect 20622 3544 20628 3596
rect 20680 3544 20686 3596
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3584 20959 3587
rect 21266 3584 21272 3596
rect 20947 3556 21272 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 21910 3544 21916 3596
rect 21968 3584 21974 3596
rect 22649 3587 22707 3593
rect 21968 3556 22140 3584
rect 21968 3544 21974 3556
rect 19659 3488 20116 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 13998 3448 14004 3460
rect 13280 3420 14004 3448
rect 12989 3411 13047 3417
rect 10152 3352 11100 3380
rect 12802 3340 12808 3392
rect 12860 3340 12866 3392
rect 13004 3380 13032 3411
rect 13998 3408 14004 3420
rect 14056 3408 14062 3460
rect 14090 3408 14096 3460
rect 14148 3408 14154 3460
rect 14277 3451 14335 3457
rect 14277 3417 14289 3451
rect 14323 3448 14335 3451
rect 14366 3448 14372 3460
rect 14323 3420 14372 3448
rect 14323 3417 14335 3420
rect 14277 3411 14335 3417
rect 14366 3408 14372 3420
rect 14424 3448 14430 3460
rect 14424 3420 14596 3448
rect 14424 3408 14430 3420
rect 13446 3380 13452 3392
rect 13004 3352 13452 3380
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 14458 3340 14464 3392
rect 14516 3340 14522 3392
rect 14568 3380 14596 3420
rect 14826 3408 14832 3460
rect 14884 3408 14890 3460
rect 14918 3408 14924 3460
rect 14976 3408 14982 3460
rect 16298 3448 16304 3460
rect 16054 3420 16304 3448
rect 16298 3408 16304 3420
rect 16356 3408 16362 3460
rect 17586 3408 17592 3460
rect 17644 3408 17650 3460
rect 22112 3448 22140 3556
rect 22649 3553 22661 3587
rect 22695 3584 22707 3587
rect 22756 3584 22784 3680
rect 23584 3652 23612 3680
rect 24397 3655 24455 3661
rect 24397 3652 24409 3655
rect 23584 3624 24409 3652
rect 24397 3621 24409 3624
rect 24443 3621 24455 3655
rect 24397 3615 24455 3621
rect 22695 3556 22784 3584
rect 23569 3587 23627 3593
rect 22695 3553 22707 3556
rect 22649 3547 22707 3553
rect 23569 3553 23581 3587
rect 23615 3584 23627 3587
rect 24578 3584 24584 3596
rect 23615 3556 24584 3584
rect 23615 3553 23627 3556
rect 23569 3547 23627 3553
rect 24578 3544 24584 3556
rect 24636 3544 24642 3596
rect 24964 3593 24992 3692
rect 25314 3680 25320 3732
rect 25372 3680 25378 3732
rect 24949 3587 25007 3593
rect 24949 3553 24961 3587
rect 24995 3553 25007 3587
rect 25332 3584 25360 3680
rect 25593 3587 25651 3593
rect 25593 3584 25605 3587
rect 25332 3556 25605 3584
rect 24949 3547 25007 3553
rect 25593 3553 25605 3556
rect 25639 3553 25651 3587
rect 25593 3547 25651 3553
rect 23014 3476 23020 3528
rect 23072 3516 23078 3528
rect 23707 3519 23765 3525
rect 23707 3516 23719 3519
rect 23072 3488 23719 3516
rect 23072 3476 23078 3488
rect 23707 3485 23719 3488
rect 23753 3485 23765 3519
rect 23707 3479 23765 3485
rect 23842 3476 23848 3528
rect 23900 3476 23906 3528
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3516 24087 3519
rect 24854 3516 24860 3528
rect 24075 3488 24860 3516
rect 24075 3485 24087 3488
rect 24029 3479 24087 3485
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 24964 3516 24992 3547
rect 24964 3488 25268 3516
rect 23937 3451 23995 3457
rect 22112 3434 23796 3448
rect 22126 3420 23796 3434
rect 14936 3380 14964 3408
rect 23768 3392 23796 3420
rect 23937 3417 23949 3451
rect 23983 3448 23995 3451
rect 25240 3448 25268 3488
rect 25314 3476 25320 3528
rect 25372 3476 25378 3528
rect 25406 3476 25412 3528
rect 25464 3476 25470 3528
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3485 25559 3519
rect 25501 3479 25559 3485
rect 25516 3448 25544 3479
rect 23983 3420 25176 3448
rect 25240 3420 25544 3448
rect 23983 3417 23995 3420
rect 23937 3411 23995 3417
rect 14568 3352 14964 3380
rect 16390 3340 16396 3392
rect 16448 3340 16454 3392
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 19061 3383 19119 3389
rect 19061 3380 19073 3383
rect 17460 3352 19073 3380
rect 17460 3340 17466 3352
rect 19061 3349 19073 3352
rect 19107 3380 19119 3383
rect 19334 3380 19340 3392
rect 19107 3352 19340 3380
rect 19107 3349 19119 3352
rect 19061 3343 19119 3349
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 23750 3340 23756 3392
rect 23808 3340 23814 3392
rect 25148 3389 25176 3420
rect 25133 3383 25191 3389
rect 25133 3349 25145 3383
rect 25179 3349 25191 3383
rect 25133 3343 25191 3349
rect 1104 3290 26656 3312
rect 1104 3238 7298 3290
rect 7350 3238 7362 3290
rect 7414 3238 7426 3290
rect 7478 3238 7490 3290
rect 7542 3238 7554 3290
rect 7606 3238 13646 3290
rect 13698 3238 13710 3290
rect 13762 3238 13774 3290
rect 13826 3238 13838 3290
rect 13890 3238 13902 3290
rect 13954 3238 19994 3290
rect 20046 3238 20058 3290
rect 20110 3238 20122 3290
rect 20174 3238 20186 3290
rect 20238 3238 20250 3290
rect 20302 3238 26342 3290
rect 26394 3238 26406 3290
rect 26458 3238 26470 3290
rect 26522 3238 26534 3290
rect 26586 3238 26598 3290
rect 26650 3238 26656 3290
rect 1104 3216 26656 3238
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1820 3148 2145 3176
rect 1820 3136 1826 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 2682 3136 2688 3188
rect 2740 3136 2746 3188
rect 3234 3176 3240 3188
rect 3068 3148 3240 3176
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2700 3040 2728 3136
rect 3068 3117 3096 3148
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 4522 3136 4528 3188
rect 4580 3136 4586 3188
rect 4614 3136 4620 3188
rect 4672 3136 4678 3188
rect 4706 3136 4712 3188
rect 4764 3136 4770 3188
rect 4893 3179 4951 3185
rect 4893 3145 4905 3179
rect 4939 3176 4951 3179
rect 5166 3176 5172 3188
rect 4939 3148 5172 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 6086 3136 6092 3188
rect 6144 3176 6150 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 6144 3148 6377 3176
rect 6144 3136 6150 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 8110 3176 8116 3188
rect 7064 3148 8116 3176
rect 7064 3136 7070 3148
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8202 3136 8208 3188
rect 8260 3136 8266 3188
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8573 3179 8631 3185
rect 8573 3176 8585 3179
rect 8444 3148 8585 3176
rect 8444 3136 8450 3148
rect 8573 3145 8585 3148
rect 8619 3145 8631 3179
rect 8573 3139 8631 3145
rect 9214 3136 9220 3188
rect 9272 3136 9278 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10689 3179 10747 3185
rect 9824 3148 10640 3176
rect 9824 3136 9830 3148
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3077 3111 3111
rect 3053 3071 3111 3077
rect 2363 3012 2728 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4632 3040 4660 3136
rect 4724 3108 4752 3136
rect 4724 3080 4936 3108
rect 4908 3049 4936 3080
rect 6270 3068 6276 3120
rect 6328 3108 6334 3120
rect 7837 3111 7895 3117
rect 6328 3080 6670 3108
rect 6328 3068 6334 3080
rect 7837 3077 7849 3111
rect 7883 3108 7895 3111
rect 7926 3108 7932 3120
rect 7883 3080 7932 3108
rect 7883 3077 7895 3080
rect 7837 3071 7895 3077
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 4709 3043 4767 3049
rect 4709 3040 4721 3043
rect 4120 3026 4186 3040
rect 4120 3012 4200 3026
rect 4632 3012 4721 3040
rect 4120 3000 4126 3012
rect 4172 2972 4200 3012
rect 4709 3009 4721 3012
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 6288 2972 6316 3068
rect 8128 3049 8156 3136
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3009 8171 3043
rect 8312 3040 8340 3136
rect 9232 3108 9260 3136
rect 8680 3080 9260 3108
rect 8680 3049 8708 3080
rect 9490 3068 9496 3120
rect 9548 3068 9554 3120
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 8312 3012 8401 3040
rect 8113 3003 8171 3009
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 8754 3000 8760 3052
rect 8812 3000 8818 3052
rect 10612 3049 10640 3148
rect 10689 3145 10701 3179
rect 10735 3176 10747 3179
rect 10870 3176 10876 3188
rect 10735 3148 10876 3176
rect 10735 3145 10747 3148
rect 10689 3139 10747 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 11149 3179 11207 3185
rect 11149 3176 11161 3179
rect 11020 3148 11161 3176
rect 11020 3136 11026 3148
rect 11149 3145 11161 3148
rect 11195 3145 11207 3179
rect 11149 3139 11207 3145
rect 11790 3136 11796 3188
rect 11848 3136 11854 3188
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 12860 3148 13676 3176
rect 12860 3136 12866 3148
rect 11808 3108 11836 3136
rect 11348 3080 11836 3108
rect 11348 3049 11376 3080
rect 13354 3068 13360 3120
rect 13412 3068 13418 3120
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3009 11391 3043
rect 11333 3003 11391 3009
rect 11514 3000 11520 3052
rect 11572 3000 11578 3052
rect 12894 3000 12900 3052
rect 12952 3000 12958 3052
rect 13372 3040 13400 3068
rect 13648 3049 13676 3148
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14277 3179 14335 3185
rect 14277 3176 14289 3179
rect 13872 3148 14289 3176
rect 13872 3136 13878 3148
rect 14277 3145 14289 3148
rect 14323 3145 14335 3179
rect 15654 3176 15660 3188
rect 14277 3139 14335 3145
rect 15218 3148 15660 3176
rect 13955 3111 14013 3117
rect 13955 3077 13967 3111
rect 14001 3108 14013 3111
rect 14550 3108 14556 3120
rect 14001 3080 14556 3108
rect 14001 3077 14013 3080
rect 13955 3071 14013 3077
rect 14550 3068 14556 3080
rect 14608 3068 14614 3120
rect 15010 3068 15016 3120
rect 15068 3068 15074 3120
rect 15102 3068 15108 3120
rect 15160 3117 15166 3120
rect 15160 3111 15189 3117
rect 15177 3077 15189 3111
rect 15160 3071 15189 3077
rect 15160 3068 15166 3071
rect 13633 3043 13691 3049
rect 13372 3012 13584 3040
rect 4172 2944 6316 2972
rect 9030 2932 9036 2984
rect 9088 2932 9094 2984
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10505 2975 10563 2981
rect 10505 2972 10517 2975
rect 10284 2944 10517 2972
rect 10284 2932 10290 2944
rect 10505 2941 10517 2944
rect 10551 2941 10563 2975
rect 10505 2935 10563 2941
rect 11793 2975 11851 2981
rect 11793 2941 11805 2975
rect 11839 2972 11851 2975
rect 13449 2975 13507 2981
rect 13449 2972 13461 2975
rect 11839 2944 13461 2972
rect 11839 2941 11851 2944
rect 11793 2935 11851 2941
rect 13449 2941 13461 2944
rect 13495 2941 13507 2975
rect 13556 2972 13584 3012
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3040 14151 3043
rect 14274 3040 14280 3052
rect 14139 3012 14280 3040
rect 14139 3009 14151 3012
rect 14093 3003 14151 3009
rect 13740 2972 13768 3003
rect 13556 2944 13768 2972
rect 13832 2972 13860 3003
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3038 14979 3043
rect 15218 3040 15246 3148
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16390 3136 16396 3188
rect 16448 3136 16454 3188
rect 16666 3136 16672 3188
rect 16724 3136 16730 3188
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17644 3148 17785 3176
rect 17644 3136 17650 3148
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 20346 3176 20352 3188
rect 17773 3139 17831 3145
rect 20088 3148 20352 3176
rect 16408 3108 16436 3136
rect 15304 3080 16436 3108
rect 15304 3049 15332 3080
rect 18690 3068 18696 3120
rect 18748 3108 18754 3120
rect 20088 3117 20116 3148
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 21269 3179 21327 3185
rect 21269 3176 21281 3179
rect 20956 3148 21281 3176
rect 20956 3136 20962 3148
rect 21269 3145 21281 3148
rect 21315 3145 21327 3179
rect 21269 3139 21327 3145
rect 21818 3136 21824 3188
rect 21876 3136 21882 3188
rect 22646 3176 22652 3188
rect 22480 3148 22652 3176
rect 20073 3111 20131 3117
rect 18748 3080 18906 3108
rect 18748 3068 18754 3080
rect 20073 3077 20085 3111
rect 20119 3077 20131 3111
rect 20073 3071 20131 3077
rect 15120 3038 15246 3040
rect 14967 3012 15246 3038
rect 15289 3043 15347 3049
rect 14967 3010 15148 3012
rect 14967 3009 14979 3010
rect 14921 3003 14979 3009
rect 15289 3009 15301 3043
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 14182 2972 14188 2984
rect 13832 2944 14188 2972
rect 13449 2935 13507 2941
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 13262 2864 13268 2916
rect 13320 2864 13326 2916
rect 13998 2864 14004 2916
rect 14056 2904 14062 2916
rect 14384 2904 14412 3003
rect 14844 2972 14872 3003
rect 15838 3000 15844 3052
rect 15896 3000 15902 3052
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3040 16083 3043
rect 16114 3040 16120 3052
rect 16071 3012 16120 3040
rect 16071 3009 16083 3012
rect 16025 3003 16083 3009
rect 16040 2972 16068 3003
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17126 3000 17132 3052
rect 17184 3000 17190 3052
rect 20349 3043 20407 3049
rect 20349 3009 20361 3043
rect 20395 3040 20407 3043
rect 20622 3040 20628 3052
rect 20395 3012 20628 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 21453 3043 21511 3049
rect 21453 3009 21465 3043
rect 21499 3040 21511 3043
rect 21836 3040 21864 3136
rect 22480 3117 22508 3148
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 25682 3176 25688 3188
rect 23808 3148 25688 3176
rect 23808 3136 23814 3148
rect 25682 3136 25688 3148
rect 25740 3136 25746 3188
rect 22465 3111 22523 3117
rect 22465 3077 22477 3111
rect 22511 3077 22523 3111
rect 23768 3108 23796 3136
rect 23690 3080 23796 3108
rect 24213 3111 24271 3117
rect 22465 3071 22523 3077
rect 24213 3077 24225 3111
rect 24259 3108 24271 3111
rect 24302 3108 24308 3120
rect 24259 3080 24308 3108
rect 24259 3077 24271 3080
rect 24213 3071 24271 3077
rect 24302 3068 24308 3080
rect 24360 3068 24366 3120
rect 21499 3012 21864 3040
rect 21499 3009 21511 3012
rect 21453 3003 21511 3009
rect 14844 2944 16068 2972
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2972 17003 2975
rect 17402 2972 17408 2984
rect 16991 2944 17408 2972
rect 16991 2941 17003 2944
rect 16945 2935 17003 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 18322 2932 18328 2984
rect 18380 2932 18386 2984
rect 20640 2972 20668 3000
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 20640 2944 22201 2972
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 22189 2935 22247 2941
rect 14056 2876 14412 2904
rect 14645 2907 14703 2913
rect 14056 2864 14062 2876
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 14826 2904 14832 2916
rect 14691 2876 14832 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 17770 2904 17776 2916
rect 17052 2876 17776 2904
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 6178 2836 6184 2848
rect 3292 2808 6184 2836
rect 3292 2796 3298 2808
rect 6178 2796 6184 2808
rect 6236 2796 6242 2848
rect 16022 2796 16028 2848
rect 16080 2796 16086 2848
rect 17052 2845 17080 2876
rect 17770 2864 17776 2876
rect 17828 2904 17834 2916
rect 18601 2907 18659 2913
rect 18601 2904 18613 2907
rect 17828 2876 18613 2904
rect 17828 2864 17834 2876
rect 18601 2873 18613 2876
rect 18647 2873 18659 2907
rect 18601 2867 18659 2873
rect 17037 2839 17095 2845
rect 17037 2805 17049 2839
rect 17083 2805 17095 2839
rect 17037 2799 17095 2805
rect 17313 2839 17371 2845
rect 17313 2805 17325 2839
rect 17359 2836 17371 2839
rect 18506 2836 18512 2848
rect 17359 2808 18512 2836
rect 17359 2805 17371 2808
rect 17313 2799 17371 2805
rect 18506 2796 18512 2808
rect 18564 2796 18570 2848
rect 1104 2746 26496 2768
rect 1104 2694 4124 2746
rect 4176 2694 4188 2746
rect 4240 2694 4252 2746
rect 4304 2694 4316 2746
rect 4368 2694 4380 2746
rect 4432 2694 10472 2746
rect 10524 2694 10536 2746
rect 10588 2694 10600 2746
rect 10652 2694 10664 2746
rect 10716 2694 10728 2746
rect 10780 2694 16820 2746
rect 16872 2694 16884 2746
rect 16936 2694 16948 2746
rect 17000 2694 17012 2746
rect 17064 2694 17076 2746
rect 17128 2694 23168 2746
rect 23220 2694 23232 2746
rect 23284 2694 23296 2746
rect 23348 2694 23360 2746
rect 23412 2694 23424 2746
rect 23476 2694 26496 2746
rect 1104 2672 26496 2694
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 9088 2604 9137 2632
rect 9088 2592 9094 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 14553 2635 14611 2641
rect 14553 2601 14565 2635
rect 14599 2632 14611 2635
rect 14734 2632 14740 2644
rect 14599 2604 14740 2632
rect 14599 2601 14611 2604
rect 14553 2595 14611 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 17865 2635 17923 2641
rect 17865 2601 17877 2635
rect 17911 2632 17923 2635
rect 18322 2632 18328 2644
rect 17911 2604 18328 2632
rect 17911 2601 17923 2604
rect 17865 2595 17923 2601
rect 18322 2592 18328 2604
rect 18380 2592 18386 2644
rect 14090 2524 14096 2576
rect 14148 2564 14154 2576
rect 14369 2567 14427 2573
rect 14369 2564 14381 2567
rect 14148 2536 14381 2564
rect 14148 2524 14154 2536
rect 14369 2533 14381 2536
rect 14415 2533 14427 2567
rect 14369 2527 14427 2533
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10042 2496 10048 2508
rect 9815 2468 10048 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 14918 2456 14924 2508
rect 14976 2456 14982 2508
rect 16022 2456 16028 2508
rect 16080 2496 16086 2508
rect 18509 2499 18567 2505
rect 16080 2468 18184 2496
rect 16080 2456 16086 2468
rect 10410 2388 10416 2440
rect 10468 2388 10474 2440
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2428 14151 2431
rect 14936 2428 14964 2456
rect 18156 2440 18184 2468
rect 18509 2465 18521 2499
rect 18555 2496 18567 2499
rect 18782 2496 18788 2508
rect 18555 2468 18788 2496
rect 18555 2465 18567 2468
rect 18509 2459 18567 2465
rect 18782 2456 18788 2468
rect 18840 2456 18846 2508
rect 14139 2400 14964 2428
rect 14139 2397 14151 2400
rect 14093 2391 14151 2397
rect 18046 2388 18052 2440
rect 18104 2388 18110 2440
rect 18138 2388 18144 2440
rect 18196 2388 18202 2440
rect 18230 2388 18236 2440
rect 18288 2388 18294 2440
rect 19150 2428 19156 2440
rect 18340 2400 19156 2428
rect 18340 2369 18368 2400
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 25774 2388 25780 2440
rect 25832 2388 25838 2440
rect 18340 2363 18409 2369
rect 18340 2332 18363 2363
rect 18351 2329 18363 2332
rect 18397 2329 18409 2363
rect 18351 2323 18409 2329
rect 18506 2320 18512 2372
rect 18564 2360 18570 2372
rect 18693 2363 18751 2369
rect 18693 2360 18705 2363
rect 18564 2332 18705 2360
rect 18564 2320 18570 2332
rect 18693 2329 18705 2332
rect 18739 2329 18751 2363
rect 18693 2323 18751 2329
rect 26142 2320 26148 2372
rect 26200 2320 26206 2372
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18104 2264 18797 2292
rect 18104 2252 18110 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 1104 2202 26656 2224
rect 1104 2150 7298 2202
rect 7350 2150 7362 2202
rect 7414 2150 7426 2202
rect 7478 2150 7490 2202
rect 7542 2150 7554 2202
rect 7606 2150 13646 2202
rect 13698 2150 13710 2202
rect 13762 2150 13774 2202
rect 13826 2150 13838 2202
rect 13890 2150 13902 2202
rect 13954 2150 19994 2202
rect 20046 2150 20058 2202
rect 20110 2150 20122 2202
rect 20174 2150 20186 2202
rect 20238 2150 20250 2202
rect 20302 2150 26342 2202
rect 26394 2150 26406 2202
rect 26458 2150 26470 2202
rect 26522 2150 26534 2202
rect 26586 2150 26598 2202
rect 26650 2150 26656 2202
rect 1104 2128 26656 2150
<< via1 >>
rect 7298 27174 7350 27226
rect 7362 27174 7414 27226
rect 7426 27174 7478 27226
rect 7490 27174 7542 27226
rect 7554 27174 7606 27226
rect 13646 27174 13698 27226
rect 13710 27174 13762 27226
rect 13774 27174 13826 27226
rect 13838 27174 13890 27226
rect 13902 27174 13954 27226
rect 19994 27174 20046 27226
rect 20058 27174 20110 27226
rect 20122 27174 20174 27226
rect 20186 27174 20238 27226
rect 20250 27174 20302 27226
rect 26342 27174 26394 27226
rect 26406 27174 26458 27226
rect 26470 27174 26522 27226
rect 26534 27174 26586 27226
rect 26598 27174 26650 27226
rect 21180 27072 21232 27124
rect 17500 27004 17552 27056
rect 3884 26936 3936 26988
rect 11060 26979 11112 26988
rect 11060 26945 11069 26979
rect 11069 26945 11103 26979
rect 11103 26945 11112 26979
rect 11060 26936 11112 26945
rect 14832 26936 14884 26988
rect 16580 26936 16632 26988
rect 17224 26936 17276 26988
rect 21088 26936 21140 26988
rect 940 26868 992 26920
rect 20996 26911 21048 26920
rect 20996 26877 21005 26911
rect 21005 26877 21039 26911
rect 21039 26877 21048 26911
rect 20996 26868 21048 26877
rect 21456 26868 21508 26920
rect 21640 26868 21692 26920
rect 21824 26868 21876 26920
rect 16672 26732 16724 26784
rect 22560 26800 22612 26852
rect 4124 26630 4176 26682
rect 4188 26630 4240 26682
rect 4252 26630 4304 26682
rect 4316 26630 4368 26682
rect 4380 26630 4432 26682
rect 10472 26630 10524 26682
rect 10536 26630 10588 26682
rect 10600 26630 10652 26682
rect 10664 26630 10716 26682
rect 10728 26630 10780 26682
rect 16820 26630 16872 26682
rect 16884 26630 16936 26682
rect 16948 26630 17000 26682
rect 17012 26630 17064 26682
rect 17076 26630 17128 26682
rect 23168 26630 23220 26682
rect 23232 26630 23284 26682
rect 23296 26630 23348 26682
rect 23360 26630 23412 26682
rect 23424 26630 23476 26682
rect 16212 26392 16264 26444
rect 16580 26528 16632 26580
rect 17408 26528 17460 26580
rect 17500 26571 17552 26580
rect 17500 26537 17509 26571
rect 17509 26537 17543 26571
rect 17543 26537 17552 26571
rect 17500 26528 17552 26537
rect 20996 26528 21048 26580
rect 21456 26528 21508 26580
rect 16580 26392 16632 26444
rect 22100 26392 22152 26444
rect 9496 26367 9548 26376
rect 9496 26333 9505 26367
rect 9505 26333 9539 26367
rect 9539 26333 9548 26367
rect 9496 26324 9548 26333
rect 11428 26367 11480 26376
rect 11428 26333 11437 26367
rect 11437 26333 11471 26367
rect 11471 26333 11480 26367
rect 11428 26324 11480 26333
rect 12532 26367 12584 26376
rect 12532 26333 12541 26367
rect 12541 26333 12575 26367
rect 12575 26333 12584 26367
rect 12532 26324 12584 26333
rect 12900 26324 12952 26376
rect 16028 26367 16080 26376
rect 16028 26333 16037 26367
rect 16037 26333 16071 26367
rect 16071 26333 16080 26367
rect 16028 26324 16080 26333
rect 16120 26367 16172 26376
rect 16120 26333 16129 26367
rect 16129 26333 16163 26367
rect 16163 26333 16172 26367
rect 16120 26324 16172 26333
rect 16764 26367 16816 26376
rect 16764 26333 16773 26367
rect 16773 26333 16807 26367
rect 16807 26333 16816 26367
rect 16764 26324 16816 26333
rect 18052 26367 18104 26376
rect 18052 26333 18061 26367
rect 18061 26333 18095 26367
rect 18095 26333 18104 26367
rect 18052 26324 18104 26333
rect 19616 26324 19668 26376
rect 19708 26367 19760 26376
rect 19708 26333 19717 26367
rect 19717 26333 19751 26367
rect 19751 26333 19760 26367
rect 19708 26324 19760 26333
rect 21272 26367 21324 26376
rect 16488 26299 16540 26308
rect 16488 26265 16513 26299
rect 16513 26265 16540 26299
rect 21272 26333 21281 26367
rect 21281 26333 21315 26367
rect 21315 26333 21324 26367
rect 21272 26324 21324 26333
rect 22376 26367 22428 26376
rect 22376 26333 22385 26367
rect 22385 26333 22419 26367
rect 22419 26333 22428 26367
rect 22376 26324 22428 26333
rect 16488 26256 16540 26265
rect 9312 26231 9364 26240
rect 9312 26197 9321 26231
rect 9321 26197 9355 26231
rect 9355 26197 9364 26231
rect 9312 26188 9364 26197
rect 10324 26188 10376 26240
rect 12624 26231 12676 26240
rect 12624 26197 12633 26231
rect 12633 26197 12667 26231
rect 12667 26197 12676 26231
rect 12624 26188 12676 26197
rect 15660 26231 15712 26240
rect 15660 26197 15669 26231
rect 15669 26197 15703 26231
rect 15703 26197 15712 26231
rect 15660 26188 15712 26197
rect 19248 26231 19300 26240
rect 19248 26197 19257 26231
rect 19257 26197 19291 26231
rect 19291 26197 19300 26231
rect 19248 26188 19300 26197
rect 19892 26188 19944 26240
rect 21732 26231 21784 26240
rect 21732 26197 21741 26231
rect 21741 26197 21775 26231
rect 21775 26197 21784 26231
rect 21732 26188 21784 26197
rect 22468 26231 22520 26240
rect 22468 26197 22477 26231
rect 22477 26197 22511 26231
rect 22511 26197 22520 26231
rect 22468 26188 22520 26197
rect 7298 26086 7350 26138
rect 7362 26086 7414 26138
rect 7426 26086 7478 26138
rect 7490 26086 7542 26138
rect 7554 26086 7606 26138
rect 13646 26086 13698 26138
rect 13710 26086 13762 26138
rect 13774 26086 13826 26138
rect 13838 26086 13890 26138
rect 13902 26086 13954 26138
rect 19994 26086 20046 26138
rect 20058 26086 20110 26138
rect 20122 26086 20174 26138
rect 20186 26086 20238 26138
rect 20250 26086 20302 26138
rect 26342 26086 26394 26138
rect 26406 26086 26458 26138
rect 26470 26086 26522 26138
rect 26534 26086 26586 26138
rect 26598 26086 26650 26138
rect 8116 25848 8168 25900
rect 9312 25848 9364 25900
rect 9956 25891 10008 25900
rect 9956 25857 9990 25891
rect 9990 25857 10008 25891
rect 9956 25848 10008 25857
rect 10968 25848 11020 25900
rect 11336 25891 11388 25900
rect 11336 25857 11345 25891
rect 11345 25857 11379 25891
rect 11379 25857 11388 25891
rect 11336 25848 11388 25857
rect 12348 25891 12400 25900
rect 12348 25857 12357 25891
rect 12357 25857 12391 25891
rect 12391 25857 12400 25891
rect 12348 25848 12400 25857
rect 11244 25780 11296 25832
rect 12256 25780 12308 25832
rect 11428 25712 11480 25764
rect 12440 25712 12492 25764
rect 9864 25644 9916 25696
rect 11152 25687 11204 25696
rect 11152 25653 11161 25687
rect 11161 25653 11195 25687
rect 11195 25653 11204 25687
rect 11152 25644 11204 25653
rect 11796 25687 11848 25696
rect 11796 25653 11805 25687
rect 11805 25653 11839 25687
rect 11839 25653 11848 25687
rect 11796 25644 11848 25653
rect 11980 25644 12032 25696
rect 12256 25644 12308 25696
rect 13360 25891 13412 25900
rect 13360 25857 13366 25891
rect 13366 25857 13400 25891
rect 13400 25857 13412 25891
rect 13360 25848 13412 25857
rect 13544 25959 13596 25968
rect 13544 25925 13553 25959
rect 13553 25925 13587 25959
rect 13587 25925 13596 25959
rect 13544 25916 13596 25925
rect 15936 25984 15988 26036
rect 14556 25916 14608 25968
rect 15752 25916 15804 25968
rect 16120 25916 16172 25968
rect 15016 25848 15068 25900
rect 16028 25848 16080 25900
rect 16212 25891 16264 25900
rect 16212 25857 16221 25891
rect 16221 25857 16255 25891
rect 16255 25857 16264 25891
rect 16212 25848 16264 25857
rect 13544 25712 13596 25764
rect 14464 25823 14516 25832
rect 14464 25789 14473 25823
rect 14473 25789 14507 25823
rect 14507 25789 14516 25823
rect 14464 25780 14516 25789
rect 13636 25687 13688 25696
rect 13636 25653 13645 25687
rect 13645 25653 13679 25687
rect 13679 25653 13688 25687
rect 13636 25644 13688 25653
rect 14280 25644 14332 25696
rect 14832 25687 14884 25696
rect 14832 25653 14841 25687
rect 14841 25653 14875 25687
rect 14875 25653 14884 25687
rect 14832 25644 14884 25653
rect 14924 25687 14976 25696
rect 14924 25653 14933 25687
rect 14933 25653 14967 25687
rect 14967 25653 14976 25687
rect 14924 25644 14976 25653
rect 16396 25644 16448 25696
rect 16764 25984 16816 26036
rect 21732 25984 21784 26036
rect 21824 26027 21876 26036
rect 21824 25993 21833 26027
rect 21833 25993 21867 26027
rect 21867 25993 21876 26027
rect 21824 25984 21876 25993
rect 19248 25916 19300 25968
rect 17500 25848 17552 25900
rect 19156 25848 19208 25900
rect 22468 25916 22520 25968
rect 22560 25916 22612 25968
rect 22744 25916 22796 25968
rect 20352 25848 20404 25900
rect 20812 25780 20864 25832
rect 21088 25891 21140 25900
rect 21088 25857 21097 25891
rect 21097 25857 21131 25891
rect 21131 25857 21140 25891
rect 21088 25848 21140 25857
rect 21180 25891 21232 25900
rect 21180 25857 21189 25891
rect 21189 25857 21223 25891
rect 21223 25857 21232 25891
rect 21180 25848 21232 25857
rect 21272 25891 21324 25900
rect 21272 25857 21281 25891
rect 21281 25857 21315 25891
rect 21315 25857 21324 25891
rect 21272 25848 21324 25857
rect 21824 25848 21876 25900
rect 19708 25644 19760 25696
rect 19892 25644 19944 25696
rect 21456 25712 21508 25764
rect 20812 25687 20864 25696
rect 20812 25653 20821 25687
rect 20821 25653 20855 25687
rect 20855 25653 20864 25687
rect 20812 25644 20864 25653
rect 21088 25644 21140 25696
rect 4124 25542 4176 25594
rect 4188 25542 4240 25594
rect 4252 25542 4304 25594
rect 4316 25542 4368 25594
rect 4380 25542 4432 25594
rect 10472 25542 10524 25594
rect 10536 25542 10588 25594
rect 10600 25542 10652 25594
rect 10664 25542 10716 25594
rect 10728 25542 10780 25594
rect 16820 25542 16872 25594
rect 16884 25542 16936 25594
rect 16948 25542 17000 25594
rect 17012 25542 17064 25594
rect 17076 25542 17128 25594
rect 23168 25542 23220 25594
rect 23232 25542 23284 25594
rect 23296 25542 23348 25594
rect 23360 25542 23412 25594
rect 23424 25542 23476 25594
rect 9496 25483 9548 25492
rect 9496 25449 9505 25483
rect 9505 25449 9539 25483
rect 9539 25449 9548 25483
rect 9496 25440 9548 25449
rect 9772 25440 9824 25492
rect 9956 25483 10008 25492
rect 9956 25449 9965 25483
rect 9965 25449 9999 25483
rect 9999 25449 10008 25483
rect 9956 25440 10008 25449
rect 12440 25440 12492 25492
rect 14280 25440 14332 25492
rect 10232 25279 10284 25288
rect 10232 25245 10241 25279
rect 10241 25245 10275 25279
rect 10275 25245 10284 25279
rect 10232 25236 10284 25245
rect 10416 25279 10468 25288
rect 10416 25245 10425 25279
rect 10425 25245 10459 25279
rect 10459 25245 10468 25279
rect 10416 25236 10468 25245
rect 9864 25211 9916 25220
rect 9864 25177 9873 25211
rect 9873 25177 9907 25211
rect 9907 25177 9916 25211
rect 9864 25168 9916 25177
rect 10140 25168 10192 25220
rect 10324 25168 10376 25220
rect 11244 25236 11296 25288
rect 12624 25236 12676 25288
rect 11152 25168 11204 25220
rect 14188 25304 14240 25356
rect 14556 25372 14608 25424
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 14464 25279 14516 25288
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 15016 25440 15068 25492
rect 16028 25372 16080 25424
rect 18052 25440 18104 25492
rect 20720 25440 20772 25492
rect 20812 25440 20864 25492
rect 22376 25440 22428 25492
rect 14740 25279 14792 25288
rect 14740 25245 14749 25279
rect 14749 25245 14783 25279
rect 14783 25245 14792 25279
rect 14740 25236 14792 25245
rect 16120 25236 16172 25288
rect 16304 25236 16356 25288
rect 10600 25100 10652 25152
rect 10784 25100 10836 25152
rect 12256 25100 12308 25152
rect 13452 25143 13504 25152
rect 13452 25109 13461 25143
rect 13461 25109 13495 25143
rect 13495 25109 13504 25143
rect 13452 25100 13504 25109
rect 14004 25100 14056 25152
rect 14832 25168 14884 25220
rect 15660 25168 15712 25220
rect 16212 25100 16264 25152
rect 16672 25168 16724 25220
rect 17316 25236 17368 25288
rect 19156 25236 19208 25288
rect 19340 25236 19392 25288
rect 20628 25236 20680 25288
rect 18052 25143 18104 25152
rect 18052 25109 18061 25143
rect 18061 25109 18095 25143
rect 18095 25109 18104 25143
rect 18052 25100 18104 25109
rect 18604 25143 18656 25152
rect 18604 25109 18613 25143
rect 18613 25109 18647 25143
rect 18647 25109 18656 25143
rect 18604 25100 18656 25109
rect 19524 25211 19576 25220
rect 19524 25177 19558 25211
rect 19558 25177 19576 25211
rect 19524 25168 19576 25177
rect 19800 25168 19852 25220
rect 20904 25279 20956 25288
rect 20904 25245 20913 25279
rect 20913 25245 20947 25279
rect 20947 25245 20956 25279
rect 20904 25236 20956 25245
rect 21088 25279 21140 25288
rect 21088 25245 21097 25279
rect 21097 25245 21131 25279
rect 21131 25245 21140 25279
rect 21088 25236 21140 25245
rect 22744 25236 22796 25288
rect 20352 25100 20404 25152
rect 20996 25100 21048 25152
rect 7298 24998 7350 25050
rect 7362 24998 7414 25050
rect 7426 24998 7478 25050
rect 7490 24998 7542 25050
rect 7554 24998 7606 25050
rect 13646 24998 13698 25050
rect 13710 24998 13762 25050
rect 13774 24998 13826 25050
rect 13838 24998 13890 25050
rect 13902 24998 13954 25050
rect 19994 24998 20046 25050
rect 20058 24998 20110 25050
rect 20122 24998 20174 25050
rect 20186 24998 20238 25050
rect 20250 24998 20302 25050
rect 26342 24998 26394 25050
rect 26406 24998 26458 25050
rect 26470 24998 26522 25050
rect 26534 24998 26586 25050
rect 26598 24998 26650 25050
rect 10600 24939 10652 24948
rect 10600 24905 10609 24939
rect 10609 24905 10643 24939
rect 10643 24905 10652 24939
rect 10600 24896 10652 24905
rect 11336 24939 11388 24948
rect 11336 24905 11345 24939
rect 11345 24905 11379 24939
rect 11379 24905 11388 24939
rect 11336 24896 11388 24905
rect 12624 24896 12676 24948
rect 13360 24896 13412 24948
rect 14464 24896 14516 24948
rect 14924 24896 14976 24948
rect 15752 24939 15804 24948
rect 15752 24905 15761 24939
rect 15761 24905 15795 24939
rect 15795 24905 15804 24939
rect 15752 24896 15804 24905
rect 15936 24939 15988 24948
rect 15936 24905 15945 24939
rect 15945 24905 15979 24939
rect 15979 24905 15988 24939
rect 15936 24896 15988 24905
rect 16028 24896 16080 24948
rect 16212 24896 16264 24948
rect 16396 24896 16448 24948
rect 17500 24896 17552 24948
rect 19340 24896 19392 24948
rect 21088 24896 21140 24948
rect 9864 24828 9916 24880
rect 10232 24828 10284 24880
rect 9128 24803 9180 24812
rect 9128 24769 9137 24803
rect 9137 24769 9171 24803
rect 9171 24769 9180 24803
rect 9128 24760 9180 24769
rect 9588 24803 9640 24812
rect 9588 24769 9597 24803
rect 9597 24769 9631 24803
rect 9631 24769 9640 24803
rect 9588 24760 9640 24769
rect 9680 24692 9732 24744
rect 10232 24692 10284 24744
rect 10048 24624 10100 24676
rect 11980 24760 12032 24812
rect 12256 24803 12308 24812
rect 12256 24769 12265 24803
rect 12265 24769 12299 24803
rect 12299 24769 12308 24803
rect 12256 24760 12308 24769
rect 13084 24871 13136 24880
rect 13084 24837 13093 24871
rect 13093 24837 13127 24871
rect 13127 24837 13136 24871
rect 13084 24828 13136 24837
rect 10876 24692 10928 24744
rect 9956 24599 10008 24608
rect 9956 24565 9965 24599
rect 9965 24565 9999 24599
rect 9999 24565 10008 24599
rect 9956 24556 10008 24565
rect 10140 24599 10192 24608
rect 10140 24565 10149 24599
rect 10149 24565 10183 24599
rect 10183 24565 10192 24599
rect 10140 24556 10192 24565
rect 10968 24556 11020 24608
rect 11152 24556 11204 24608
rect 12532 24692 12584 24744
rect 12624 24735 12676 24744
rect 12624 24701 12633 24735
rect 12633 24701 12667 24735
rect 12667 24701 12676 24735
rect 12624 24692 12676 24701
rect 12716 24735 12768 24744
rect 12716 24701 12725 24735
rect 12725 24701 12759 24735
rect 12759 24701 12768 24735
rect 12716 24692 12768 24701
rect 13360 24692 13412 24744
rect 13452 24624 13504 24676
rect 14280 24760 14332 24812
rect 14648 24803 14700 24812
rect 14648 24769 14682 24803
rect 14682 24769 14700 24803
rect 14648 24760 14700 24769
rect 17224 24871 17276 24880
rect 17224 24837 17233 24871
rect 17233 24837 17267 24871
rect 17267 24837 17276 24871
rect 17224 24828 17276 24837
rect 18604 24871 18656 24880
rect 18604 24837 18638 24871
rect 18638 24837 18656 24871
rect 18604 24828 18656 24837
rect 19892 24828 19944 24880
rect 16580 24760 16632 24812
rect 17592 24760 17644 24812
rect 18052 24760 18104 24812
rect 19156 24760 19208 24812
rect 22376 24896 22428 24948
rect 14740 24556 14792 24608
rect 16120 24556 16172 24608
rect 18328 24735 18380 24744
rect 18328 24701 18337 24735
rect 18337 24701 18371 24735
rect 18371 24701 18380 24735
rect 18328 24692 18380 24701
rect 17408 24667 17460 24676
rect 17408 24633 17417 24667
rect 17417 24633 17451 24667
rect 17451 24633 17460 24667
rect 17408 24624 17460 24633
rect 20536 24692 20588 24744
rect 18144 24556 18196 24608
rect 20536 24599 20588 24608
rect 20536 24565 20545 24599
rect 20545 24565 20579 24599
rect 20579 24565 20588 24599
rect 20536 24556 20588 24565
rect 21180 24692 21232 24744
rect 22284 24624 22336 24676
rect 23020 24624 23072 24676
rect 22008 24599 22060 24608
rect 22008 24565 22017 24599
rect 22017 24565 22051 24599
rect 22051 24565 22060 24599
rect 22008 24556 22060 24565
rect 4124 24454 4176 24506
rect 4188 24454 4240 24506
rect 4252 24454 4304 24506
rect 4316 24454 4368 24506
rect 4380 24454 4432 24506
rect 10472 24454 10524 24506
rect 10536 24454 10588 24506
rect 10600 24454 10652 24506
rect 10664 24454 10716 24506
rect 10728 24454 10780 24506
rect 16820 24454 16872 24506
rect 16884 24454 16936 24506
rect 16948 24454 17000 24506
rect 17012 24454 17064 24506
rect 17076 24454 17128 24506
rect 23168 24454 23220 24506
rect 23232 24454 23284 24506
rect 23296 24454 23348 24506
rect 23360 24454 23412 24506
rect 23424 24454 23476 24506
rect 9128 24352 9180 24404
rect 9680 24352 9732 24404
rect 10140 24352 10192 24404
rect 12900 24395 12952 24404
rect 12900 24361 12909 24395
rect 12909 24361 12943 24395
rect 12943 24361 12952 24395
rect 12900 24352 12952 24361
rect 13084 24352 13136 24404
rect 13360 24352 13412 24404
rect 14648 24395 14700 24404
rect 14648 24361 14657 24395
rect 14657 24361 14691 24395
rect 14691 24361 14700 24395
rect 14648 24352 14700 24361
rect 16120 24395 16172 24404
rect 16120 24361 16129 24395
rect 16129 24361 16163 24395
rect 16163 24361 16172 24395
rect 16120 24352 16172 24361
rect 19524 24352 19576 24404
rect 19616 24352 19668 24404
rect 20536 24352 20588 24404
rect 9588 24284 9640 24336
rect 9772 24284 9824 24336
rect 10876 24284 10928 24336
rect 10968 24284 11020 24336
rect 12532 24284 12584 24336
rect 8116 24148 8168 24200
rect 9404 24148 9456 24200
rect 10232 24191 10284 24200
rect 10232 24157 10241 24191
rect 10241 24157 10275 24191
rect 10275 24157 10284 24191
rect 10232 24148 10284 24157
rect 11796 24259 11848 24268
rect 11796 24225 11805 24259
rect 11805 24225 11839 24259
rect 11839 24225 11848 24259
rect 11796 24216 11848 24225
rect 11152 24148 11204 24200
rect 12624 24191 12676 24200
rect 12624 24157 12633 24191
rect 12633 24157 12667 24191
rect 12667 24157 12676 24191
rect 12624 24148 12676 24157
rect 16304 24284 16356 24336
rect 14004 24216 14056 24268
rect 16212 24216 16264 24268
rect 16488 24216 16540 24268
rect 19708 24284 19760 24336
rect 19524 24216 19576 24268
rect 20628 24216 20680 24268
rect 7748 24080 7800 24132
rect 12716 24123 12768 24132
rect 12716 24089 12725 24123
rect 12725 24089 12759 24123
rect 12759 24089 12768 24123
rect 12716 24080 12768 24089
rect 19800 24148 19852 24200
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 19892 24080 19944 24132
rect 19800 24012 19852 24064
rect 22376 24148 22428 24200
rect 23020 24148 23072 24200
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 23296 24191 23348 24200
rect 23296 24157 23305 24191
rect 23305 24157 23339 24191
rect 23339 24157 23348 24191
rect 23296 24148 23348 24157
rect 26148 24191 26200 24200
rect 26148 24157 26157 24191
rect 26157 24157 26191 24191
rect 26191 24157 26200 24191
rect 26148 24148 26200 24157
rect 22468 24012 22520 24064
rect 7298 23910 7350 23962
rect 7362 23910 7414 23962
rect 7426 23910 7478 23962
rect 7490 23910 7542 23962
rect 7554 23910 7606 23962
rect 13646 23910 13698 23962
rect 13710 23910 13762 23962
rect 13774 23910 13826 23962
rect 13838 23910 13890 23962
rect 13902 23910 13954 23962
rect 19994 23910 20046 23962
rect 20058 23910 20110 23962
rect 20122 23910 20174 23962
rect 20186 23910 20238 23962
rect 20250 23910 20302 23962
rect 26342 23910 26394 23962
rect 26406 23910 26458 23962
rect 26470 23910 26522 23962
rect 26534 23910 26586 23962
rect 26598 23910 26650 23962
rect 7748 23851 7800 23860
rect 7748 23817 7757 23851
rect 7757 23817 7791 23851
rect 7791 23817 7800 23851
rect 7748 23808 7800 23817
rect 9772 23808 9824 23860
rect 10048 23808 10100 23860
rect 8116 23672 8168 23724
rect 10324 23715 10376 23724
rect 10324 23681 10333 23715
rect 10333 23681 10367 23715
rect 10367 23681 10376 23715
rect 10324 23672 10376 23681
rect 16028 23672 16080 23724
rect 22468 23740 22520 23792
rect 9404 23511 9456 23520
rect 9404 23477 9413 23511
rect 9413 23477 9447 23511
rect 9447 23477 9456 23511
rect 9404 23468 9456 23477
rect 9956 23536 10008 23588
rect 10140 23536 10192 23588
rect 14556 23604 14608 23656
rect 15384 23647 15436 23656
rect 15384 23613 15393 23647
rect 15393 23613 15427 23647
rect 15427 23613 15436 23647
rect 15384 23604 15436 23613
rect 20352 23604 20404 23656
rect 22284 23715 22336 23724
rect 22284 23681 22293 23715
rect 22293 23681 22327 23715
rect 22327 23681 22336 23715
rect 22284 23672 22336 23681
rect 22376 23715 22428 23724
rect 22376 23681 22385 23715
rect 22385 23681 22419 23715
rect 22419 23681 22428 23715
rect 22376 23672 22428 23681
rect 23296 23808 23348 23860
rect 23572 23808 23624 23860
rect 15476 23536 15528 23588
rect 14648 23511 14700 23520
rect 14648 23477 14657 23511
rect 14657 23477 14691 23511
rect 14691 23477 14700 23511
rect 14648 23468 14700 23477
rect 15108 23468 15160 23520
rect 18144 23468 18196 23520
rect 19064 23511 19116 23520
rect 19064 23477 19073 23511
rect 19073 23477 19107 23511
rect 19107 23477 19116 23511
rect 19064 23468 19116 23477
rect 24768 23715 24820 23724
rect 24768 23681 24777 23715
rect 24777 23681 24811 23715
rect 24811 23681 24820 23715
rect 24768 23672 24820 23681
rect 22744 23647 22796 23656
rect 22744 23613 22753 23647
rect 22753 23613 22787 23647
rect 22787 23613 22796 23647
rect 22744 23604 22796 23613
rect 4124 23366 4176 23418
rect 4188 23366 4240 23418
rect 4252 23366 4304 23418
rect 4316 23366 4368 23418
rect 4380 23366 4432 23418
rect 10472 23366 10524 23418
rect 10536 23366 10588 23418
rect 10600 23366 10652 23418
rect 10664 23366 10716 23418
rect 10728 23366 10780 23418
rect 16820 23366 16872 23418
rect 16884 23366 16936 23418
rect 16948 23366 17000 23418
rect 17012 23366 17064 23418
rect 17076 23366 17128 23418
rect 23168 23366 23220 23418
rect 23232 23366 23284 23418
rect 23296 23366 23348 23418
rect 23360 23366 23412 23418
rect 23424 23366 23476 23418
rect 10048 23196 10100 23248
rect 9404 23171 9456 23180
rect 9404 23137 9413 23171
rect 9413 23137 9447 23171
rect 9447 23137 9456 23171
rect 9404 23128 9456 23137
rect 10232 23128 10284 23180
rect 9588 23060 9640 23112
rect 11152 23239 11204 23248
rect 11152 23205 11161 23239
rect 11161 23205 11195 23239
rect 11195 23205 11204 23239
rect 11152 23196 11204 23205
rect 14280 23264 14332 23316
rect 15108 23264 15160 23316
rect 13084 23196 13136 23248
rect 9956 22992 10008 23044
rect 11152 23060 11204 23112
rect 11704 23103 11756 23112
rect 11704 23069 11713 23103
rect 11713 23069 11747 23103
rect 11747 23069 11756 23103
rect 11704 23060 11756 23069
rect 11796 23060 11848 23112
rect 12164 23103 12216 23112
rect 12164 23069 12173 23103
rect 12173 23069 12207 23103
rect 12207 23069 12216 23103
rect 12164 23060 12216 23069
rect 9680 22967 9732 22976
rect 9680 22933 9689 22967
rect 9689 22933 9723 22967
rect 9723 22933 9732 22967
rect 9680 22924 9732 22933
rect 12992 22992 13044 23044
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 14188 23103 14240 23112
rect 14188 23069 14197 23103
rect 14197 23069 14231 23103
rect 14231 23069 14240 23103
rect 14188 23060 14240 23069
rect 14924 23103 14976 23112
rect 14924 23069 14933 23103
rect 14933 23069 14967 23103
rect 14967 23069 14976 23103
rect 14924 23060 14976 23069
rect 15568 23103 15620 23112
rect 15568 23069 15577 23103
rect 15577 23069 15611 23103
rect 15611 23069 15620 23103
rect 15568 23060 15620 23069
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 20904 23264 20956 23316
rect 23296 23264 23348 23316
rect 19524 23196 19576 23248
rect 21916 23196 21968 23248
rect 22284 23196 22336 23248
rect 22652 23196 22704 23248
rect 19892 23128 19944 23180
rect 16488 22992 16540 23044
rect 17684 22992 17736 23044
rect 18052 23060 18104 23112
rect 18144 23103 18196 23112
rect 18144 23069 18153 23103
rect 18153 23069 18187 23103
rect 18187 23069 18196 23103
rect 18144 23060 18196 23069
rect 18236 23060 18288 23112
rect 19064 23060 19116 23112
rect 20352 23103 20404 23112
rect 20352 23069 20361 23103
rect 20361 23069 20395 23103
rect 20395 23069 20404 23103
rect 20352 23060 20404 23069
rect 20812 23060 20864 23112
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 22100 23103 22152 23112
rect 22100 23069 22114 23103
rect 22114 23069 22148 23103
rect 22148 23069 22152 23103
rect 22100 23060 22152 23069
rect 22284 23060 22336 23112
rect 21916 23035 21968 23044
rect 21916 23001 21925 23035
rect 21925 23001 21959 23035
rect 21959 23001 21968 23035
rect 21916 22992 21968 23001
rect 22192 22992 22244 23044
rect 22560 23103 22612 23112
rect 22560 23069 22569 23103
rect 22569 23069 22603 23103
rect 22603 23069 22612 23103
rect 22560 23060 22612 23069
rect 22744 23060 22796 23112
rect 24032 23128 24084 23180
rect 24768 23171 24820 23180
rect 24768 23137 24777 23171
rect 24777 23137 24811 23171
rect 24811 23137 24820 23171
rect 24768 23128 24820 23137
rect 24676 23103 24728 23112
rect 24676 23069 24685 23103
rect 24685 23069 24719 23103
rect 24719 23069 24728 23103
rect 24676 23060 24728 23069
rect 22928 23035 22980 23044
rect 22928 23001 22962 23035
rect 22962 23001 22980 23035
rect 22928 22992 22980 23001
rect 25320 23103 25372 23112
rect 25320 23069 25329 23103
rect 25329 23069 25363 23103
rect 25363 23069 25372 23103
rect 25320 23060 25372 23069
rect 11980 22967 12032 22976
rect 11980 22933 11989 22967
rect 11989 22933 12023 22967
rect 12023 22933 12032 22967
rect 11980 22924 12032 22933
rect 15016 22967 15068 22976
rect 15016 22933 15025 22967
rect 15025 22933 15059 22967
rect 15059 22933 15068 22967
rect 15016 22924 15068 22933
rect 16212 22924 16264 22976
rect 16672 22924 16724 22976
rect 17408 22924 17460 22976
rect 17960 22924 18012 22976
rect 19248 22967 19300 22976
rect 19248 22933 19257 22967
rect 19257 22933 19291 22967
rect 19291 22933 19300 22967
rect 19248 22924 19300 22933
rect 20444 22967 20496 22976
rect 20444 22933 20453 22967
rect 20453 22933 20487 22967
rect 20487 22933 20496 22967
rect 20444 22924 20496 22933
rect 22284 22967 22336 22976
rect 22284 22933 22293 22967
rect 22293 22933 22327 22967
rect 22327 22933 22336 22967
rect 22284 22924 22336 22933
rect 22468 22967 22520 22976
rect 22468 22933 22477 22967
rect 22477 22933 22511 22967
rect 22511 22933 22520 22967
rect 22468 22924 22520 22933
rect 22836 22924 22888 22976
rect 23664 22924 23716 22976
rect 24952 22992 25004 23044
rect 24124 22924 24176 22976
rect 25136 22967 25188 22976
rect 25136 22933 25145 22967
rect 25145 22933 25179 22967
rect 25179 22933 25188 22967
rect 25136 22924 25188 22933
rect 7298 22822 7350 22874
rect 7362 22822 7414 22874
rect 7426 22822 7478 22874
rect 7490 22822 7542 22874
rect 7554 22822 7606 22874
rect 13646 22822 13698 22874
rect 13710 22822 13762 22874
rect 13774 22822 13826 22874
rect 13838 22822 13890 22874
rect 13902 22822 13954 22874
rect 19994 22822 20046 22874
rect 20058 22822 20110 22874
rect 20122 22822 20174 22874
rect 20186 22822 20238 22874
rect 20250 22822 20302 22874
rect 26342 22822 26394 22874
rect 26406 22822 26458 22874
rect 26470 22822 26522 22874
rect 26534 22822 26586 22874
rect 26598 22822 26650 22874
rect 9680 22720 9732 22772
rect 9956 22763 10008 22772
rect 9956 22729 9965 22763
rect 9965 22729 9999 22763
rect 9999 22729 10008 22763
rect 9956 22720 10008 22729
rect 11152 22720 11204 22772
rect 11796 22720 11848 22772
rect 11980 22720 12032 22772
rect 12164 22720 12216 22772
rect 13360 22720 13412 22772
rect 8116 22584 8168 22636
rect 9312 22584 9364 22636
rect 9956 22584 10008 22636
rect 11244 22584 11296 22636
rect 11704 22584 11756 22636
rect 12532 22652 12584 22704
rect 13452 22652 13504 22704
rect 12164 22584 12216 22636
rect 15568 22720 15620 22772
rect 16028 22720 16080 22772
rect 15384 22652 15436 22704
rect 20444 22720 20496 22772
rect 14004 22627 14056 22636
rect 14004 22593 14038 22627
rect 14038 22593 14056 22627
rect 12992 22516 13044 22568
rect 14004 22584 14056 22593
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 16212 22584 16264 22636
rect 16672 22584 16724 22636
rect 18328 22652 18380 22704
rect 19248 22584 19300 22636
rect 19800 22584 19852 22636
rect 13728 22559 13780 22568
rect 13728 22525 13737 22559
rect 13737 22525 13771 22559
rect 13771 22525 13780 22559
rect 13728 22516 13780 22525
rect 22008 22652 22060 22704
rect 22284 22720 22336 22772
rect 22468 22720 22520 22772
rect 22560 22720 22612 22772
rect 23572 22763 23624 22772
rect 23572 22729 23581 22763
rect 23581 22729 23615 22763
rect 23615 22729 23624 22763
rect 23572 22720 23624 22729
rect 23664 22763 23716 22772
rect 23664 22729 23673 22763
rect 23673 22729 23707 22763
rect 23707 22729 23716 22763
rect 23664 22720 23716 22729
rect 24216 22720 24268 22772
rect 24492 22720 24544 22772
rect 25780 22720 25832 22772
rect 16580 22516 16632 22568
rect 16764 22559 16816 22568
rect 16764 22525 16773 22559
rect 16773 22525 16807 22559
rect 16807 22525 16816 22559
rect 16764 22516 16816 22525
rect 21272 22516 21324 22568
rect 22284 22584 22336 22636
rect 24032 22652 24084 22704
rect 22652 22516 22704 22568
rect 22836 22627 22888 22636
rect 22836 22593 22845 22627
rect 22845 22593 22879 22627
rect 22879 22593 22888 22627
rect 22836 22584 22888 22593
rect 10048 22423 10100 22432
rect 10048 22389 10057 22423
rect 10057 22389 10091 22423
rect 10091 22389 10100 22423
rect 10048 22380 10100 22389
rect 12532 22380 12584 22432
rect 16120 22380 16172 22432
rect 18236 22448 18288 22500
rect 20812 22448 20864 22500
rect 20996 22448 21048 22500
rect 18052 22380 18104 22432
rect 21180 22423 21232 22432
rect 21180 22389 21189 22423
rect 21189 22389 21223 22423
rect 21223 22389 21232 22423
rect 21180 22380 21232 22389
rect 21456 22448 21508 22500
rect 22192 22380 22244 22432
rect 23756 22584 23808 22636
rect 23112 22516 23164 22568
rect 23296 22516 23348 22568
rect 24400 22652 24452 22704
rect 24952 22652 25004 22704
rect 24860 22627 24912 22636
rect 24860 22593 24883 22627
rect 24883 22593 24912 22627
rect 24860 22584 24912 22593
rect 24492 22448 24544 22500
rect 24768 22380 24820 22432
rect 4124 22278 4176 22330
rect 4188 22278 4240 22330
rect 4252 22278 4304 22330
rect 4316 22278 4368 22330
rect 4380 22278 4432 22330
rect 10472 22278 10524 22330
rect 10536 22278 10588 22330
rect 10600 22278 10652 22330
rect 10664 22278 10716 22330
rect 10728 22278 10780 22330
rect 16820 22278 16872 22330
rect 16884 22278 16936 22330
rect 16948 22278 17000 22330
rect 17012 22278 17064 22330
rect 17076 22278 17128 22330
rect 23168 22278 23220 22330
rect 23232 22278 23284 22330
rect 23296 22278 23348 22330
rect 23360 22278 23412 22330
rect 23424 22278 23476 22330
rect 9312 22219 9364 22228
rect 9312 22185 9321 22219
rect 9321 22185 9355 22219
rect 9355 22185 9364 22219
rect 9312 22176 9364 22185
rect 13544 22176 13596 22228
rect 14004 22176 14056 22228
rect 16120 22219 16172 22228
rect 16120 22185 16129 22219
rect 16129 22185 16163 22219
rect 16163 22185 16172 22219
rect 16120 22176 16172 22185
rect 16488 22176 16540 22228
rect 18144 22176 18196 22228
rect 19800 22219 19852 22228
rect 19800 22185 19809 22219
rect 19809 22185 19843 22219
rect 19843 22185 19852 22219
rect 19800 22176 19852 22185
rect 19892 22219 19944 22228
rect 19892 22185 19901 22219
rect 19901 22185 19935 22219
rect 19935 22185 19944 22219
rect 19892 22176 19944 22185
rect 13728 22040 13780 22092
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 16212 22040 16264 22092
rect 10048 21972 10100 22024
rect 12348 21904 12400 21956
rect 11704 21836 11756 21888
rect 13636 21972 13688 22024
rect 14280 22015 14332 22024
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 14556 22015 14608 22024
rect 14556 21981 14565 22015
rect 14565 21981 14599 22015
rect 14599 21981 14608 22015
rect 14556 21972 14608 21981
rect 16672 21972 16724 22024
rect 14648 21904 14700 21956
rect 15384 21904 15436 21956
rect 16396 21947 16448 21956
rect 16396 21913 16423 21947
rect 16423 21913 16448 21947
rect 16396 21904 16448 21913
rect 22744 22176 22796 22228
rect 22928 22176 22980 22228
rect 24860 22176 24912 22228
rect 18144 22040 18196 22092
rect 21272 22083 21324 22092
rect 21272 22049 21281 22083
rect 21281 22049 21315 22083
rect 21315 22049 21324 22083
rect 21272 22040 21324 22049
rect 20996 22015 21048 22024
rect 20996 21981 21014 22015
rect 21014 21981 21048 22015
rect 20996 21972 21048 21981
rect 21640 21972 21692 22024
rect 24124 22040 24176 22092
rect 21180 21904 21232 21956
rect 21364 21947 21416 21956
rect 21364 21913 21373 21947
rect 21373 21913 21407 21947
rect 21407 21913 21416 21947
rect 21364 21904 21416 21913
rect 23664 21904 23716 21956
rect 17316 21836 17368 21888
rect 17776 21836 17828 21888
rect 18972 21879 19024 21888
rect 18972 21845 18981 21879
rect 18981 21845 19015 21879
rect 19015 21845 19024 21879
rect 18972 21836 19024 21845
rect 22928 21836 22980 21888
rect 24032 22015 24084 22024
rect 24032 21981 24041 22015
rect 24041 21981 24075 22015
rect 24075 21981 24084 22015
rect 25136 22040 25188 22092
rect 25780 22083 25832 22092
rect 25780 22049 25789 22083
rect 25789 22049 25823 22083
rect 25823 22049 25832 22083
rect 25780 22040 25832 22049
rect 24032 21972 24084 21981
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 7298 21734 7350 21786
rect 7362 21734 7414 21786
rect 7426 21734 7478 21786
rect 7490 21734 7542 21786
rect 7554 21734 7606 21786
rect 13646 21734 13698 21786
rect 13710 21734 13762 21786
rect 13774 21734 13826 21786
rect 13838 21734 13890 21786
rect 13902 21734 13954 21786
rect 19994 21734 20046 21786
rect 20058 21734 20110 21786
rect 20122 21734 20174 21786
rect 20186 21734 20238 21786
rect 20250 21734 20302 21786
rect 26342 21734 26394 21786
rect 26406 21734 26458 21786
rect 26470 21734 26522 21786
rect 26534 21734 26586 21786
rect 26598 21734 26650 21786
rect 8116 21632 8168 21684
rect 12348 21632 12400 21684
rect 14740 21632 14792 21684
rect 15384 21632 15436 21684
rect 15936 21632 15988 21684
rect 16028 21675 16080 21684
rect 16028 21641 16037 21675
rect 16037 21641 16071 21675
rect 16071 21641 16080 21675
rect 16028 21632 16080 21641
rect 17316 21675 17368 21684
rect 17316 21641 17325 21675
rect 17325 21641 17359 21675
rect 17359 21641 17368 21675
rect 17316 21632 17368 21641
rect 17408 21632 17460 21684
rect 9036 21496 9088 21548
rect 12164 21539 12216 21548
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 13084 21496 13136 21548
rect 15016 21564 15068 21616
rect 16580 21564 16632 21616
rect 17684 21675 17736 21684
rect 17684 21641 17693 21675
rect 17693 21641 17727 21675
rect 17727 21641 17736 21675
rect 17684 21632 17736 21641
rect 18052 21632 18104 21684
rect 18236 21632 18288 21684
rect 18972 21632 19024 21684
rect 21916 21632 21968 21684
rect 16212 21496 16264 21548
rect 16764 21539 16816 21548
rect 16764 21505 16773 21539
rect 16773 21505 16807 21539
rect 16807 21505 16816 21539
rect 16764 21496 16816 21505
rect 17408 21496 17460 21548
rect 17592 21496 17644 21548
rect 19892 21607 19944 21616
rect 19892 21573 19901 21607
rect 19901 21573 19935 21607
rect 19935 21573 19944 21607
rect 19892 21564 19944 21573
rect 22652 21632 22704 21684
rect 23664 21632 23716 21684
rect 24768 21632 24820 21684
rect 25320 21632 25372 21684
rect 17868 21496 17920 21548
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 18328 21539 18380 21548
rect 18328 21505 18337 21539
rect 18337 21505 18371 21539
rect 18371 21505 18380 21539
rect 18328 21496 18380 21505
rect 20628 21496 20680 21548
rect 20812 21496 20864 21548
rect 21456 21496 21508 21548
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 22100 21496 22152 21548
rect 7932 21471 7984 21480
rect 7932 21437 7941 21471
rect 7941 21437 7975 21471
rect 7975 21437 7984 21471
rect 7932 21428 7984 21437
rect 23664 21496 23716 21548
rect 23940 21539 23992 21548
rect 23940 21505 23949 21539
rect 23949 21505 23983 21539
rect 23983 21505 23992 21539
rect 23940 21496 23992 21505
rect 24124 21496 24176 21548
rect 25780 21539 25832 21548
rect 25780 21505 25789 21539
rect 25789 21505 25823 21539
rect 25823 21505 25832 21539
rect 25780 21496 25832 21505
rect 23572 21471 23624 21480
rect 23572 21437 23581 21471
rect 23581 21437 23615 21471
rect 23615 21437 23624 21471
rect 23572 21428 23624 21437
rect 25320 21471 25372 21480
rect 25320 21437 25329 21471
rect 25329 21437 25363 21471
rect 25363 21437 25372 21471
rect 25320 21428 25372 21437
rect 17224 21403 17276 21412
rect 17224 21369 17233 21403
rect 17233 21369 17267 21403
rect 17267 21369 17276 21403
rect 17224 21360 17276 21369
rect 18052 21360 18104 21412
rect 18604 21403 18656 21412
rect 18604 21369 18613 21403
rect 18613 21369 18647 21403
rect 18647 21369 18656 21403
rect 18604 21360 18656 21369
rect 22560 21360 22612 21412
rect 24032 21360 24084 21412
rect 9588 21292 9640 21344
rect 17500 21292 17552 21344
rect 22100 21292 22152 21344
rect 22836 21335 22888 21344
rect 22836 21301 22845 21335
rect 22845 21301 22879 21335
rect 22879 21301 22888 21335
rect 22836 21292 22888 21301
rect 24216 21292 24268 21344
rect 4124 21190 4176 21242
rect 4188 21190 4240 21242
rect 4252 21190 4304 21242
rect 4316 21190 4368 21242
rect 4380 21190 4432 21242
rect 10472 21190 10524 21242
rect 10536 21190 10588 21242
rect 10600 21190 10652 21242
rect 10664 21190 10716 21242
rect 10728 21190 10780 21242
rect 16820 21190 16872 21242
rect 16884 21190 16936 21242
rect 16948 21190 17000 21242
rect 17012 21190 17064 21242
rect 17076 21190 17128 21242
rect 23168 21190 23220 21242
rect 23232 21190 23284 21242
rect 23296 21190 23348 21242
rect 23360 21190 23412 21242
rect 23424 21190 23476 21242
rect 8576 20884 8628 20936
rect 8760 20927 8812 20936
rect 8760 20893 8769 20927
rect 8769 20893 8803 20927
rect 8803 20893 8812 20927
rect 8760 20884 8812 20893
rect 8392 20816 8444 20868
rect 9588 20884 9640 20936
rect 11336 20952 11388 21004
rect 14740 20952 14792 21004
rect 16488 21020 16540 21072
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 17040 21020 17092 21072
rect 17132 21020 17184 21072
rect 17868 21088 17920 21140
rect 18236 21088 18288 21140
rect 22008 21088 22060 21140
rect 23204 21088 23256 21140
rect 25320 21088 25372 21140
rect 11244 20816 11296 20868
rect 7840 20748 7892 20800
rect 8300 20791 8352 20800
rect 8300 20757 8309 20791
rect 8309 20757 8343 20791
rect 8343 20757 8352 20791
rect 8300 20748 8352 20757
rect 8668 20791 8720 20800
rect 8668 20757 8677 20791
rect 8677 20757 8711 20791
rect 8711 20757 8720 20791
rect 8668 20748 8720 20757
rect 8852 20748 8904 20800
rect 8944 20791 8996 20800
rect 8944 20757 8953 20791
rect 8953 20757 8987 20791
rect 8987 20757 8996 20791
rect 8944 20748 8996 20757
rect 9404 20748 9456 20800
rect 9680 20791 9732 20800
rect 9680 20757 9689 20791
rect 9689 20757 9723 20791
rect 9723 20757 9732 20791
rect 9680 20748 9732 20757
rect 12624 20816 12676 20868
rect 17040 20884 17092 20936
rect 18144 20884 18196 20936
rect 18604 20927 18656 20936
rect 18604 20893 18613 20927
rect 18613 20893 18647 20927
rect 18647 20893 18656 20927
rect 18604 20884 18656 20893
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 22744 20884 22796 20936
rect 22928 20927 22980 20936
rect 22928 20893 22937 20927
rect 22937 20893 22971 20927
rect 22971 20893 22980 20927
rect 22928 20884 22980 20893
rect 23204 20884 23256 20936
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 16948 20859 17000 20868
rect 16948 20825 16957 20859
rect 16957 20825 16991 20859
rect 16991 20825 17000 20859
rect 16948 20816 17000 20825
rect 12808 20791 12860 20800
rect 12808 20757 12817 20791
rect 12817 20757 12851 20791
rect 12851 20757 12860 20791
rect 12808 20748 12860 20757
rect 16580 20791 16632 20800
rect 16580 20757 16589 20791
rect 16589 20757 16623 20791
rect 16623 20757 16632 20791
rect 16580 20748 16632 20757
rect 16672 20748 16724 20800
rect 17040 20791 17092 20800
rect 17040 20757 17042 20791
rect 17042 20757 17076 20791
rect 17076 20757 17092 20791
rect 17040 20748 17092 20757
rect 22192 20859 22244 20868
rect 22192 20825 22201 20859
rect 22201 20825 22235 20859
rect 22235 20825 22244 20859
rect 23572 20884 23624 20936
rect 24216 20884 24268 20936
rect 22192 20816 22244 20825
rect 18236 20748 18288 20800
rect 18328 20791 18380 20800
rect 18328 20757 18337 20791
rect 18337 20757 18371 20791
rect 18371 20757 18380 20791
rect 18328 20748 18380 20757
rect 18420 20791 18472 20800
rect 18420 20757 18429 20791
rect 18429 20757 18463 20791
rect 18463 20757 18472 20791
rect 18420 20748 18472 20757
rect 22744 20748 22796 20800
rect 23756 20748 23808 20800
rect 7298 20646 7350 20698
rect 7362 20646 7414 20698
rect 7426 20646 7478 20698
rect 7490 20646 7542 20698
rect 7554 20646 7606 20698
rect 13646 20646 13698 20698
rect 13710 20646 13762 20698
rect 13774 20646 13826 20698
rect 13838 20646 13890 20698
rect 13902 20646 13954 20698
rect 19994 20646 20046 20698
rect 20058 20646 20110 20698
rect 20122 20646 20174 20698
rect 20186 20646 20238 20698
rect 20250 20646 20302 20698
rect 26342 20646 26394 20698
rect 26406 20646 26458 20698
rect 26470 20646 26522 20698
rect 26534 20646 26586 20698
rect 26598 20646 26650 20698
rect 8668 20544 8720 20596
rect 11336 20544 11388 20596
rect 11980 20587 12032 20596
rect 11980 20553 11989 20587
rect 11989 20553 12023 20587
rect 12023 20553 12032 20587
rect 11980 20544 12032 20553
rect 9036 20476 9088 20528
rect 11244 20476 11296 20528
rect 11612 20476 11664 20528
rect 15108 20544 15160 20596
rect 7564 20451 7616 20460
rect 7564 20417 7573 20451
rect 7573 20417 7607 20451
rect 7607 20417 7616 20451
rect 7564 20408 7616 20417
rect 7840 20408 7892 20460
rect 8024 20451 8076 20460
rect 8024 20417 8033 20451
rect 8033 20417 8067 20451
rect 8067 20417 8076 20451
rect 8024 20408 8076 20417
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 11888 20451 11940 20460
rect 11888 20417 11897 20451
rect 11897 20417 11931 20451
rect 11931 20417 11940 20451
rect 11888 20408 11940 20417
rect 9036 20340 9088 20392
rect 10048 20340 10100 20392
rect 12808 20476 12860 20528
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 16580 20476 16632 20528
rect 16764 20476 16816 20528
rect 13176 20408 13228 20417
rect 14096 20408 14148 20460
rect 14556 20408 14608 20460
rect 15292 20451 15344 20460
rect 15292 20417 15301 20451
rect 15301 20417 15335 20451
rect 15335 20417 15344 20451
rect 15292 20408 15344 20417
rect 17132 20408 17184 20460
rect 17408 20451 17460 20460
rect 17408 20417 17417 20451
rect 17417 20417 17451 20451
rect 17451 20417 17460 20451
rect 17408 20408 17460 20417
rect 18512 20587 18564 20596
rect 18512 20553 18521 20587
rect 18521 20553 18555 20587
rect 18555 20553 18564 20587
rect 18512 20544 18564 20553
rect 22744 20544 22796 20596
rect 23664 20544 23716 20596
rect 23940 20587 23992 20596
rect 23940 20553 23949 20587
rect 23949 20553 23983 20587
rect 23983 20553 23992 20587
rect 23940 20544 23992 20553
rect 24952 20587 25004 20596
rect 22100 20519 22152 20528
rect 22100 20485 22112 20519
rect 22112 20485 22152 20519
rect 22100 20476 22152 20485
rect 12808 20340 12860 20392
rect 18328 20408 18380 20460
rect 18604 20408 18656 20460
rect 19340 20408 19392 20460
rect 20536 20408 20588 20460
rect 20904 20408 20956 20460
rect 22560 20408 22612 20460
rect 23204 20408 23256 20460
rect 23480 20476 23532 20528
rect 13452 20272 13504 20324
rect 17776 20340 17828 20392
rect 8944 20204 8996 20256
rect 9404 20204 9456 20256
rect 13544 20247 13596 20256
rect 13544 20213 13553 20247
rect 13553 20213 13587 20247
rect 13587 20213 13596 20247
rect 13544 20204 13596 20213
rect 15936 20204 15988 20256
rect 17316 20204 17368 20256
rect 17684 20204 17736 20256
rect 20260 20204 20312 20256
rect 21640 20272 21692 20324
rect 20812 20247 20864 20256
rect 20812 20213 20821 20247
rect 20821 20213 20855 20247
rect 20855 20213 20864 20247
rect 20812 20204 20864 20213
rect 22928 20340 22980 20392
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 23664 20408 23716 20417
rect 24952 20553 24969 20587
rect 24969 20553 25004 20587
rect 24952 20544 25004 20553
rect 23572 20340 23624 20392
rect 23388 20272 23440 20324
rect 22192 20204 22244 20256
rect 23480 20204 23532 20256
rect 23664 20204 23716 20256
rect 24124 20204 24176 20256
rect 4124 20102 4176 20154
rect 4188 20102 4240 20154
rect 4252 20102 4304 20154
rect 4316 20102 4368 20154
rect 4380 20102 4432 20154
rect 10472 20102 10524 20154
rect 10536 20102 10588 20154
rect 10600 20102 10652 20154
rect 10664 20102 10716 20154
rect 10728 20102 10780 20154
rect 16820 20102 16872 20154
rect 16884 20102 16936 20154
rect 16948 20102 17000 20154
rect 17012 20102 17064 20154
rect 17076 20102 17128 20154
rect 23168 20102 23220 20154
rect 23232 20102 23284 20154
rect 23296 20102 23348 20154
rect 23360 20102 23412 20154
rect 23424 20102 23476 20154
rect 7564 20000 7616 20052
rect 7932 20000 7984 20052
rect 8760 20000 8812 20052
rect 9220 20000 9272 20052
rect 10048 20000 10100 20052
rect 12624 20000 12676 20052
rect 15292 20000 15344 20052
rect 16580 20000 16632 20052
rect 17408 20000 17460 20052
rect 18604 20000 18656 20052
rect 20812 20000 20864 20052
rect 20904 20000 20956 20052
rect 23572 20043 23624 20052
rect 23572 20009 23581 20043
rect 23581 20009 23615 20043
rect 23615 20009 23624 20043
rect 23572 20000 23624 20009
rect 7656 19796 7708 19848
rect 8024 19728 8076 19780
rect 7012 19660 7064 19712
rect 7932 19703 7984 19712
rect 7932 19669 7941 19703
rect 7941 19669 7975 19703
rect 7975 19669 7984 19703
rect 7932 19660 7984 19669
rect 8300 19864 8352 19916
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 8852 19796 8904 19848
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 12440 19932 12492 19984
rect 10508 19864 10560 19916
rect 14464 19864 14516 19916
rect 9312 19796 9364 19848
rect 9404 19839 9456 19848
rect 9404 19805 9413 19839
rect 9413 19805 9447 19839
rect 9447 19805 9456 19839
rect 9404 19796 9456 19805
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 9680 19796 9732 19848
rect 12808 19796 12860 19848
rect 14648 19839 14700 19848
rect 14648 19805 14657 19839
rect 14657 19805 14691 19839
rect 14691 19805 14700 19839
rect 14648 19796 14700 19805
rect 15108 19796 15160 19848
rect 16304 19796 16356 19848
rect 17684 19839 17736 19848
rect 17684 19805 17718 19839
rect 17718 19805 17736 19839
rect 17684 19796 17736 19805
rect 18972 19796 19024 19848
rect 22192 19907 22244 19916
rect 22192 19873 22201 19907
rect 22201 19873 22235 19907
rect 22235 19873 22244 19907
rect 22192 19864 22244 19873
rect 11244 19728 11296 19780
rect 11612 19728 11664 19780
rect 12624 19728 12676 19780
rect 16580 19771 16632 19780
rect 16580 19737 16589 19771
rect 16589 19737 16623 19771
rect 16623 19737 16632 19771
rect 16580 19728 16632 19737
rect 18420 19728 18472 19780
rect 12808 19703 12860 19712
rect 12808 19669 12817 19703
rect 12817 19669 12851 19703
rect 12851 19669 12860 19703
rect 12808 19660 12860 19669
rect 12900 19660 12952 19712
rect 14004 19660 14056 19712
rect 15200 19660 15252 19712
rect 16672 19660 16724 19712
rect 17500 19660 17552 19712
rect 17592 19660 17644 19712
rect 22744 19728 22796 19780
rect 20260 19660 20312 19712
rect 7298 19558 7350 19610
rect 7362 19558 7414 19610
rect 7426 19558 7478 19610
rect 7490 19558 7542 19610
rect 7554 19558 7606 19610
rect 13646 19558 13698 19610
rect 13710 19558 13762 19610
rect 13774 19558 13826 19610
rect 13838 19558 13890 19610
rect 13902 19558 13954 19610
rect 19994 19558 20046 19610
rect 20058 19558 20110 19610
rect 20122 19558 20174 19610
rect 20186 19558 20238 19610
rect 20250 19558 20302 19610
rect 26342 19558 26394 19610
rect 26406 19558 26458 19610
rect 26470 19558 26522 19610
rect 26534 19558 26586 19610
rect 26598 19558 26650 19610
rect 7656 19456 7708 19508
rect 7932 19456 7984 19508
rect 8760 19456 8812 19508
rect 8944 19456 8996 19508
rect 9128 19456 9180 19508
rect 9496 19456 9548 19508
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 7104 19320 7156 19372
rect 9404 19388 9456 19440
rect 9036 19320 9088 19372
rect 8392 19252 8444 19304
rect 9496 19320 9548 19372
rect 9956 19456 10008 19508
rect 11612 19388 11664 19440
rect 11888 19431 11940 19440
rect 11888 19397 11897 19431
rect 11897 19397 11931 19431
rect 11931 19397 11940 19431
rect 12532 19456 12584 19508
rect 13176 19456 13228 19508
rect 11888 19388 11940 19397
rect 10324 19320 10376 19372
rect 10508 19363 10560 19372
rect 10508 19329 10517 19363
rect 10517 19329 10551 19363
rect 10551 19329 10560 19363
rect 10508 19320 10560 19329
rect 11060 19320 11112 19372
rect 11152 19363 11204 19372
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11152 19320 11204 19329
rect 11336 19363 11388 19372
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 11428 19320 11480 19372
rect 9036 19184 9088 19236
rect 10876 19252 10928 19304
rect 11980 19363 12032 19372
rect 11980 19329 12015 19363
rect 12015 19329 12032 19363
rect 11980 19320 12032 19329
rect 12256 19363 12308 19372
rect 12256 19329 12265 19363
rect 12265 19329 12299 19363
rect 12299 19329 12308 19363
rect 12256 19320 12308 19329
rect 12348 19320 12400 19372
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 12624 19320 12676 19372
rect 14924 19320 14976 19372
rect 11888 19252 11940 19304
rect 12900 19252 12952 19304
rect 13360 19252 13412 19304
rect 15476 19252 15528 19304
rect 16488 19456 16540 19508
rect 18512 19456 18564 19508
rect 17224 19388 17276 19440
rect 16580 19252 16632 19304
rect 940 19116 992 19168
rect 6552 19159 6604 19168
rect 6552 19125 6561 19159
rect 6561 19125 6595 19159
rect 6595 19125 6604 19159
rect 6552 19116 6604 19125
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 8576 19116 8628 19168
rect 10232 19184 10284 19236
rect 10416 19227 10468 19236
rect 10416 19193 10425 19227
rect 10425 19193 10459 19227
rect 10459 19193 10468 19227
rect 10416 19184 10468 19193
rect 11336 19184 11388 19236
rect 12348 19184 12400 19236
rect 18328 19320 18380 19372
rect 18420 19320 18472 19372
rect 18972 19388 19024 19440
rect 20904 19388 20956 19440
rect 21640 19456 21692 19508
rect 22744 19499 22796 19508
rect 22744 19465 22753 19499
rect 22753 19465 22787 19499
rect 22787 19465 22796 19499
rect 22744 19456 22796 19465
rect 19340 19295 19392 19304
rect 19340 19261 19349 19295
rect 19349 19261 19383 19295
rect 19383 19261 19392 19295
rect 22192 19320 22244 19372
rect 23664 19320 23716 19372
rect 19340 19252 19392 19261
rect 22836 19252 22888 19304
rect 18328 19184 18380 19236
rect 9588 19116 9640 19168
rect 12072 19116 12124 19168
rect 12164 19116 12216 19168
rect 13636 19116 13688 19168
rect 14096 19116 14148 19168
rect 15200 19116 15252 19168
rect 17500 19116 17552 19168
rect 19800 19184 19852 19236
rect 4124 19014 4176 19066
rect 4188 19014 4240 19066
rect 4252 19014 4304 19066
rect 4316 19014 4368 19066
rect 4380 19014 4432 19066
rect 10472 19014 10524 19066
rect 10536 19014 10588 19066
rect 10600 19014 10652 19066
rect 10664 19014 10716 19066
rect 10728 19014 10780 19066
rect 16820 19014 16872 19066
rect 16884 19014 16936 19066
rect 16948 19014 17000 19066
rect 17012 19014 17064 19066
rect 17076 19014 17128 19066
rect 23168 19014 23220 19066
rect 23232 19014 23284 19066
rect 23296 19014 23348 19066
rect 23360 19014 23412 19066
rect 23424 19014 23476 19066
rect 7104 18912 7156 18964
rect 8392 18912 8444 18964
rect 6368 18776 6420 18828
rect 8300 18776 8352 18828
rect 6920 18640 6972 18692
rect 8668 18708 8720 18760
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 9496 18912 9548 18964
rect 11152 18912 11204 18964
rect 11704 18844 11756 18896
rect 11888 18844 11940 18896
rect 12440 18912 12492 18964
rect 13360 18912 13412 18964
rect 13544 18912 13596 18964
rect 14648 18912 14700 18964
rect 18420 18955 18472 18964
rect 18420 18921 18429 18955
rect 18429 18921 18463 18955
rect 18463 18921 18472 18955
rect 18420 18912 18472 18921
rect 12716 18844 12768 18896
rect 12624 18776 12676 18828
rect 14280 18844 14332 18896
rect 19340 18844 19392 18896
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 10416 18751 10468 18760
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 11152 18708 11204 18760
rect 8208 18640 8260 18692
rect 9864 18640 9916 18692
rect 11244 18683 11296 18692
rect 11244 18649 11253 18683
rect 11253 18649 11287 18683
rect 11287 18649 11296 18683
rect 11244 18640 11296 18649
rect 7012 18572 7064 18624
rect 8116 18572 8168 18624
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 12348 18751 12400 18760
rect 12348 18717 12357 18751
rect 12357 18717 12391 18751
rect 12391 18717 12400 18751
rect 12348 18708 12400 18717
rect 13176 18751 13228 18760
rect 13176 18717 13185 18751
rect 13185 18717 13219 18751
rect 13219 18717 13228 18751
rect 13176 18708 13228 18717
rect 13544 18751 13596 18760
rect 13544 18717 13553 18751
rect 13553 18717 13587 18751
rect 13587 18717 13596 18751
rect 13544 18708 13596 18717
rect 15936 18819 15988 18828
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 12164 18683 12216 18692
rect 12164 18649 12173 18683
rect 12173 18649 12207 18683
rect 12207 18649 12216 18683
rect 12164 18640 12216 18649
rect 13084 18640 13136 18692
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 14648 18708 14700 18760
rect 16580 18708 16632 18760
rect 17316 18751 17368 18760
rect 17316 18717 17350 18751
rect 17350 18717 17368 18751
rect 17316 18708 17368 18717
rect 20352 18708 20404 18760
rect 20720 18708 20772 18760
rect 22836 18751 22888 18760
rect 22836 18717 22845 18751
rect 22845 18717 22879 18751
rect 22879 18717 22888 18751
rect 22836 18708 22888 18717
rect 13452 18572 13504 18624
rect 14188 18640 14240 18692
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 14924 18572 14976 18624
rect 15660 18640 15712 18692
rect 17500 18640 17552 18692
rect 19708 18572 19760 18624
rect 23296 18572 23348 18624
rect 7298 18470 7350 18522
rect 7362 18470 7414 18522
rect 7426 18470 7478 18522
rect 7490 18470 7542 18522
rect 7554 18470 7606 18522
rect 13646 18470 13698 18522
rect 13710 18470 13762 18522
rect 13774 18470 13826 18522
rect 13838 18470 13890 18522
rect 13902 18470 13954 18522
rect 19994 18470 20046 18522
rect 20058 18470 20110 18522
rect 20122 18470 20174 18522
rect 20186 18470 20238 18522
rect 20250 18470 20302 18522
rect 26342 18470 26394 18522
rect 26406 18470 26458 18522
rect 26470 18470 26522 18522
rect 26534 18470 26586 18522
rect 26598 18470 26650 18522
rect 1768 18368 1820 18420
rect 8116 18411 8168 18420
rect 8116 18377 8125 18411
rect 8125 18377 8159 18411
rect 8159 18377 8168 18411
rect 8116 18368 8168 18377
rect 8300 18368 8352 18420
rect 6552 18300 6604 18352
rect 7932 18232 7984 18284
rect 6368 18207 6420 18216
rect 6368 18173 6377 18207
rect 6377 18173 6411 18207
rect 6411 18173 6420 18207
rect 6368 18164 6420 18173
rect 7104 18028 7156 18080
rect 8576 18300 8628 18352
rect 11244 18368 11296 18420
rect 11428 18368 11480 18420
rect 14096 18368 14148 18420
rect 14372 18368 14424 18420
rect 15476 18368 15528 18420
rect 19708 18368 19760 18420
rect 9036 18300 9088 18352
rect 9956 18232 10008 18284
rect 10048 18232 10100 18284
rect 8944 18164 8996 18216
rect 9404 18164 9456 18216
rect 10324 18232 10376 18284
rect 10692 18232 10744 18284
rect 11060 18232 11112 18284
rect 11336 18275 11388 18284
rect 11336 18241 11345 18275
rect 11345 18241 11379 18275
rect 11379 18241 11388 18275
rect 11336 18232 11388 18241
rect 12072 18275 12124 18284
rect 12072 18241 12081 18275
rect 12081 18241 12115 18275
rect 12115 18241 12124 18275
rect 12072 18232 12124 18241
rect 12440 18300 12492 18352
rect 10968 18164 11020 18216
rect 10416 18139 10468 18148
rect 10416 18105 10425 18139
rect 10425 18105 10459 18139
rect 10459 18105 10468 18139
rect 10416 18096 10468 18105
rect 11336 18096 11388 18148
rect 12072 18096 12124 18148
rect 11060 18071 11112 18080
rect 11060 18037 11069 18071
rect 11069 18037 11103 18071
rect 11103 18037 11112 18071
rect 11060 18028 11112 18037
rect 11520 18071 11572 18080
rect 11520 18037 11529 18071
rect 11529 18037 11563 18071
rect 11563 18037 11572 18071
rect 11520 18028 11572 18037
rect 12256 18232 12308 18284
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 13452 18232 13504 18284
rect 13544 18232 13596 18284
rect 14004 18232 14056 18284
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 18972 18232 19024 18284
rect 20536 18232 20588 18284
rect 12256 18096 12308 18148
rect 22192 18232 22244 18284
rect 22744 18275 22796 18284
rect 22744 18241 22753 18275
rect 22753 18241 22787 18275
rect 22787 18241 22796 18275
rect 22744 18232 22796 18241
rect 23296 18300 23348 18352
rect 22008 18164 22060 18216
rect 22928 18164 22980 18216
rect 23388 18164 23440 18216
rect 25136 18207 25188 18216
rect 25136 18173 25145 18207
rect 25145 18173 25179 18207
rect 25179 18173 25188 18207
rect 25136 18164 25188 18173
rect 13176 18028 13228 18080
rect 13544 18071 13596 18080
rect 13544 18037 13553 18071
rect 13553 18037 13587 18071
rect 13587 18037 13596 18071
rect 13544 18028 13596 18037
rect 14464 18028 14516 18080
rect 20904 18071 20956 18080
rect 20904 18037 20913 18071
rect 20913 18037 20947 18071
rect 20947 18037 20956 18071
rect 20904 18028 20956 18037
rect 22560 18071 22612 18080
rect 22560 18037 22569 18071
rect 22569 18037 22603 18071
rect 22603 18037 22612 18071
rect 22560 18028 22612 18037
rect 24124 18028 24176 18080
rect 4124 17926 4176 17978
rect 4188 17926 4240 17978
rect 4252 17926 4304 17978
rect 4316 17926 4368 17978
rect 4380 17926 4432 17978
rect 10472 17926 10524 17978
rect 10536 17926 10588 17978
rect 10600 17926 10652 17978
rect 10664 17926 10716 17978
rect 10728 17926 10780 17978
rect 16820 17926 16872 17978
rect 16884 17926 16936 17978
rect 16948 17926 17000 17978
rect 17012 17926 17064 17978
rect 17076 17926 17128 17978
rect 23168 17926 23220 17978
rect 23232 17926 23284 17978
rect 23296 17926 23348 17978
rect 23360 17926 23412 17978
rect 23424 17926 23476 17978
rect 8208 17824 8260 17876
rect 8392 17867 8444 17876
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 8576 17824 8628 17876
rect 9128 17867 9180 17876
rect 9128 17833 9137 17867
rect 9137 17833 9171 17867
rect 9171 17833 9180 17867
rect 9128 17824 9180 17833
rect 6000 17688 6052 17740
rect 11980 17824 12032 17876
rect 5816 17620 5868 17672
rect 8484 17620 8536 17672
rect 9956 17688 10008 17740
rect 11060 17688 11112 17740
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 4620 17484 4672 17536
rect 6644 17484 6696 17536
rect 7932 17484 7984 17536
rect 9772 17620 9824 17672
rect 12348 17867 12400 17876
rect 12348 17833 12357 17867
rect 12357 17833 12391 17867
rect 12391 17833 12400 17867
rect 12348 17824 12400 17833
rect 22100 17824 22152 17876
rect 22836 17824 22888 17876
rect 12532 17799 12584 17808
rect 12532 17765 12541 17799
rect 12541 17765 12575 17799
rect 12575 17765 12584 17799
rect 12532 17756 12584 17765
rect 9312 17484 9364 17536
rect 10048 17484 10100 17536
rect 11152 17552 11204 17604
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 11520 17620 11572 17672
rect 12072 17663 12124 17672
rect 12072 17629 12081 17663
rect 12081 17629 12115 17663
rect 12115 17629 12124 17663
rect 12072 17620 12124 17629
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 14556 17620 14608 17629
rect 15660 17620 15712 17672
rect 18604 17620 18656 17672
rect 18788 17620 18840 17672
rect 18880 17620 18932 17672
rect 20536 17620 20588 17672
rect 21088 17688 21140 17740
rect 22192 17688 22244 17740
rect 24860 17824 24912 17876
rect 23572 17756 23624 17808
rect 11612 17552 11664 17604
rect 12716 17595 12768 17604
rect 12716 17561 12725 17595
rect 12725 17561 12759 17595
rect 12759 17561 12768 17595
rect 12716 17552 12768 17561
rect 11428 17484 11480 17536
rect 12256 17484 12308 17536
rect 14832 17527 14884 17536
rect 14832 17493 14841 17527
rect 14841 17493 14875 17527
rect 14875 17493 14884 17527
rect 14832 17484 14884 17493
rect 17224 17484 17276 17536
rect 18420 17484 18472 17536
rect 19064 17484 19116 17536
rect 22100 17552 22152 17604
rect 22376 17620 22428 17672
rect 22928 17663 22980 17672
rect 22928 17629 22937 17663
rect 22937 17629 22971 17663
rect 22971 17629 22980 17663
rect 22928 17620 22980 17629
rect 24124 17688 24176 17740
rect 20996 17484 21048 17536
rect 21088 17484 21140 17536
rect 22836 17552 22888 17604
rect 22284 17484 22336 17536
rect 23020 17484 23072 17536
rect 23664 17527 23716 17536
rect 23664 17493 23673 17527
rect 23673 17493 23707 17527
rect 23707 17493 23716 17527
rect 23664 17484 23716 17493
rect 23756 17484 23808 17536
rect 24032 17484 24084 17536
rect 24952 17552 25004 17604
rect 25044 17484 25096 17536
rect 26148 17527 26200 17536
rect 26148 17493 26157 17527
rect 26157 17493 26191 17527
rect 26191 17493 26200 17527
rect 26148 17484 26200 17493
rect 7298 17382 7350 17434
rect 7362 17382 7414 17434
rect 7426 17382 7478 17434
rect 7490 17382 7542 17434
rect 7554 17382 7606 17434
rect 13646 17382 13698 17434
rect 13710 17382 13762 17434
rect 13774 17382 13826 17434
rect 13838 17382 13890 17434
rect 13902 17382 13954 17434
rect 19994 17382 20046 17434
rect 20058 17382 20110 17434
rect 20122 17382 20174 17434
rect 20186 17382 20238 17434
rect 20250 17382 20302 17434
rect 26342 17382 26394 17434
rect 26406 17382 26458 17434
rect 26470 17382 26522 17434
rect 26534 17382 26586 17434
rect 26598 17382 26650 17434
rect 11612 17323 11664 17332
rect 11612 17289 11621 17323
rect 11621 17289 11655 17323
rect 11655 17289 11664 17323
rect 11612 17280 11664 17289
rect 12716 17280 12768 17332
rect 14556 17280 14608 17332
rect 17224 17280 17276 17332
rect 18420 17323 18472 17332
rect 18420 17289 18429 17323
rect 18429 17289 18463 17323
rect 18463 17289 18472 17323
rect 18420 17280 18472 17289
rect 18880 17323 18932 17332
rect 18880 17289 18889 17323
rect 18889 17289 18923 17323
rect 18923 17289 18932 17323
rect 18880 17280 18932 17289
rect 19064 17280 19116 17332
rect 3976 17144 4028 17196
rect 6276 17144 6328 17196
rect 9864 17144 9916 17196
rect 2412 17119 2464 17128
rect 2412 17085 2421 17119
rect 2421 17085 2455 17119
rect 2455 17085 2464 17119
rect 2412 17076 2464 17085
rect 3240 17076 3292 17128
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 5540 17076 5592 17128
rect 6460 17119 6512 17128
rect 6460 17085 6469 17119
rect 6469 17085 6503 17119
rect 6503 17085 6512 17119
rect 6460 17076 6512 17085
rect 10232 17076 10284 17128
rect 10968 17076 11020 17128
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 12900 17144 12952 17196
rect 12992 17144 13044 17196
rect 14280 17212 14332 17264
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 22284 17280 22336 17332
rect 22836 17280 22888 17332
rect 24216 17280 24268 17332
rect 25044 17323 25096 17332
rect 25044 17289 25053 17323
rect 25053 17289 25087 17323
rect 25087 17289 25096 17323
rect 25044 17280 25096 17289
rect 20536 17212 20588 17264
rect 22468 17212 22520 17264
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 12164 17008 12216 17060
rect 14556 17008 14608 17060
rect 4528 16940 4580 16992
rect 7564 16940 7616 16992
rect 11428 16940 11480 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 15292 17076 15344 17128
rect 16580 17076 16632 17128
rect 18696 17144 18748 17196
rect 20904 17144 20956 17196
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 14832 17008 14884 17060
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 19248 17076 19300 17128
rect 20628 17076 20680 17128
rect 21180 17076 21232 17128
rect 22008 17076 22060 17128
rect 22284 17187 22336 17196
rect 22284 17153 22293 17187
rect 22293 17153 22327 17187
rect 22327 17153 22336 17187
rect 22284 17144 22336 17153
rect 22652 17187 22704 17196
rect 22652 17153 22661 17187
rect 22661 17153 22695 17187
rect 22695 17153 22704 17187
rect 22652 17144 22704 17153
rect 23296 17187 23348 17196
rect 23296 17153 23305 17187
rect 23305 17153 23339 17187
rect 23339 17153 23348 17187
rect 23296 17144 23348 17153
rect 24860 17144 24912 17196
rect 25320 17144 25372 17196
rect 26148 17144 26200 17196
rect 22744 17076 22796 17128
rect 22928 17076 22980 17128
rect 22652 17008 22704 17060
rect 23572 17119 23624 17128
rect 23572 17085 23581 17119
rect 23581 17085 23615 17119
rect 23615 17085 23624 17119
rect 23572 17076 23624 17085
rect 15752 16940 15804 16992
rect 18696 16983 18748 16992
rect 18696 16949 18705 16983
rect 18705 16949 18739 16983
rect 18739 16949 18748 16983
rect 18696 16940 18748 16949
rect 18880 16940 18932 16992
rect 19340 16940 19392 16992
rect 20812 16983 20864 16992
rect 20812 16949 20821 16983
rect 20821 16949 20855 16983
rect 20855 16949 20864 16983
rect 20812 16940 20864 16949
rect 22376 16940 22428 16992
rect 22928 16983 22980 16992
rect 22928 16949 22937 16983
rect 22937 16949 22971 16983
rect 22971 16949 22980 16983
rect 22928 16940 22980 16949
rect 24216 16940 24268 16992
rect 25964 16983 26016 16992
rect 25964 16949 25973 16983
rect 25973 16949 26007 16983
rect 26007 16949 26016 16983
rect 25964 16940 26016 16949
rect 4124 16838 4176 16890
rect 4188 16838 4240 16890
rect 4252 16838 4304 16890
rect 4316 16838 4368 16890
rect 4380 16838 4432 16890
rect 10472 16838 10524 16890
rect 10536 16838 10588 16890
rect 10600 16838 10652 16890
rect 10664 16838 10716 16890
rect 10728 16838 10780 16890
rect 16820 16838 16872 16890
rect 16884 16838 16936 16890
rect 16948 16838 17000 16890
rect 17012 16838 17064 16890
rect 17076 16838 17128 16890
rect 23168 16838 23220 16890
rect 23232 16838 23284 16890
rect 23296 16838 23348 16890
rect 23360 16838 23412 16890
rect 23424 16838 23476 16890
rect 2412 16736 2464 16788
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 7564 16736 7616 16788
rect 11428 16736 11480 16788
rect 12072 16668 12124 16720
rect 6368 16600 6420 16652
rect 7012 16600 7064 16652
rect 10324 16600 10376 16652
rect 11244 16600 11296 16652
rect 14372 16736 14424 16788
rect 14556 16736 14608 16788
rect 20444 16736 20496 16788
rect 20720 16736 20772 16788
rect 21640 16779 21692 16788
rect 21640 16745 21649 16779
rect 21649 16745 21683 16779
rect 21683 16745 21692 16779
rect 21640 16736 21692 16745
rect 23572 16736 23624 16788
rect 4436 16575 4488 16584
rect 4436 16541 4445 16575
rect 4445 16541 4479 16575
rect 4479 16541 4488 16575
rect 4436 16532 4488 16541
rect 4528 16532 4580 16584
rect 6920 16532 6972 16584
rect 4252 16464 4304 16516
rect 6368 16464 6420 16516
rect 6000 16396 6052 16448
rect 10784 16464 10836 16516
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 8944 16396 8996 16405
rect 10140 16396 10192 16448
rect 10968 16396 11020 16448
rect 12532 16575 12584 16584
rect 12532 16541 12541 16575
rect 12541 16541 12575 16575
rect 12575 16541 12584 16575
rect 18604 16668 18656 16720
rect 12532 16532 12584 16541
rect 12624 16396 12676 16448
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 13268 16439 13320 16448
rect 13268 16405 13277 16439
rect 13277 16405 13311 16439
rect 13311 16405 13320 16439
rect 13268 16396 13320 16405
rect 13544 16396 13596 16448
rect 14832 16464 14884 16516
rect 16580 16600 16632 16652
rect 18696 16600 18748 16652
rect 18328 16532 18380 16584
rect 18788 16532 18840 16584
rect 19340 16600 19392 16652
rect 20812 16668 20864 16720
rect 21548 16668 21600 16720
rect 22928 16668 22980 16720
rect 24952 16736 25004 16788
rect 19248 16575 19300 16584
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19248 16532 19300 16541
rect 19800 16532 19852 16584
rect 19892 16532 19944 16584
rect 21732 16600 21784 16652
rect 21916 16600 21968 16652
rect 22560 16600 22612 16652
rect 22652 16643 22704 16652
rect 22652 16609 22661 16643
rect 22661 16609 22695 16643
rect 22695 16609 22704 16643
rect 22652 16600 22704 16609
rect 22836 16600 22888 16652
rect 20904 16532 20956 16584
rect 20996 16532 21048 16584
rect 17500 16464 17552 16516
rect 22008 16575 22060 16584
rect 22008 16541 22017 16575
rect 22017 16541 22051 16575
rect 22051 16541 22060 16575
rect 22008 16532 22060 16541
rect 23940 16600 23992 16652
rect 25504 16668 25556 16720
rect 25044 16643 25096 16652
rect 25044 16609 25053 16643
rect 25053 16609 25087 16643
rect 25087 16609 25096 16643
rect 25044 16600 25096 16609
rect 25964 16600 26016 16652
rect 19524 16396 19576 16448
rect 20904 16439 20956 16448
rect 20904 16405 20913 16439
rect 20913 16405 20947 16439
rect 20947 16405 20956 16439
rect 20904 16396 20956 16405
rect 22376 16464 22428 16516
rect 22744 16464 22796 16516
rect 22928 16464 22980 16516
rect 23388 16507 23440 16516
rect 23388 16473 23397 16507
rect 23397 16473 23431 16507
rect 23431 16473 23440 16507
rect 23388 16464 23440 16473
rect 23480 16507 23532 16516
rect 23480 16473 23489 16507
rect 23489 16473 23523 16507
rect 23523 16473 23532 16507
rect 23480 16464 23532 16473
rect 23572 16507 23624 16516
rect 23572 16473 23607 16507
rect 23607 16473 23624 16507
rect 23572 16464 23624 16473
rect 23112 16396 23164 16448
rect 24032 16507 24084 16516
rect 24032 16473 24041 16507
rect 24041 16473 24075 16507
rect 24075 16473 24084 16507
rect 24032 16464 24084 16473
rect 25412 16507 25464 16516
rect 25412 16473 25421 16507
rect 25421 16473 25455 16507
rect 25455 16473 25464 16507
rect 25412 16464 25464 16473
rect 25504 16507 25556 16516
rect 25504 16473 25514 16507
rect 25514 16473 25548 16507
rect 25548 16473 25556 16507
rect 25504 16464 25556 16473
rect 25688 16464 25740 16516
rect 25872 16575 25924 16584
rect 25872 16541 25881 16575
rect 25881 16541 25915 16575
rect 25915 16541 25924 16575
rect 25872 16532 25924 16541
rect 7298 16294 7350 16346
rect 7362 16294 7414 16346
rect 7426 16294 7478 16346
rect 7490 16294 7542 16346
rect 7554 16294 7606 16346
rect 13646 16294 13698 16346
rect 13710 16294 13762 16346
rect 13774 16294 13826 16346
rect 13838 16294 13890 16346
rect 13902 16294 13954 16346
rect 19994 16294 20046 16346
rect 20058 16294 20110 16346
rect 20122 16294 20174 16346
rect 20186 16294 20238 16346
rect 20250 16294 20302 16346
rect 26342 16294 26394 16346
rect 26406 16294 26458 16346
rect 26470 16294 26522 16346
rect 26534 16294 26586 16346
rect 26598 16294 26650 16346
rect 3976 16192 4028 16244
rect 3148 16124 3200 16176
rect 5816 16192 5868 16244
rect 6460 16192 6512 16244
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 6276 16124 6328 16176
rect 6920 16124 6972 16176
rect 7012 16124 7064 16176
rect 8944 16192 8996 16244
rect 10232 16192 10284 16244
rect 11244 16192 11296 16244
rect 12900 16192 12952 16244
rect 13452 16192 13504 16244
rect 7472 16056 7524 16108
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 3424 15988 3476 16040
rect 1676 15852 1728 15904
rect 4252 15988 4304 16040
rect 6460 15988 6512 16040
rect 10048 16056 10100 16108
rect 9772 15988 9824 16040
rect 12716 16124 12768 16176
rect 14832 16124 14884 16176
rect 12072 16056 12124 16108
rect 15476 16056 15528 16108
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 13544 16031 13596 16040
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 13820 16031 13872 16040
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 18604 16192 18656 16244
rect 19248 16192 19300 16244
rect 17500 16124 17552 16176
rect 19800 16235 19852 16244
rect 19800 16201 19809 16235
rect 19809 16201 19843 16235
rect 19843 16201 19852 16235
rect 19800 16192 19852 16201
rect 19892 16192 19944 16244
rect 20904 16192 20956 16244
rect 22376 16192 22428 16244
rect 23020 16192 23072 16244
rect 23388 16192 23440 16244
rect 24032 16192 24084 16244
rect 16396 16099 16448 16108
rect 16396 16065 16405 16099
rect 16405 16065 16439 16099
rect 16439 16065 16448 16099
rect 16396 16056 16448 16065
rect 16580 16056 16632 16108
rect 18420 16056 18472 16108
rect 19524 16056 19576 16108
rect 23480 16124 23532 16176
rect 23756 16124 23808 16176
rect 9680 15920 9732 15972
rect 5540 15852 5592 15904
rect 11980 15895 12032 15904
rect 11980 15861 11989 15895
rect 11989 15861 12023 15895
rect 12023 15861 12032 15895
rect 11980 15852 12032 15861
rect 13912 15852 13964 15904
rect 14004 15852 14056 15904
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 22008 15988 22060 16040
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 24952 16192 25004 16244
rect 25412 16192 25464 16244
rect 25504 16192 25556 16244
rect 25136 16124 25188 16176
rect 25596 16124 25648 16176
rect 25044 16056 25096 16108
rect 25412 16099 25464 16108
rect 25412 16065 25421 16099
rect 25421 16065 25455 16099
rect 25455 16065 25464 16099
rect 25412 16056 25464 16065
rect 16212 15963 16264 15972
rect 16212 15929 16221 15963
rect 16221 15929 16255 15963
rect 16255 15929 16264 15963
rect 16212 15920 16264 15929
rect 16672 15920 16724 15972
rect 22928 15920 22980 15972
rect 15292 15852 15344 15861
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 24584 15852 24636 15904
rect 25320 15852 25372 15904
rect 25412 15852 25464 15904
rect 25872 15920 25924 15972
rect 25780 15895 25832 15904
rect 25780 15861 25789 15895
rect 25789 15861 25823 15895
rect 25823 15861 25832 15895
rect 25780 15852 25832 15861
rect 4124 15750 4176 15802
rect 4188 15750 4240 15802
rect 4252 15750 4304 15802
rect 4316 15750 4368 15802
rect 4380 15750 4432 15802
rect 10472 15750 10524 15802
rect 10536 15750 10588 15802
rect 10600 15750 10652 15802
rect 10664 15750 10716 15802
rect 10728 15750 10780 15802
rect 16820 15750 16872 15802
rect 16884 15750 16936 15802
rect 16948 15750 17000 15802
rect 17012 15750 17064 15802
rect 17076 15750 17128 15802
rect 23168 15750 23220 15802
rect 23232 15750 23284 15802
rect 23296 15750 23348 15802
rect 23360 15750 23412 15802
rect 23424 15750 23476 15802
rect 1860 15648 1912 15700
rect 3148 15648 3200 15700
rect 5724 15648 5776 15700
rect 7748 15648 7800 15700
rect 10140 15648 10192 15700
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 5540 15512 5592 15564
rect 6736 15555 6788 15564
rect 6736 15521 6745 15555
rect 6745 15521 6779 15555
rect 6779 15521 6788 15555
rect 6736 15512 6788 15521
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 11244 15512 11296 15564
rect 4896 15444 4948 15496
rect 6368 15487 6420 15496
rect 6368 15453 6377 15487
rect 6377 15453 6411 15487
rect 6411 15453 6420 15487
rect 6368 15444 6420 15453
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 12900 15648 12952 15700
rect 13268 15648 13320 15700
rect 13544 15648 13596 15700
rect 13820 15648 13872 15700
rect 13912 15648 13964 15700
rect 14556 15648 14608 15700
rect 15016 15648 15068 15700
rect 16672 15648 16724 15700
rect 18512 15648 18564 15700
rect 21088 15648 21140 15700
rect 12624 15444 12676 15496
rect 14832 15512 14884 15564
rect 15568 15512 15620 15564
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 14004 15444 14056 15496
rect 18328 15512 18380 15564
rect 4896 15351 4948 15360
rect 4896 15317 4905 15351
rect 4905 15317 4939 15351
rect 4939 15317 4948 15351
rect 4896 15308 4948 15317
rect 7472 15376 7524 15428
rect 10140 15308 10192 15360
rect 10324 15351 10376 15360
rect 10324 15317 10333 15351
rect 10333 15317 10367 15351
rect 10367 15317 10376 15351
rect 10324 15308 10376 15317
rect 10968 15376 11020 15428
rect 12256 15351 12308 15360
rect 12256 15317 12265 15351
rect 12265 15317 12299 15351
rect 12299 15317 12308 15351
rect 12256 15308 12308 15317
rect 14556 15308 14608 15360
rect 14832 15376 14884 15428
rect 18420 15376 18472 15428
rect 18604 15487 18656 15496
rect 18604 15453 18613 15487
rect 18613 15453 18647 15487
rect 18647 15453 18656 15487
rect 18604 15444 18656 15453
rect 19892 15512 19944 15564
rect 19248 15487 19300 15496
rect 19248 15453 19257 15487
rect 19257 15453 19291 15487
rect 19291 15453 19300 15487
rect 19248 15444 19300 15453
rect 20904 15512 20956 15564
rect 21180 15487 21232 15496
rect 21180 15453 21189 15487
rect 21189 15453 21223 15487
rect 21223 15453 21232 15487
rect 21180 15444 21232 15453
rect 22376 15487 22428 15496
rect 22376 15453 22385 15487
rect 22385 15453 22419 15487
rect 22419 15453 22428 15487
rect 22376 15444 22428 15453
rect 23112 15512 23164 15564
rect 24584 15512 24636 15564
rect 23940 15444 23992 15496
rect 25780 15512 25832 15564
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 24952 15444 25004 15453
rect 26056 15487 26108 15496
rect 26056 15453 26065 15487
rect 26065 15453 26099 15487
rect 26099 15453 26108 15487
rect 26056 15444 26108 15453
rect 19616 15376 19668 15428
rect 24216 15376 24268 15428
rect 15200 15308 15252 15360
rect 18788 15351 18840 15360
rect 18788 15317 18797 15351
rect 18797 15317 18831 15351
rect 18831 15317 18840 15351
rect 18788 15308 18840 15317
rect 21088 15308 21140 15360
rect 24492 15351 24544 15360
rect 24492 15317 24501 15351
rect 24501 15317 24535 15351
rect 24535 15317 24544 15351
rect 24492 15308 24544 15317
rect 7298 15206 7350 15258
rect 7362 15206 7414 15258
rect 7426 15206 7478 15258
rect 7490 15206 7542 15258
rect 7554 15206 7606 15258
rect 13646 15206 13698 15258
rect 13710 15206 13762 15258
rect 13774 15206 13826 15258
rect 13838 15206 13890 15258
rect 13902 15206 13954 15258
rect 19994 15206 20046 15258
rect 20058 15206 20110 15258
rect 20122 15206 20174 15258
rect 20186 15206 20238 15258
rect 20250 15206 20302 15258
rect 26342 15206 26394 15258
rect 26406 15206 26458 15258
rect 26470 15206 26522 15258
rect 26534 15206 26586 15258
rect 26598 15206 26650 15258
rect 6460 15104 6512 15156
rect 3148 15036 3200 15088
rect 9680 15104 9732 15156
rect 10324 15104 10376 15156
rect 10416 15147 10468 15156
rect 10416 15113 10425 15147
rect 10425 15113 10459 15147
rect 10459 15113 10468 15147
rect 10416 15104 10468 15113
rect 10876 15147 10928 15156
rect 10876 15113 10885 15147
rect 10885 15113 10919 15147
rect 10919 15113 10928 15147
rect 10876 15104 10928 15113
rect 6736 14968 6788 15020
rect 2412 14900 2464 14952
rect 3240 14900 3292 14952
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 8760 14832 8812 14884
rect 10048 14968 10100 15020
rect 10140 14968 10192 15020
rect 12256 15104 12308 15156
rect 1676 14764 1728 14816
rect 8668 14764 8720 14816
rect 9588 14900 9640 14952
rect 11520 14900 11572 14952
rect 13452 15036 13504 15088
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 17500 15104 17552 15156
rect 19248 15104 19300 15156
rect 17960 15036 18012 15088
rect 19340 15011 19392 15020
rect 19340 14977 19349 15011
rect 19349 14977 19383 15011
rect 19383 14977 19392 15011
rect 19340 14968 19392 14977
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 22376 15104 22428 15156
rect 22836 15104 22888 15156
rect 23664 15104 23716 15156
rect 18880 14900 18932 14909
rect 20904 15036 20956 15088
rect 22284 15036 22336 15088
rect 22652 15036 22704 15088
rect 23848 15079 23900 15088
rect 23848 15045 23857 15079
rect 23857 15045 23891 15079
rect 23891 15045 23900 15079
rect 23848 15036 23900 15045
rect 24952 15104 25004 15156
rect 26056 15147 26108 15156
rect 26056 15113 26065 15147
rect 26065 15113 26099 15147
rect 26099 15113 26108 15147
rect 26056 15104 26108 15113
rect 24492 15036 24544 15088
rect 24860 15036 24912 15088
rect 9956 14764 10008 14816
rect 12348 14807 12400 14816
rect 12348 14773 12357 14807
rect 12357 14773 12391 14807
rect 12391 14773 12400 14807
rect 12348 14764 12400 14773
rect 15108 14807 15160 14816
rect 15108 14773 15117 14807
rect 15117 14773 15151 14807
rect 15151 14773 15160 14807
rect 15108 14764 15160 14773
rect 23020 14943 23072 14952
rect 23020 14909 23029 14943
rect 23029 14909 23063 14943
rect 23063 14909 23072 14943
rect 23020 14900 23072 14909
rect 23664 14832 23716 14884
rect 24124 14968 24176 15020
rect 25596 14968 25648 15020
rect 24308 14943 24360 14952
rect 24308 14909 24317 14943
rect 24317 14909 24351 14943
rect 24351 14909 24360 14943
rect 24308 14900 24360 14909
rect 25228 14900 25280 14952
rect 19892 14764 19944 14816
rect 21364 14807 21416 14816
rect 21364 14773 21373 14807
rect 21373 14773 21407 14807
rect 21407 14773 21416 14807
rect 21364 14764 21416 14773
rect 23112 14807 23164 14816
rect 23112 14773 23121 14807
rect 23121 14773 23155 14807
rect 23155 14773 23164 14807
rect 23112 14764 23164 14773
rect 23572 14807 23624 14816
rect 23572 14773 23581 14807
rect 23581 14773 23615 14807
rect 23615 14773 23624 14807
rect 23572 14764 23624 14773
rect 23848 14764 23900 14816
rect 24124 14764 24176 14816
rect 25136 14764 25188 14816
rect 25688 14764 25740 14816
rect 4124 14662 4176 14714
rect 4188 14662 4240 14714
rect 4252 14662 4304 14714
rect 4316 14662 4368 14714
rect 4380 14662 4432 14714
rect 10472 14662 10524 14714
rect 10536 14662 10588 14714
rect 10600 14662 10652 14714
rect 10664 14662 10716 14714
rect 10728 14662 10780 14714
rect 16820 14662 16872 14714
rect 16884 14662 16936 14714
rect 16948 14662 17000 14714
rect 17012 14662 17064 14714
rect 17076 14662 17128 14714
rect 23168 14662 23220 14714
rect 23232 14662 23284 14714
rect 23296 14662 23348 14714
rect 23360 14662 23412 14714
rect 23424 14662 23476 14714
rect 2320 14603 2372 14612
rect 2320 14569 2329 14603
rect 2329 14569 2363 14603
rect 2363 14569 2372 14603
rect 2320 14560 2372 14569
rect 6644 14560 6696 14612
rect 7656 14560 7708 14612
rect 1952 14331 2004 14340
rect 1952 14297 1961 14331
rect 1961 14297 1995 14331
rect 1995 14297 2004 14331
rect 1952 14288 2004 14297
rect 3240 14356 3292 14408
rect 3424 14356 3476 14408
rect 4712 14424 4764 14476
rect 5448 14424 5500 14476
rect 3056 14288 3108 14340
rect 2228 14263 2280 14272
rect 2228 14229 2237 14263
rect 2237 14229 2271 14263
rect 2271 14229 2280 14263
rect 2228 14220 2280 14229
rect 2688 14263 2740 14272
rect 2688 14229 2697 14263
rect 2697 14229 2731 14263
rect 2731 14229 2740 14263
rect 2688 14220 2740 14229
rect 2872 14220 2924 14272
rect 3148 14263 3200 14272
rect 3148 14229 3157 14263
rect 3157 14229 3191 14263
rect 3191 14229 3200 14263
rect 3148 14220 3200 14229
rect 4804 14288 4856 14340
rect 5724 14356 5776 14408
rect 6000 14356 6052 14408
rect 9588 14560 9640 14612
rect 12348 14603 12400 14612
rect 12348 14569 12378 14603
rect 12378 14569 12400 14603
rect 12348 14560 12400 14569
rect 15016 14560 15068 14612
rect 16396 14560 16448 14612
rect 17408 14560 17460 14612
rect 18880 14560 18932 14612
rect 19340 14560 19392 14612
rect 22836 14603 22888 14612
rect 22836 14569 22845 14603
rect 22845 14569 22879 14603
rect 22879 14569 22888 14603
rect 22836 14560 22888 14569
rect 9772 14492 9824 14544
rect 18420 14492 18472 14544
rect 8760 14424 8812 14476
rect 11244 14424 11296 14476
rect 8300 14356 8352 14408
rect 9680 14356 9732 14408
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 6828 14288 6880 14340
rect 9864 14288 9916 14340
rect 10140 14288 10192 14340
rect 12624 14288 12676 14340
rect 15292 14424 15344 14476
rect 22192 14492 22244 14544
rect 23756 14560 23808 14612
rect 23848 14603 23900 14612
rect 23848 14569 23857 14603
rect 23857 14569 23891 14603
rect 23891 14569 23900 14603
rect 23848 14560 23900 14569
rect 24032 14560 24084 14612
rect 15936 14356 15988 14408
rect 14648 14288 14700 14340
rect 17592 14356 17644 14408
rect 21364 14424 21416 14476
rect 23020 14467 23072 14476
rect 23020 14433 23029 14467
rect 23029 14433 23063 14467
rect 23063 14433 23072 14467
rect 23020 14424 23072 14433
rect 18788 14399 18840 14408
rect 18788 14365 18797 14399
rect 18797 14365 18831 14399
rect 18831 14365 18840 14399
rect 18788 14356 18840 14365
rect 19616 14356 19668 14408
rect 20628 14399 20680 14408
rect 20628 14365 20637 14399
rect 20637 14365 20671 14399
rect 20671 14365 20680 14399
rect 20628 14356 20680 14365
rect 21088 14356 21140 14408
rect 19524 14288 19576 14340
rect 23572 14356 23624 14408
rect 24216 14356 24268 14408
rect 25412 14399 25464 14408
rect 25412 14365 25421 14399
rect 25421 14365 25455 14399
rect 25455 14365 25464 14399
rect 25412 14356 25464 14365
rect 3608 14220 3660 14272
rect 5356 14263 5408 14272
rect 5356 14229 5365 14263
rect 5365 14229 5399 14263
rect 5399 14229 5408 14263
rect 5356 14220 5408 14229
rect 5540 14220 5592 14272
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 8392 14263 8444 14272
rect 8392 14229 8401 14263
rect 8401 14229 8435 14263
rect 8435 14229 8444 14263
rect 8392 14220 8444 14229
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 8760 14220 8812 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 12440 14220 12492 14272
rect 14096 14220 14148 14272
rect 14188 14220 14240 14272
rect 15476 14220 15528 14272
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 16856 14263 16908 14272
rect 16856 14229 16865 14263
rect 16865 14229 16899 14263
rect 16899 14229 16908 14263
rect 16856 14220 16908 14229
rect 19340 14263 19392 14272
rect 19340 14229 19349 14263
rect 19349 14229 19383 14263
rect 19383 14229 19392 14263
rect 19340 14220 19392 14229
rect 20904 14220 20956 14272
rect 22652 14220 22704 14272
rect 24032 14288 24084 14340
rect 24952 14288 25004 14340
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 24768 14263 24820 14272
rect 24768 14229 24777 14263
rect 24777 14229 24811 14263
rect 24811 14229 24820 14263
rect 24768 14220 24820 14229
rect 25504 14220 25556 14272
rect 7298 14118 7350 14170
rect 7362 14118 7414 14170
rect 7426 14118 7478 14170
rect 7490 14118 7542 14170
rect 7554 14118 7606 14170
rect 13646 14118 13698 14170
rect 13710 14118 13762 14170
rect 13774 14118 13826 14170
rect 13838 14118 13890 14170
rect 13902 14118 13954 14170
rect 19994 14118 20046 14170
rect 20058 14118 20110 14170
rect 20122 14118 20174 14170
rect 20186 14118 20238 14170
rect 20250 14118 20302 14170
rect 26342 14118 26394 14170
rect 26406 14118 26458 14170
rect 26470 14118 26522 14170
rect 26534 14118 26586 14170
rect 26598 14118 26650 14170
rect 1952 14016 2004 14068
rect 2228 14016 2280 14068
rect 2412 14016 2464 14068
rect 3148 14016 3200 14068
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 3608 13991 3660 14000
rect 3608 13957 3617 13991
rect 3617 13957 3651 13991
rect 3651 13957 3660 13991
rect 3608 13948 3660 13957
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 2872 13880 2924 13932
rect 3240 13923 3292 13932
rect 3240 13889 3249 13923
rect 3249 13889 3283 13923
rect 3283 13889 3292 13923
rect 3240 13880 3292 13889
rect 3608 13812 3660 13864
rect 4712 13812 4764 13864
rect 5356 14016 5408 14068
rect 5540 14016 5592 14068
rect 6736 14016 6788 14068
rect 7104 13948 7156 14000
rect 8760 13948 8812 14000
rect 5172 13923 5224 13932
rect 5172 13889 5181 13923
rect 5181 13889 5215 13923
rect 5215 13889 5224 13923
rect 5172 13880 5224 13889
rect 5356 13923 5408 13932
rect 5356 13889 5391 13923
rect 5391 13889 5408 13923
rect 5356 13880 5408 13889
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 11980 13948 12032 14000
rect 5908 13812 5960 13864
rect 10048 13812 10100 13864
rect 11520 13923 11572 13932
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 15384 14016 15436 14068
rect 15936 14059 15988 14068
rect 15936 14025 15945 14059
rect 15945 14025 15979 14059
rect 15979 14025 15988 14059
rect 15936 14016 15988 14025
rect 16672 14016 16724 14068
rect 16856 14016 16908 14068
rect 19248 14016 19300 14068
rect 12624 13812 12676 13864
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 15568 13880 15620 13932
rect 10876 13787 10928 13796
rect 10876 13753 10885 13787
rect 10885 13753 10919 13787
rect 10919 13753 10928 13787
rect 10876 13744 10928 13753
rect 13912 13744 13964 13796
rect 2780 13676 2832 13728
rect 3240 13676 3292 13728
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 4988 13676 5040 13728
rect 5356 13676 5408 13728
rect 5632 13719 5684 13728
rect 5632 13685 5641 13719
rect 5641 13685 5675 13719
rect 5675 13685 5684 13719
rect 5632 13676 5684 13685
rect 7012 13676 7064 13728
rect 9128 13676 9180 13728
rect 11612 13719 11664 13728
rect 11612 13685 11621 13719
rect 11621 13685 11655 13719
rect 11655 13685 11664 13719
rect 11612 13676 11664 13685
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 17960 13880 18012 13932
rect 20812 13948 20864 14000
rect 22192 13923 22244 13932
rect 18052 13812 18104 13864
rect 19892 13812 19944 13864
rect 20444 13812 20496 13864
rect 20628 13812 20680 13864
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 23020 13948 23072 14000
rect 23940 14016 23992 14068
rect 24768 14016 24820 14068
rect 23664 13948 23716 14000
rect 23940 13880 23992 13932
rect 25504 13948 25556 14000
rect 19340 13744 19392 13796
rect 21732 13744 21784 13796
rect 22652 13812 22704 13864
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 24952 13880 25004 13932
rect 25228 13812 25280 13864
rect 24860 13744 24912 13796
rect 14556 13676 14608 13728
rect 17316 13719 17368 13728
rect 17316 13685 17325 13719
rect 17325 13685 17359 13719
rect 17359 13685 17368 13719
rect 17316 13676 17368 13685
rect 17592 13719 17644 13728
rect 17592 13685 17601 13719
rect 17601 13685 17635 13719
rect 17635 13685 17644 13719
rect 17592 13676 17644 13685
rect 19248 13676 19300 13728
rect 21364 13676 21416 13728
rect 22652 13676 22704 13728
rect 23848 13676 23900 13728
rect 24032 13676 24084 13728
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 4124 13574 4176 13626
rect 4188 13574 4240 13626
rect 4252 13574 4304 13626
rect 4316 13574 4368 13626
rect 4380 13574 4432 13626
rect 10472 13574 10524 13626
rect 10536 13574 10588 13626
rect 10600 13574 10652 13626
rect 10664 13574 10716 13626
rect 10728 13574 10780 13626
rect 16820 13574 16872 13626
rect 16884 13574 16936 13626
rect 16948 13574 17000 13626
rect 17012 13574 17064 13626
rect 17076 13574 17128 13626
rect 23168 13574 23220 13626
rect 23232 13574 23284 13626
rect 23296 13574 23348 13626
rect 23360 13574 23412 13626
rect 23424 13574 23476 13626
rect 2688 13472 2740 13524
rect 3516 13472 3568 13524
rect 5080 13472 5132 13524
rect 5172 13472 5224 13524
rect 6368 13472 6420 13524
rect 8208 13472 8260 13524
rect 8392 13472 8444 13524
rect 14464 13472 14516 13524
rect 15384 13515 15436 13524
rect 15384 13481 15393 13515
rect 15393 13481 15427 13515
rect 15427 13481 15436 13515
rect 15384 13472 15436 13481
rect 3608 13404 3660 13456
rect 4436 13404 4488 13456
rect 9864 13404 9916 13456
rect 1676 13336 1728 13388
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 5540 13336 5592 13388
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 2964 13200 3016 13252
rect 3516 13200 3568 13252
rect 4436 13311 4488 13320
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 7012 13336 7064 13388
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 9772 13336 9824 13388
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 11244 13336 11296 13388
rect 11612 13336 11664 13388
rect 12900 13336 12952 13388
rect 13912 13336 13964 13388
rect 14648 13336 14700 13388
rect 4712 13200 4764 13252
rect 5080 13200 5132 13252
rect 6828 13243 6880 13252
rect 6828 13209 6837 13243
rect 6837 13209 6871 13243
rect 6871 13209 6880 13243
rect 6828 13200 6880 13209
rect 8944 13268 8996 13320
rect 9956 13268 10008 13320
rect 10876 13268 10928 13320
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 15292 13268 15344 13320
rect 18052 13472 18104 13524
rect 17592 13404 17644 13456
rect 17316 13336 17368 13388
rect 17500 13379 17552 13388
rect 17500 13345 17509 13379
rect 17509 13345 17543 13379
rect 17543 13345 17552 13379
rect 17500 13336 17552 13345
rect 18420 13472 18472 13524
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 20628 13472 20680 13524
rect 23664 13472 23716 13524
rect 24216 13472 24268 13524
rect 24492 13472 24544 13524
rect 19524 13336 19576 13388
rect 12624 13200 12676 13252
rect 3148 13132 3200 13184
rect 4620 13132 4672 13184
rect 4988 13132 5040 13184
rect 5908 13132 5960 13184
rect 11152 13132 11204 13184
rect 13176 13132 13228 13184
rect 14096 13132 14148 13184
rect 15568 13200 15620 13252
rect 20904 13268 20956 13320
rect 21364 13336 21416 13388
rect 23848 13336 23900 13388
rect 24400 13268 24452 13320
rect 20444 13200 20496 13252
rect 24032 13243 24084 13252
rect 24032 13209 24041 13243
rect 24041 13209 24075 13243
rect 24075 13209 24084 13243
rect 24032 13200 24084 13209
rect 24216 13243 24268 13252
rect 24216 13209 24225 13243
rect 24225 13209 24259 13243
rect 24259 13209 24268 13243
rect 24216 13200 24268 13209
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 19800 13132 19852 13184
rect 23020 13132 23072 13184
rect 24124 13132 24176 13184
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 25044 13311 25096 13320
rect 25044 13277 25053 13311
rect 25053 13277 25087 13311
rect 25087 13277 25096 13311
rect 25044 13268 25096 13277
rect 24676 13243 24728 13252
rect 24676 13209 24685 13243
rect 24685 13209 24719 13243
rect 24719 13209 24728 13243
rect 24676 13200 24728 13209
rect 24768 13243 24820 13252
rect 24768 13209 24777 13243
rect 24777 13209 24811 13243
rect 24811 13209 24820 13243
rect 24768 13200 24820 13209
rect 26148 13311 26200 13320
rect 26148 13277 26157 13311
rect 26157 13277 26191 13311
rect 26191 13277 26200 13311
rect 26148 13268 26200 13277
rect 25228 13243 25280 13252
rect 25228 13209 25237 13243
rect 25237 13209 25271 13243
rect 25271 13209 25280 13243
rect 25228 13200 25280 13209
rect 25504 13200 25556 13252
rect 25964 13175 26016 13184
rect 25964 13141 25973 13175
rect 25973 13141 26007 13175
rect 26007 13141 26016 13175
rect 25964 13132 26016 13141
rect 7298 13030 7350 13082
rect 7362 13030 7414 13082
rect 7426 13030 7478 13082
rect 7490 13030 7542 13082
rect 7554 13030 7606 13082
rect 13646 13030 13698 13082
rect 13710 13030 13762 13082
rect 13774 13030 13826 13082
rect 13838 13030 13890 13082
rect 13902 13030 13954 13082
rect 19994 13030 20046 13082
rect 20058 13030 20110 13082
rect 20122 13030 20174 13082
rect 20186 13030 20238 13082
rect 20250 13030 20302 13082
rect 26342 13030 26394 13082
rect 26406 13030 26458 13082
rect 26470 13030 26522 13082
rect 26534 13030 26586 13082
rect 26598 13030 26650 13082
rect 1676 12928 1728 12980
rect 4896 12928 4948 12980
rect 2872 12860 2924 12912
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 2780 12724 2832 12776
rect 3148 12724 3200 12776
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 3332 12767 3384 12776
rect 3332 12733 3341 12767
rect 3341 12733 3375 12767
rect 3375 12733 3384 12767
rect 3332 12724 3384 12733
rect 3056 12656 3108 12708
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5632 12860 5684 12912
rect 7012 12928 7064 12980
rect 7104 12928 7156 12980
rect 9128 12928 9180 12980
rect 9772 12928 9824 12980
rect 14556 12928 14608 12980
rect 6276 12860 6328 12912
rect 9220 12860 9272 12912
rect 12440 12860 12492 12912
rect 15568 12860 15620 12912
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 8852 12792 8904 12844
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 4436 12656 4488 12708
rect 5540 12656 5592 12708
rect 6000 12656 6052 12708
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 9680 12792 9732 12844
rect 14096 12792 14148 12844
rect 17408 12860 17460 12912
rect 17960 12928 18012 12980
rect 19248 12928 19300 12980
rect 23848 12928 23900 12980
rect 10048 12724 10100 12776
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 5632 12588 5684 12640
rect 6368 12631 6420 12640
rect 6368 12597 6377 12631
rect 6377 12597 6411 12631
rect 6411 12597 6420 12631
rect 6368 12588 6420 12597
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 8944 12588 8996 12640
rect 10140 12588 10192 12640
rect 11888 12767 11940 12776
rect 11888 12733 11897 12767
rect 11897 12733 11931 12767
rect 11931 12733 11940 12767
rect 11888 12724 11940 12733
rect 23940 12903 23992 12912
rect 23940 12869 23949 12903
rect 23949 12869 23983 12903
rect 23983 12869 23992 12903
rect 23940 12860 23992 12869
rect 24676 12928 24728 12980
rect 24768 12928 24820 12980
rect 24584 12860 24636 12912
rect 20444 12835 20496 12844
rect 20444 12801 20453 12835
rect 20453 12801 20487 12835
rect 20487 12801 20496 12835
rect 20444 12792 20496 12801
rect 20904 12835 20956 12844
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 19432 12724 19484 12776
rect 20812 12724 20864 12776
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 21732 12792 21784 12844
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 23572 12835 23624 12844
rect 23572 12801 23581 12835
rect 23581 12801 23615 12835
rect 23615 12801 23624 12835
rect 23572 12792 23624 12801
rect 25044 12792 25096 12844
rect 25136 12792 25188 12844
rect 21548 12724 21600 12776
rect 24032 12724 24084 12776
rect 24492 12724 24544 12776
rect 26056 12792 26108 12844
rect 22652 12656 22704 12708
rect 12992 12588 13044 12640
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 21916 12631 21968 12640
rect 21916 12597 21925 12631
rect 21925 12597 21959 12631
rect 21959 12597 21968 12631
rect 21916 12588 21968 12597
rect 23664 12631 23716 12640
rect 23664 12597 23673 12631
rect 23673 12597 23707 12631
rect 23707 12597 23716 12631
rect 23664 12588 23716 12597
rect 4124 12486 4176 12538
rect 4188 12486 4240 12538
rect 4252 12486 4304 12538
rect 4316 12486 4368 12538
rect 4380 12486 4432 12538
rect 10472 12486 10524 12538
rect 10536 12486 10588 12538
rect 10600 12486 10652 12538
rect 10664 12486 10716 12538
rect 10728 12486 10780 12538
rect 16820 12486 16872 12538
rect 16884 12486 16936 12538
rect 16948 12486 17000 12538
rect 17012 12486 17064 12538
rect 17076 12486 17128 12538
rect 23168 12486 23220 12538
rect 23232 12486 23284 12538
rect 23296 12486 23348 12538
rect 23360 12486 23412 12538
rect 23424 12486 23476 12538
rect 4988 12427 5040 12436
rect 4988 12393 4997 12427
rect 4997 12393 5031 12427
rect 5031 12393 5040 12427
rect 4988 12384 5040 12393
rect 6276 12427 6328 12436
rect 6276 12393 6285 12427
rect 6285 12393 6319 12427
rect 6319 12393 6328 12427
rect 6276 12384 6328 12393
rect 6644 12384 6696 12436
rect 11888 12384 11940 12436
rect 14280 12384 14332 12436
rect 15200 12384 15252 12436
rect 19248 12384 19300 12436
rect 20904 12384 20956 12436
rect 23848 12384 23900 12436
rect 26056 12384 26108 12436
rect 7748 12316 7800 12368
rect 11520 12316 11572 12368
rect 4620 12248 4672 12300
rect 3884 12223 3936 12232
rect 3884 12189 3893 12223
rect 3893 12189 3927 12223
rect 3927 12189 3936 12223
rect 3884 12180 3936 12189
rect 4528 12180 4580 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 5632 12112 5684 12164
rect 6000 12112 6052 12164
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 6828 12180 6880 12232
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 8116 12180 8168 12232
rect 9496 12248 9548 12300
rect 11060 12248 11112 12300
rect 9588 12223 9640 12232
rect 9588 12189 9597 12223
rect 9597 12189 9631 12223
rect 9631 12189 9640 12223
rect 9588 12180 9640 12189
rect 14556 12248 14608 12300
rect 9312 12112 9364 12164
rect 3424 12044 3476 12096
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 8760 12044 8812 12096
rect 11244 12112 11296 12164
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 15660 12316 15712 12368
rect 20444 12316 20496 12368
rect 19340 12248 19392 12300
rect 19892 12248 19944 12300
rect 20904 12248 20956 12300
rect 22744 12248 22796 12300
rect 24308 12248 24360 12300
rect 14188 12112 14240 12164
rect 15476 12180 15528 12232
rect 16396 12180 16448 12232
rect 19248 12223 19300 12232
rect 19248 12189 19257 12223
rect 19257 12189 19291 12223
rect 19291 12189 19300 12223
rect 19248 12180 19300 12189
rect 19524 12223 19576 12232
rect 19524 12189 19533 12223
rect 19533 12189 19567 12223
rect 19567 12189 19576 12223
rect 19524 12180 19576 12189
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 19616 12180 19668 12189
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 19800 12180 19852 12232
rect 15200 12112 15252 12164
rect 21824 12180 21876 12232
rect 20812 12155 20864 12164
rect 20812 12121 20821 12155
rect 20821 12121 20855 12155
rect 20855 12121 20864 12155
rect 20812 12112 20864 12121
rect 21548 12112 21600 12164
rect 10508 12044 10560 12096
rect 14464 12044 14516 12096
rect 15568 12044 15620 12096
rect 16304 12044 16356 12096
rect 19340 12044 19392 12096
rect 19708 12044 19760 12096
rect 19892 12087 19944 12096
rect 19892 12053 19901 12087
rect 19901 12053 19935 12087
rect 19935 12053 19944 12087
rect 19892 12044 19944 12053
rect 20260 12044 20312 12096
rect 20444 12044 20496 12096
rect 21180 12044 21232 12096
rect 21732 12044 21784 12096
rect 23020 12112 23072 12164
rect 23756 12112 23808 12164
rect 24124 12112 24176 12164
rect 23480 12044 23532 12096
rect 7298 11942 7350 11994
rect 7362 11942 7414 11994
rect 7426 11942 7478 11994
rect 7490 11942 7542 11994
rect 7554 11942 7606 11994
rect 13646 11942 13698 11994
rect 13710 11942 13762 11994
rect 13774 11942 13826 11994
rect 13838 11942 13890 11994
rect 13902 11942 13954 11994
rect 19994 11942 20046 11994
rect 20058 11942 20110 11994
rect 20122 11942 20174 11994
rect 20186 11942 20238 11994
rect 20250 11942 20302 11994
rect 26342 11942 26394 11994
rect 26406 11942 26458 11994
rect 26470 11942 26522 11994
rect 26534 11942 26586 11994
rect 26598 11942 26650 11994
rect 3516 11840 3568 11892
rect 2872 11815 2924 11824
rect 2872 11781 2881 11815
rect 2881 11781 2915 11815
rect 2915 11781 2924 11815
rect 2872 11772 2924 11781
rect 4804 11840 4856 11892
rect 7104 11840 7156 11892
rect 9312 11840 9364 11892
rect 9588 11840 9640 11892
rect 10508 11840 10560 11892
rect 11244 11840 11296 11892
rect 12716 11840 12768 11892
rect 12992 11840 13044 11892
rect 15476 11840 15528 11892
rect 15660 11840 15712 11892
rect 18144 11840 18196 11892
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 4436 11747 4488 11756
rect 4436 11713 4445 11747
rect 4445 11713 4479 11747
rect 4479 11713 4488 11747
rect 4436 11704 4488 11713
rect 4712 11704 4764 11756
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 5264 11704 5316 11756
rect 5724 11747 5776 11756
rect 5724 11713 5733 11747
rect 5733 11713 5767 11747
rect 5767 11713 5776 11747
rect 5724 11704 5776 11713
rect 6552 11704 6604 11756
rect 8852 11772 8904 11824
rect 6368 11636 6420 11688
rect 6828 11636 6880 11688
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 8484 11704 8536 11756
rect 8944 11747 8996 11756
rect 8944 11713 8953 11747
rect 8953 11713 8987 11747
rect 8987 11713 8996 11747
rect 8944 11704 8996 11713
rect 9680 11815 9732 11824
rect 9680 11781 9689 11815
rect 9689 11781 9723 11815
rect 9723 11781 9732 11815
rect 9680 11772 9732 11781
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 11152 11704 11204 11756
rect 8116 11636 8168 11688
rect 3056 11568 3108 11620
rect 4436 11568 4488 11620
rect 2136 11500 2188 11552
rect 3148 11500 3200 11552
rect 5080 11500 5132 11552
rect 5264 11500 5316 11552
rect 9220 11568 9272 11620
rect 10048 11636 10100 11688
rect 13176 11704 13228 11756
rect 13544 11704 13596 11756
rect 14188 11772 14240 11824
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 8852 11500 8904 11552
rect 14096 11568 14148 11620
rect 14464 11772 14516 11824
rect 14648 11704 14700 11756
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 16396 11772 16448 11824
rect 17408 11772 17460 11824
rect 18696 11815 18748 11824
rect 18696 11781 18705 11815
rect 18705 11781 18739 11815
rect 18739 11781 18748 11815
rect 18696 11772 18748 11781
rect 19524 11840 19576 11892
rect 20352 11840 20404 11892
rect 22744 11840 22796 11892
rect 24492 11840 24544 11892
rect 15936 11747 15988 11756
rect 15936 11713 15969 11747
rect 15969 11713 15988 11747
rect 15936 11704 15988 11713
rect 17224 11704 17276 11756
rect 16488 11636 16540 11688
rect 17960 11747 18012 11756
rect 17960 11713 17969 11747
rect 17969 11713 18003 11747
rect 18003 11713 18012 11747
rect 17960 11704 18012 11713
rect 19616 11747 19668 11756
rect 19616 11713 19625 11747
rect 19625 11713 19659 11747
rect 19659 11713 19668 11747
rect 19616 11704 19668 11713
rect 19708 11747 19760 11756
rect 19708 11713 19717 11747
rect 19717 11713 19751 11747
rect 19751 11713 19760 11747
rect 19708 11704 19760 11713
rect 21180 11747 21232 11756
rect 21180 11713 21189 11747
rect 21189 11713 21223 11747
rect 21223 11713 21232 11747
rect 21180 11704 21232 11713
rect 18052 11636 18104 11688
rect 18512 11636 18564 11688
rect 20444 11568 20496 11620
rect 14188 11500 14240 11552
rect 14556 11543 14608 11552
rect 14556 11509 14565 11543
rect 14565 11509 14599 11543
rect 14599 11509 14608 11543
rect 14556 11500 14608 11509
rect 14648 11543 14700 11552
rect 14648 11509 14657 11543
rect 14657 11509 14691 11543
rect 14691 11509 14700 11543
rect 14648 11500 14700 11509
rect 15292 11500 15344 11552
rect 15568 11500 15620 11552
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 16028 11543 16080 11552
rect 16028 11509 16037 11543
rect 16037 11509 16071 11543
rect 16071 11509 16080 11543
rect 16028 11500 16080 11509
rect 18236 11500 18288 11552
rect 19616 11500 19668 11552
rect 21272 11500 21324 11552
rect 23480 11772 23532 11824
rect 23664 11636 23716 11688
rect 25964 11568 26016 11620
rect 4124 11398 4176 11450
rect 4188 11398 4240 11450
rect 4252 11398 4304 11450
rect 4316 11398 4368 11450
rect 4380 11398 4432 11450
rect 10472 11398 10524 11450
rect 10536 11398 10588 11450
rect 10600 11398 10652 11450
rect 10664 11398 10716 11450
rect 10728 11398 10780 11450
rect 16820 11398 16872 11450
rect 16884 11398 16936 11450
rect 16948 11398 17000 11450
rect 17012 11398 17064 11450
rect 17076 11398 17128 11450
rect 23168 11398 23220 11450
rect 23232 11398 23284 11450
rect 23296 11398 23348 11450
rect 23360 11398 23412 11450
rect 23424 11398 23476 11450
rect 2136 11296 2188 11348
rect 2872 11296 2924 11348
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 3884 11296 3936 11348
rect 3424 11228 3476 11280
rect 4620 11339 4672 11348
rect 4620 11305 4629 11339
rect 4629 11305 4663 11339
rect 4663 11305 4672 11339
rect 4620 11296 4672 11305
rect 4988 11296 5040 11348
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 3884 11160 3936 11212
rect 4712 11228 4764 11280
rect 3148 11024 3200 11076
rect 3700 11024 3752 11076
rect 4804 11160 4856 11212
rect 5540 11271 5592 11280
rect 5540 11237 5549 11271
rect 5549 11237 5583 11271
rect 5583 11237 5592 11271
rect 5540 11228 5592 11237
rect 5448 11092 5500 11144
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 4528 11024 4580 11076
rect 5724 11092 5776 11144
rect 4344 10956 4396 11008
rect 5172 10956 5224 11008
rect 6184 11024 6236 11076
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 8116 11296 8168 11348
rect 9680 11296 9732 11348
rect 9772 11296 9824 11348
rect 15200 11296 15252 11348
rect 15844 11296 15896 11348
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 17960 11296 18012 11348
rect 8576 11160 8628 11212
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 8852 11092 8904 11144
rect 9220 11024 9272 11076
rect 14464 11092 14516 11144
rect 14740 11092 14792 11144
rect 15568 11160 15620 11212
rect 13544 11024 13596 11076
rect 16028 11228 16080 11280
rect 18236 11228 18288 11280
rect 18696 11228 18748 11280
rect 17868 11203 17920 11212
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 18144 11160 18196 11212
rect 19616 11160 19668 11212
rect 21272 11203 21324 11212
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 22744 11296 22796 11348
rect 8300 10999 8352 11008
rect 8300 10965 8309 10999
rect 8309 10965 8343 10999
rect 8343 10965 8352 10999
rect 8300 10956 8352 10965
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 15476 11024 15528 11076
rect 15200 10956 15252 11008
rect 15292 10956 15344 11008
rect 16304 11024 16356 11076
rect 16488 11067 16540 11076
rect 16488 11033 16497 11067
rect 16497 11033 16531 11067
rect 16531 11033 16540 11067
rect 16488 11024 16540 11033
rect 16672 11067 16724 11076
rect 16672 11033 16681 11067
rect 16681 11033 16715 11067
rect 16715 11033 16724 11067
rect 16672 11024 16724 11033
rect 17224 11024 17276 11076
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 19156 11092 19208 11144
rect 21640 11135 21692 11144
rect 21640 11101 21649 11135
rect 21649 11101 21683 11135
rect 21683 11101 21692 11135
rect 21640 11092 21692 11101
rect 19800 11024 19852 11076
rect 18696 10956 18748 11008
rect 19524 10956 19576 11008
rect 19616 10956 19668 11008
rect 22100 11024 22152 11076
rect 7298 10854 7350 10906
rect 7362 10854 7414 10906
rect 7426 10854 7478 10906
rect 7490 10854 7542 10906
rect 7554 10854 7606 10906
rect 13646 10854 13698 10906
rect 13710 10854 13762 10906
rect 13774 10854 13826 10906
rect 13838 10854 13890 10906
rect 13902 10854 13954 10906
rect 19994 10854 20046 10906
rect 20058 10854 20110 10906
rect 20122 10854 20174 10906
rect 20186 10854 20238 10906
rect 20250 10854 20302 10906
rect 26342 10854 26394 10906
rect 26406 10854 26458 10906
rect 26470 10854 26522 10906
rect 26534 10854 26586 10906
rect 26598 10854 26650 10906
rect 3792 10752 3844 10804
rect 4712 10752 4764 10804
rect 5264 10752 5316 10804
rect 3056 10727 3108 10736
rect 3056 10693 3065 10727
rect 3065 10693 3099 10727
rect 3099 10693 3108 10727
rect 3056 10684 3108 10693
rect 3516 10684 3568 10736
rect 3700 10659 3752 10668
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 4344 10727 4396 10736
rect 4344 10693 4353 10727
rect 4353 10693 4387 10727
rect 4387 10693 4396 10727
rect 4344 10684 4396 10693
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 4436 10659 4488 10692
rect 4436 10640 4445 10659
rect 4445 10640 4479 10659
rect 4479 10640 4488 10659
rect 4620 10684 4672 10736
rect 5172 10684 5224 10736
rect 5724 10752 5776 10804
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 8944 10752 8996 10804
rect 9680 10752 9732 10804
rect 15660 10752 15712 10804
rect 16488 10752 16540 10804
rect 6828 10684 6880 10736
rect 5080 10548 5132 10600
rect 7196 10616 7248 10668
rect 8300 10727 8352 10736
rect 8300 10693 8309 10727
rect 8309 10693 8343 10727
rect 8343 10693 8352 10727
rect 8300 10684 8352 10693
rect 12808 10684 12860 10736
rect 15384 10727 15436 10736
rect 15384 10693 15393 10727
rect 15393 10693 15427 10727
rect 15427 10693 15436 10727
rect 15384 10684 15436 10693
rect 9312 10616 9364 10668
rect 10876 10616 10928 10668
rect 6184 10591 6236 10600
rect 6184 10557 6193 10591
rect 6193 10557 6227 10591
rect 6227 10557 6236 10591
rect 6184 10548 6236 10557
rect 6644 10548 6696 10600
rect 12532 10616 12584 10668
rect 13176 10616 13228 10668
rect 14740 10616 14792 10668
rect 3608 10480 3660 10532
rect 4436 10480 4488 10532
rect 4620 10480 4672 10532
rect 5448 10480 5500 10532
rect 12716 10548 12768 10600
rect 14188 10548 14240 10600
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 15568 10659 15620 10668
rect 15568 10625 15613 10659
rect 15613 10625 15620 10659
rect 15568 10616 15620 10625
rect 16396 10659 16448 10668
rect 16396 10625 16405 10659
rect 16405 10625 16439 10659
rect 16439 10625 16448 10659
rect 16396 10616 16448 10625
rect 16672 10659 16724 10668
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 18512 10752 18564 10804
rect 17868 10727 17920 10736
rect 17868 10693 17877 10727
rect 17877 10693 17911 10727
rect 17911 10693 17920 10727
rect 17868 10684 17920 10693
rect 18328 10684 18380 10736
rect 19524 10684 19576 10736
rect 19800 10684 19852 10736
rect 21640 10684 21692 10736
rect 16304 10548 16356 10600
rect 9404 10480 9456 10532
rect 14648 10480 14700 10532
rect 15384 10480 15436 10532
rect 15568 10480 15620 10532
rect 17408 10616 17460 10668
rect 19340 10616 19392 10668
rect 19892 10659 19944 10668
rect 19892 10625 19901 10659
rect 19901 10625 19935 10659
rect 19935 10625 19944 10659
rect 19892 10616 19944 10625
rect 20352 10616 20404 10668
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2136 10412 2188 10421
rect 4528 10412 4580 10464
rect 8116 10412 8168 10464
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 12072 10412 12124 10464
rect 14280 10455 14332 10464
rect 14280 10421 14289 10455
rect 14289 10421 14323 10455
rect 14323 10421 14332 10455
rect 14280 10412 14332 10421
rect 15844 10455 15896 10464
rect 15844 10421 15853 10455
rect 15853 10421 15887 10455
rect 15887 10421 15896 10455
rect 15844 10412 15896 10421
rect 16488 10412 16540 10464
rect 18328 10548 18380 10600
rect 19616 10548 19668 10600
rect 22560 10591 22612 10600
rect 22560 10557 22569 10591
rect 22569 10557 22603 10591
rect 22603 10557 22612 10591
rect 22560 10548 22612 10557
rect 17224 10412 17276 10464
rect 18052 10412 18104 10464
rect 19248 10412 19300 10464
rect 4124 10310 4176 10362
rect 4188 10310 4240 10362
rect 4252 10310 4304 10362
rect 4316 10310 4368 10362
rect 4380 10310 4432 10362
rect 10472 10310 10524 10362
rect 10536 10310 10588 10362
rect 10600 10310 10652 10362
rect 10664 10310 10716 10362
rect 10728 10310 10780 10362
rect 16820 10310 16872 10362
rect 16884 10310 16936 10362
rect 16948 10310 17000 10362
rect 17012 10310 17064 10362
rect 17076 10310 17128 10362
rect 23168 10310 23220 10362
rect 23232 10310 23284 10362
rect 23296 10310 23348 10362
rect 23360 10310 23412 10362
rect 23424 10310 23476 10362
rect 2136 10208 2188 10260
rect 3608 10208 3660 10260
rect 4528 10208 4580 10260
rect 5540 10208 5592 10260
rect 6644 10251 6696 10260
rect 6644 10217 6653 10251
rect 6653 10217 6687 10251
rect 6687 10217 6696 10251
rect 6644 10208 6696 10217
rect 9404 10208 9456 10260
rect 9496 10208 9548 10260
rect 10968 10208 11020 10260
rect 15568 10251 15620 10260
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 15844 10208 15896 10260
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 16396 10208 16448 10260
rect 1400 10072 1452 10124
rect 1860 10072 1912 10124
rect 5540 10072 5592 10124
rect 6828 10072 6880 10124
rect 7196 10004 7248 10056
rect 7656 10004 7708 10056
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 8116 10004 8168 10056
rect 3148 9936 3200 9988
rect 3792 9936 3844 9988
rect 7012 9936 7064 9988
rect 11060 10072 11112 10124
rect 12808 10072 12860 10124
rect 13176 10072 13228 10124
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 19708 10208 19760 10260
rect 22744 10208 22796 10260
rect 16488 10072 16540 10124
rect 3884 9868 3936 9920
rect 6920 9868 6972 9920
rect 10140 9936 10192 9988
rect 11520 9979 11572 9988
rect 11520 9945 11529 9979
rect 11529 9945 11563 9979
rect 11563 9945 11572 9979
rect 11520 9936 11572 9945
rect 12900 9936 12952 9988
rect 14464 9936 14516 9988
rect 16120 10004 16172 10056
rect 17224 10072 17276 10124
rect 18880 10183 18932 10192
rect 18880 10149 18889 10183
rect 18889 10149 18923 10183
rect 18923 10149 18932 10183
rect 18880 10140 18932 10149
rect 19248 10140 19300 10192
rect 19800 10140 19852 10192
rect 18052 10004 18104 10056
rect 16304 9936 16356 9988
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 19616 10004 19668 10056
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 23756 10072 23808 10124
rect 23112 10004 23164 10056
rect 24584 10047 24636 10056
rect 24584 10013 24593 10047
rect 24593 10013 24627 10047
rect 24627 10013 24636 10047
rect 24584 10004 24636 10013
rect 25504 10047 25556 10056
rect 25504 10013 25513 10047
rect 25513 10013 25547 10047
rect 25547 10013 25556 10047
rect 25504 10004 25556 10013
rect 21180 9979 21232 9988
rect 21180 9945 21189 9979
rect 21189 9945 21223 9979
rect 21223 9945 21232 9979
rect 21180 9936 21232 9945
rect 22192 9936 22244 9988
rect 22836 9936 22888 9988
rect 24860 9936 24912 9988
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 11704 9868 11756 9920
rect 12348 9868 12400 9920
rect 12808 9868 12860 9920
rect 13360 9868 13412 9920
rect 15292 9868 15344 9920
rect 18144 9868 18196 9920
rect 20444 9868 20496 9920
rect 23020 9911 23072 9920
rect 23020 9877 23029 9911
rect 23029 9877 23063 9911
rect 23063 9877 23072 9911
rect 23020 9868 23072 9877
rect 23480 9911 23532 9920
rect 23480 9877 23505 9911
rect 23505 9877 23532 9911
rect 23480 9868 23532 9877
rect 23664 9911 23716 9920
rect 23664 9877 23673 9911
rect 23673 9877 23707 9911
rect 23707 9877 23716 9911
rect 23664 9868 23716 9877
rect 24400 9911 24452 9920
rect 24400 9877 24409 9911
rect 24409 9877 24443 9911
rect 24443 9877 24452 9911
rect 24400 9868 24452 9877
rect 25044 9868 25096 9920
rect 25320 9911 25372 9920
rect 25320 9877 25329 9911
rect 25329 9877 25363 9911
rect 25363 9877 25372 9911
rect 25320 9868 25372 9877
rect 7298 9766 7350 9818
rect 7362 9766 7414 9818
rect 7426 9766 7478 9818
rect 7490 9766 7542 9818
rect 7554 9766 7606 9818
rect 13646 9766 13698 9818
rect 13710 9766 13762 9818
rect 13774 9766 13826 9818
rect 13838 9766 13890 9818
rect 13902 9766 13954 9818
rect 19994 9766 20046 9818
rect 20058 9766 20110 9818
rect 20122 9766 20174 9818
rect 20186 9766 20238 9818
rect 20250 9766 20302 9818
rect 26342 9766 26394 9818
rect 26406 9766 26458 9818
rect 26470 9766 26522 9818
rect 26534 9766 26586 9818
rect 26598 9766 26650 9818
rect 5540 9664 5592 9716
rect 7012 9664 7064 9716
rect 7564 9664 7616 9716
rect 7656 9664 7708 9716
rect 7840 9664 7892 9716
rect 8116 9664 8168 9716
rect 9404 9664 9456 9716
rect 13268 9664 13320 9716
rect 1860 9528 1912 9580
rect 3884 9460 3936 9512
rect 3884 9324 3936 9376
rect 5172 9528 5224 9580
rect 7012 9528 7064 9580
rect 11060 9596 11112 9648
rect 18328 9596 18380 9648
rect 21180 9664 21232 9716
rect 7196 9460 7248 9512
rect 8208 9460 8260 9512
rect 8760 9460 8812 9512
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 7748 9367 7800 9376
rect 7748 9333 7757 9367
rect 7757 9333 7791 9367
rect 7791 9333 7800 9367
rect 7748 9324 7800 9333
rect 8116 9324 8168 9376
rect 8300 9324 8352 9376
rect 12900 9528 12952 9580
rect 11796 9503 11848 9512
rect 11796 9469 11805 9503
rect 11805 9469 11839 9503
rect 11839 9469 11848 9503
rect 11796 9460 11848 9469
rect 12256 9460 12308 9512
rect 13452 9460 13504 9512
rect 15200 9460 15252 9512
rect 16028 9528 16080 9580
rect 16120 9460 16172 9512
rect 10968 9392 11020 9444
rect 11336 9324 11388 9376
rect 13084 9392 13136 9444
rect 14096 9392 14148 9444
rect 14188 9324 14240 9376
rect 15292 9324 15344 9376
rect 18420 9460 18472 9512
rect 19616 9503 19668 9512
rect 19616 9469 19625 9503
rect 19625 9469 19659 9503
rect 19659 9469 19668 9503
rect 19616 9460 19668 9469
rect 20536 9392 20588 9444
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 22744 9664 22796 9716
rect 23020 9664 23072 9716
rect 24860 9664 24912 9716
rect 25044 9664 25096 9716
rect 25504 9664 25556 9716
rect 23572 9596 23624 9648
rect 22560 9503 22612 9512
rect 22560 9469 22569 9503
rect 22569 9469 22603 9503
rect 22603 9469 22612 9503
rect 22560 9460 22612 9469
rect 22836 9460 22888 9512
rect 17868 9324 17920 9376
rect 22928 9324 22980 9376
rect 24860 9571 24912 9580
rect 24860 9537 24869 9571
rect 24869 9537 24903 9571
rect 24903 9537 24912 9571
rect 24860 9528 24912 9537
rect 24308 9367 24360 9376
rect 24308 9333 24317 9367
rect 24317 9333 24351 9367
rect 24351 9333 24360 9367
rect 24308 9324 24360 9333
rect 25872 9503 25924 9512
rect 25872 9469 25881 9503
rect 25881 9469 25915 9503
rect 25915 9469 25924 9503
rect 25872 9460 25924 9469
rect 24952 9324 25004 9376
rect 4124 9222 4176 9274
rect 4188 9222 4240 9274
rect 4252 9222 4304 9274
rect 4316 9222 4368 9274
rect 4380 9222 4432 9274
rect 10472 9222 10524 9274
rect 10536 9222 10588 9274
rect 10600 9222 10652 9274
rect 10664 9222 10716 9274
rect 10728 9222 10780 9274
rect 16820 9222 16872 9274
rect 16884 9222 16936 9274
rect 16948 9222 17000 9274
rect 17012 9222 17064 9274
rect 17076 9222 17128 9274
rect 23168 9222 23220 9274
rect 23232 9222 23284 9274
rect 23296 9222 23348 9274
rect 23360 9222 23412 9274
rect 23424 9222 23476 9274
rect 5908 9120 5960 9172
rect 4160 8984 4212 9036
rect 3516 8959 3568 8968
rect 3516 8925 3525 8959
rect 3525 8925 3559 8959
rect 3559 8925 3568 8959
rect 3516 8916 3568 8925
rect 4068 8916 4120 8968
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 7012 8984 7064 9036
rect 8208 9120 8260 9172
rect 9680 9120 9732 9172
rect 12808 9120 12860 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 18420 9120 18472 9172
rect 22008 9120 22060 9172
rect 23020 9120 23072 9172
rect 6184 8891 6236 8900
rect 6184 8857 6193 8891
rect 6193 8857 6227 8891
rect 6227 8857 6236 8891
rect 6184 8848 6236 8857
rect 6552 8916 6604 8968
rect 6920 8916 6972 8968
rect 8208 8984 8260 9036
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 8024 8916 8076 8968
rect 2872 8780 2924 8832
rect 3700 8780 3752 8832
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 4712 8780 4764 8832
rect 6828 8780 6880 8832
rect 8300 8848 8352 8900
rect 10968 8916 11020 8968
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 11428 9052 11480 9104
rect 13084 9052 13136 9104
rect 11336 8984 11388 9036
rect 11888 8984 11940 9036
rect 15108 9052 15160 9104
rect 24860 9120 24912 9172
rect 14188 9027 14240 9036
rect 14188 8993 14197 9027
rect 14197 8993 14231 9027
rect 14231 8993 14240 9027
rect 14188 8984 14240 8993
rect 14280 8984 14332 9036
rect 16120 9027 16172 9036
rect 16120 8993 16129 9027
rect 16129 8993 16163 9027
rect 16163 8993 16172 9027
rect 16120 8984 16172 8993
rect 11704 8916 11756 8968
rect 12808 8916 12860 8968
rect 20536 8984 20588 9036
rect 23480 8984 23532 9036
rect 23940 9027 23992 9036
rect 23940 8993 23949 9027
rect 23949 8993 23983 9027
rect 23983 8993 23992 9027
rect 23940 8984 23992 8993
rect 24308 8984 24360 9036
rect 25320 8984 25372 9036
rect 17960 8916 18012 8968
rect 18880 8916 18932 8968
rect 10048 8848 10100 8900
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 12164 8848 12216 8900
rect 13084 8848 13136 8900
rect 17868 8891 17920 8900
rect 17868 8857 17877 8891
rect 17877 8857 17911 8891
rect 17911 8857 17920 8891
rect 17868 8848 17920 8857
rect 20628 8916 20680 8968
rect 20720 8959 20772 8968
rect 20720 8925 20729 8959
rect 20729 8925 20763 8959
rect 20763 8925 20772 8959
rect 20720 8916 20772 8925
rect 22836 8916 22888 8968
rect 23572 8916 23624 8968
rect 23664 8959 23716 8968
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 23756 8916 23808 8968
rect 21548 8848 21600 8900
rect 11612 8780 11664 8832
rect 11980 8780 12032 8832
rect 12532 8780 12584 8832
rect 12716 8823 12768 8832
rect 12716 8789 12725 8823
rect 12725 8789 12759 8823
rect 12759 8789 12768 8823
rect 12716 8780 12768 8789
rect 12900 8780 12952 8832
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 15936 8823 15988 8832
rect 15936 8789 15945 8823
rect 15945 8789 15979 8823
rect 15979 8789 15988 8823
rect 15936 8780 15988 8789
rect 17408 8780 17460 8832
rect 20444 8780 20496 8832
rect 23204 8780 23256 8832
rect 23848 8848 23900 8900
rect 24032 8848 24084 8900
rect 24676 8848 24728 8900
rect 23572 8780 23624 8832
rect 24308 8780 24360 8832
rect 24952 8780 25004 8832
rect 7298 8678 7350 8730
rect 7362 8678 7414 8730
rect 7426 8678 7478 8730
rect 7490 8678 7542 8730
rect 7554 8678 7606 8730
rect 13646 8678 13698 8730
rect 13710 8678 13762 8730
rect 13774 8678 13826 8730
rect 13838 8678 13890 8730
rect 13902 8678 13954 8730
rect 19994 8678 20046 8730
rect 20058 8678 20110 8730
rect 20122 8678 20174 8730
rect 20186 8678 20238 8730
rect 20250 8678 20302 8730
rect 26342 8678 26394 8730
rect 26406 8678 26458 8730
rect 26470 8678 26522 8730
rect 26534 8678 26586 8730
rect 26598 8678 26650 8730
rect 3884 8576 3936 8628
rect 4528 8576 4580 8628
rect 8024 8576 8076 8628
rect 9496 8576 9548 8628
rect 10232 8576 10284 8628
rect 10876 8576 10928 8628
rect 11428 8576 11480 8628
rect 4068 8551 4120 8560
rect 4068 8517 4103 8551
rect 4103 8517 4120 8551
rect 4068 8508 4120 8517
rect 5540 8508 5592 8560
rect 8116 8508 8168 8560
rect 9404 8508 9456 8560
rect 3424 8440 3476 8492
rect 3516 8440 3568 8492
rect 3608 8440 3660 8492
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 3700 8304 3752 8356
rect 5908 8440 5960 8492
rect 6828 8440 6880 8492
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 7932 8440 7984 8492
rect 4528 8372 4580 8424
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 11612 8551 11664 8560
rect 11612 8517 11621 8551
rect 11621 8517 11655 8551
rect 11655 8517 11664 8551
rect 11612 8508 11664 8517
rect 11796 8576 11848 8628
rect 13268 8619 13320 8628
rect 13268 8585 13277 8619
rect 13277 8585 13311 8619
rect 13311 8585 13320 8619
rect 13268 8576 13320 8585
rect 14924 8619 14976 8628
rect 14924 8585 14933 8619
rect 14933 8585 14967 8619
rect 14967 8585 14976 8619
rect 14924 8576 14976 8585
rect 15384 8576 15436 8628
rect 11060 8372 11112 8424
rect 1860 8236 1912 8288
rect 3332 8236 3384 8288
rect 7288 8236 7340 8288
rect 8760 8236 8812 8288
rect 11152 8304 11204 8356
rect 11520 8372 11572 8424
rect 12072 8440 12124 8492
rect 12716 8508 12768 8560
rect 15936 8576 15988 8628
rect 20352 8576 20404 8628
rect 20628 8576 20680 8628
rect 22560 8576 22612 8628
rect 23756 8576 23808 8628
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 11980 8372 12032 8424
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 16028 8551 16080 8560
rect 16028 8517 16037 8551
rect 16037 8517 16071 8551
rect 16071 8517 16080 8551
rect 16028 8508 16080 8517
rect 20720 8508 20772 8560
rect 23480 8508 23532 8560
rect 24032 8576 24084 8628
rect 25872 8576 25924 8628
rect 12256 8304 12308 8356
rect 12716 8304 12768 8356
rect 17776 8372 17828 8424
rect 19708 8415 19760 8424
rect 19708 8381 19717 8415
rect 19717 8381 19751 8415
rect 19751 8381 19760 8415
rect 19708 8372 19760 8381
rect 20352 8483 20404 8492
rect 20352 8449 20361 8483
rect 20361 8449 20395 8483
rect 20395 8449 20404 8483
rect 20352 8440 20404 8449
rect 21272 8372 21324 8424
rect 22376 8415 22428 8424
rect 22376 8381 22385 8415
rect 22385 8381 22419 8415
rect 22419 8381 22428 8415
rect 22376 8372 22428 8381
rect 23020 8440 23072 8492
rect 23204 8483 23256 8492
rect 23204 8449 23213 8483
rect 23213 8449 23247 8483
rect 23247 8449 23256 8483
rect 24400 8508 24452 8560
rect 24676 8508 24728 8560
rect 23204 8440 23256 8449
rect 23572 8372 23624 8424
rect 23756 8372 23808 8424
rect 16120 8304 16172 8356
rect 19892 8347 19944 8356
rect 19892 8313 19901 8347
rect 19901 8313 19935 8347
rect 19935 8313 19944 8347
rect 19892 8304 19944 8313
rect 20812 8304 20864 8356
rect 22928 8304 22980 8356
rect 24584 8372 24636 8424
rect 24860 8372 24912 8424
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 15292 8236 15344 8288
rect 16212 8279 16264 8288
rect 16212 8245 16221 8279
rect 16221 8245 16255 8279
rect 16255 8245 16264 8279
rect 16212 8236 16264 8245
rect 16396 8236 16448 8288
rect 18328 8236 18380 8288
rect 23664 8236 23716 8288
rect 25780 8304 25832 8356
rect 4124 8134 4176 8186
rect 4188 8134 4240 8186
rect 4252 8134 4304 8186
rect 4316 8134 4368 8186
rect 4380 8134 4432 8186
rect 10472 8134 10524 8186
rect 10536 8134 10588 8186
rect 10600 8134 10652 8186
rect 10664 8134 10716 8186
rect 10728 8134 10780 8186
rect 16820 8134 16872 8186
rect 16884 8134 16936 8186
rect 16948 8134 17000 8186
rect 17012 8134 17064 8186
rect 17076 8134 17128 8186
rect 23168 8134 23220 8186
rect 23232 8134 23284 8186
rect 23296 8134 23348 8186
rect 23360 8134 23412 8186
rect 23424 8134 23476 8186
rect 3976 8075 4028 8084
rect 3976 8041 3985 8075
rect 3985 8041 4019 8075
rect 4019 8041 4028 8075
rect 3976 8032 4028 8041
rect 4068 8032 4120 8084
rect 14004 8032 14056 8084
rect 4528 7964 4580 8016
rect 10048 8007 10100 8016
rect 10048 7973 10057 8007
rect 10057 7973 10091 8007
rect 10091 7973 10100 8007
rect 10048 7964 10100 7973
rect 12164 7964 12216 8016
rect 2872 7896 2924 7948
rect 5448 7896 5500 7948
rect 6552 7896 6604 7948
rect 7104 7896 7156 7948
rect 8300 7896 8352 7948
rect 8760 7939 8812 7948
rect 8760 7905 8769 7939
rect 8769 7905 8803 7939
rect 8803 7905 8812 7939
rect 8760 7896 8812 7905
rect 10876 7896 10928 7948
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 2780 7760 2832 7812
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4528 7828 4580 7880
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 11980 7828 12032 7880
rect 6920 7760 6972 7812
rect 7288 7760 7340 7812
rect 7656 7760 7708 7812
rect 11520 7760 11572 7812
rect 13176 7964 13228 8016
rect 13452 7896 13504 7948
rect 15200 7896 15252 7948
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 16212 8032 16264 8084
rect 23020 8032 23072 8084
rect 23572 8075 23624 8084
rect 23572 8041 23581 8075
rect 23581 8041 23615 8075
rect 23615 8041 23624 8075
rect 23572 8032 23624 8041
rect 19524 7964 19576 8016
rect 19892 7939 19944 7948
rect 17316 7828 17368 7880
rect 18880 7828 18932 7880
rect 19892 7905 19901 7939
rect 19901 7905 19935 7939
rect 19935 7905 19944 7939
rect 19892 7896 19944 7905
rect 20628 7939 20680 7948
rect 20628 7905 20637 7939
rect 20637 7905 20671 7939
rect 20671 7905 20680 7939
rect 20628 7896 20680 7905
rect 22560 7896 22612 7948
rect 15660 7760 15712 7812
rect 4620 7692 4672 7744
rect 7196 7692 7248 7744
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 12256 7692 12308 7744
rect 14556 7735 14608 7744
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 16488 7692 16540 7744
rect 18696 7760 18748 7812
rect 19800 7828 19852 7880
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 20812 7760 20864 7812
rect 21180 7760 21232 7812
rect 23388 7871 23440 7880
rect 23388 7837 23397 7871
rect 23397 7837 23431 7871
rect 23431 7837 23440 7871
rect 23388 7828 23440 7837
rect 17408 7692 17460 7744
rect 17684 7692 17736 7744
rect 19340 7692 19392 7744
rect 20536 7735 20588 7744
rect 20536 7701 20545 7735
rect 20545 7701 20579 7735
rect 20579 7701 20588 7735
rect 20536 7692 20588 7701
rect 20720 7692 20772 7744
rect 22192 7692 22244 7744
rect 22376 7735 22428 7744
rect 22376 7701 22385 7735
rect 22385 7701 22419 7735
rect 22419 7701 22428 7735
rect 22376 7692 22428 7701
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 23940 7871 23992 7880
rect 23940 7837 23949 7871
rect 23949 7837 23983 7871
rect 23983 7837 23992 7871
rect 23940 7828 23992 7837
rect 24032 7760 24084 7812
rect 23848 7692 23900 7744
rect 24216 7692 24268 7744
rect 7298 7590 7350 7642
rect 7362 7590 7414 7642
rect 7426 7590 7478 7642
rect 7490 7590 7542 7642
rect 7554 7590 7606 7642
rect 13646 7590 13698 7642
rect 13710 7590 13762 7642
rect 13774 7590 13826 7642
rect 13838 7590 13890 7642
rect 13902 7590 13954 7642
rect 19994 7590 20046 7642
rect 20058 7590 20110 7642
rect 20122 7590 20174 7642
rect 20186 7590 20238 7642
rect 20250 7590 20302 7642
rect 26342 7590 26394 7642
rect 26406 7590 26458 7642
rect 26470 7590 26522 7642
rect 26534 7590 26586 7642
rect 26598 7590 26650 7642
rect 1676 7488 1728 7540
rect 3792 7488 3844 7540
rect 3884 7463 3936 7472
rect 3884 7429 3893 7463
rect 3893 7429 3927 7463
rect 3927 7429 3936 7463
rect 3884 7420 3936 7429
rect 3516 7352 3568 7404
rect 7104 7488 7156 7540
rect 9680 7488 9732 7540
rect 12072 7488 12124 7540
rect 4712 7420 4764 7472
rect 6920 7420 6972 7472
rect 9772 7420 9824 7472
rect 12808 7488 12860 7540
rect 5908 7352 5960 7404
rect 12716 7463 12768 7472
rect 12716 7429 12725 7463
rect 12725 7429 12759 7463
rect 12759 7429 12768 7463
rect 12716 7420 12768 7429
rect 14556 7488 14608 7540
rect 16028 7488 16080 7540
rect 19524 7488 19576 7540
rect 19892 7488 19944 7540
rect 20352 7531 20404 7540
rect 20352 7497 20361 7531
rect 20361 7497 20395 7531
rect 20395 7497 20404 7531
rect 20352 7488 20404 7497
rect 20536 7488 20588 7540
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 21272 7488 21324 7540
rect 16488 7420 16540 7472
rect 18696 7420 18748 7472
rect 3332 7327 3384 7336
rect 3332 7293 3341 7327
rect 3341 7293 3375 7327
rect 3375 7293 3384 7327
rect 3332 7284 3384 7293
rect 4896 7284 4948 7336
rect 5172 7284 5224 7336
rect 10048 7327 10100 7336
rect 10048 7293 10057 7327
rect 10057 7293 10091 7327
rect 10091 7293 10100 7327
rect 10048 7284 10100 7293
rect 16120 7352 16172 7404
rect 11520 7216 11572 7268
rect 2780 7148 2832 7200
rect 4988 7148 5040 7200
rect 7932 7148 7984 7200
rect 9496 7148 9548 7200
rect 11612 7191 11664 7200
rect 11612 7157 11621 7191
rect 11621 7157 11655 7191
rect 11655 7157 11664 7191
rect 11612 7148 11664 7157
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 16028 7284 16080 7336
rect 17316 7284 17368 7336
rect 17868 7327 17920 7336
rect 17868 7293 17877 7327
rect 17877 7293 17911 7327
rect 17911 7293 17920 7327
rect 17868 7284 17920 7293
rect 17776 7259 17828 7268
rect 17776 7225 17785 7259
rect 17785 7225 17819 7259
rect 17819 7225 17828 7259
rect 17776 7216 17828 7225
rect 12900 7148 12952 7200
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 17592 7191 17644 7200
rect 17592 7157 17601 7191
rect 17601 7157 17635 7191
rect 17635 7157 17644 7191
rect 17592 7148 17644 7157
rect 18880 7148 18932 7200
rect 20812 7216 20864 7268
rect 21824 7352 21876 7404
rect 23388 7488 23440 7540
rect 24216 7488 24268 7540
rect 24308 7531 24360 7540
rect 24308 7497 24317 7531
rect 24317 7497 24351 7531
rect 24351 7497 24360 7531
rect 24308 7488 24360 7497
rect 24584 7488 24636 7540
rect 22652 7352 22704 7404
rect 22376 7284 22428 7336
rect 23020 7352 23072 7404
rect 22284 7216 22336 7268
rect 23848 7395 23900 7404
rect 23848 7361 23857 7395
rect 23857 7361 23891 7395
rect 23891 7361 23900 7395
rect 23848 7352 23900 7361
rect 21548 7191 21600 7200
rect 21548 7157 21557 7191
rect 21557 7157 21591 7191
rect 21591 7157 21600 7191
rect 21548 7148 21600 7157
rect 24492 7352 24544 7404
rect 25044 7395 25096 7404
rect 25044 7361 25053 7395
rect 25053 7361 25087 7395
rect 25087 7361 25096 7395
rect 25044 7352 25096 7361
rect 25228 7395 25280 7404
rect 25228 7361 25237 7395
rect 25237 7361 25271 7395
rect 25271 7361 25280 7395
rect 25228 7352 25280 7361
rect 24400 7148 24452 7200
rect 24860 7191 24912 7200
rect 24860 7157 24869 7191
rect 24869 7157 24903 7191
rect 24903 7157 24912 7191
rect 24860 7148 24912 7157
rect 24952 7148 25004 7200
rect 4124 7046 4176 7098
rect 4188 7046 4240 7098
rect 4252 7046 4304 7098
rect 4316 7046 4368 7098
rect 4380 7046 4432 7098
rect 10472 7046 10524 7098
rect 10536 7046 10588 7098
rect 10600 7046 10652 7098
rect 10664 7046 10716 7098
rect 10728 7046 10780 7098
rect 16820 7046 16872 7098
rect 16884 7046 16936 7098
rect 16948 7046 17000 7098
rect 17012 7046 17064 7098
rect 17076 7046 17128 7098
rect 23168 7046 23220 7098
rect 23232 7046 23284 7098
rect 23296 7046 23348 7098
rect 23360 7046 23412 7098
rect 23424 7046 23476 7098
rect 4344 6944 4396 6996
rect 3792 6919 3844 6928
rect 3792 6885 3801 6919
rect 3801 6885 3835 6919
rect 3835 6885 3844 6919
rect 3792 6876 3844 6885
rect 3424 6808 3476 6860
rect 3516 6808 3568 6860
rect 3148 6740 3200 6792
rect 4712 6783 4764 6792
rect 4712 6749 4722 6783
rect 4722 6749 4764 6783
rect 3608 6715 3660 6724
rect 3608 6681 3617 6715
rect 3617 6681 3651 6715
rect 3651 6681 3660 6715
rect 3608 6672 3660 6681
rect 3884 6672 3936 6724
rect 3976 6672 4028 6724
rect 4712 6740 4764 6749
rect 11152 6944 11204 6996
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 16028 6944 16080 6996
rect 17592 6944 17644 6996
rect 7932 6808 7984 6860
rect 15200 6876 15252 6928
rect 16396 6876 16448 6928
rect 23572 6944 23624 6996
rect 23940 6944 23992 6996
rect 24032 6944 24084 6996
rect 25044 6944 25096 6996
rect 26056 6944 26108 6996
rect 6000 6672 6052 6724
rect 4068 6604 4120 6656
rect 4344 6604 4396 6656
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 10232 6851 10284 6860
rect 10232 6817 10241 6851
rect 10241 6817 10275 6851
rect 10275 6817 10284 6851
rect 10232 6808 10284 6817
rect 11520 6808 11572 6860
rect 12440 6808 12492 6860
rect 14188 6808 14240 6860
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 10048 6740 10100 6792
rect 19708 6808 19760 6860
rect 24768 6808 24820 6860
rect 16580 6740 16632 6792
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 18696 6740 18748 6792
rect 19340 6740 19392 6792
rect 9036 6604 9088 6656
rect 9680 6604 9732 6656
rect 12348 6715 12400 6724
rect 12348 6681 12357 6715
rect 12357 6681 12391 6715
rect 12391 6681 12400 6715
rect 12348 6672 12400 6681
rect 12900 6672 12952 6724
rect 15844 6715 15896 6724
rect 15844 6681 15853 6715
rect 15853 6681 15887 6715
rect 15887 6681 15896 6715
rect 15844 6672 15896 6681
rect 17684 6672 17736 6724
rect 19800 6672 19852 6724
rect 23480 6740 23532 6792
rect 23756 6740 23808 6792
rect 23848 6740 23900 6792
rect 24308 6740 24360 6792
rect 11796 6604 11848 6656
rect 14004 6604 14056 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14464 6647 14516 6656
rect 14464 6613 14473 6647
rect 14473 6613 14507 6647
rect 14507 6613 14516 6647
rect 14464 6604 14516 6613
rect 19432 6647 19484 6656
rect 19432 6613 19441 6647
rect 19441 6613 19475 6647
rect 19475 6613 19484 6647
rect 19432 6604 19484 6613
rect 24676 6715 24728 6724
rect 24676 6681 24685 6715
rect 24685 6681 24719 6715
rect 24719 6681 24728 6715
rect 24676 6672 24728 6681
rect 25688 6672 25740 6724
rect 21732 6647 21784 6656
rect 21732 6613 21741 6647
rect 21741 6613 21775 6647
rect 21775 6613 21784 6647
rect 21732 6604 21784 6613
rect 22836 6647 22888 6656
rect 22836 6613 22845 6647
rect 22845 6613 22879 6647
rect 22879 6613 22888 6647
rect 22836 6604 22888 6613
rect 23664 6604 23716 6656
rect 7298 6502 7350 6554
rect 7362 6502 7414 6554
rect 7426 6502 7478 6554
rect 7490 6502 7542 6554
rect 7554 6502 7606 6554
rect 13646 6502 13698 6554
rect 13710 6502 13762 6554
rect 13774 6502 13826 6554
rect 13838 6502 13890 6554
rect 13902 6502 13954 6554
rect 19994 6502 20046 6554
rect 20058 6502 20110 6554
rect 20122 6502 20174 6554
rect 20186 6502 20238 6554
rect 20250 6502 20302 6554
rect 26342 6502 26394 6554
rect 26406 6502 26458 6554
rect 26470 6502 26522 6554
rect 26534 6502 26586 6554
rect 26598 6502 26650 6554
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 3516 6400 3568 6452
rect 3792 6400 3844 6452
rect 3884 6400 3936 6452
rect 2780 6264 2832 6316
rect 3608 6264 3660 6316
rect 3976 6332 4028 6384
rect 4804 6400 4856 6452
rect 4620 6332 4672 6384
rect 4896 6332 4948 6384
rect 4988 6375 5040 6384
rect 4988 6341 4997 6375
rect 4997 6341 5031 6375
rect 5031 6341 5040 6375
rect 4988 6332 5040 6341
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 4528 6196 4580 6248
rect 3700 6128 3752 6180
rect 5632 6264 5684 6316
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 8116 6400 8168 6452
rect 8208 6400 8260 6452
rect 10876 6400 10928 6452
rect 11152 6443 11204 6452
rect 11152 6409 11161 6443
rect 11161 6409 11195 6443
rect 11195 6409 11204 6443
rect 11152 6400 11204 6409
rect 11612 6400 11664 6452
rect 11796 6400 11848 6452
rect 14004 6400 14056 6452
rect 14464 6400 14516 6452
rect 18880 6443 18932 6452
rect 18880 6409 18889 6443
rect 18889 6409 18923 6443
rect 18923 6409 18932 6443
rect 18880 6400 18932 6409
rect 19340 6400 19392 6452
rect 4804 6128 4856 6180
rect 5356 6128 5408 6180
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 7932 6196 7984 6248
rect 9680 6332 9732 6384
rect 11520 6307 11572 6316
rect 11520 6273 11529 6307
rect 11529 6273 11563 6307
rect 11563 6273 11572 6307
rect 11520 6264 11572 6273
rect 19616 6400 19668 6452
rect 20628 6400 20680 6452
rect 19800 6332 19852 6384
rect 21732 6400 21784 6452
rect 21824 6443 21876 6452
rect 21824 6409 21833 6443
rect 21833 6409 21867 6443
rect 21867 6409 21876 6443
rect 21824 6400 21876 6409
rect 22560 6443 22612 6452
rect 22560 6409 22569 6443
rect 22569 6409 22603 6443
rect 22603 6409 22612 6443
rect 22560 6400 22612 6409
rect 22836 6400 22888 6452
rect 23848 6400 23900 6452
rect 24676 6400 24728 6452
rect 21180 6264 21232 6316
rect 5816 6060 5868 6112
rect 5908 6060 5960 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 8116 6060 8168 6112
rect 8576 6060 8628 6112
rect 8760 6060 8812 6112
rect 10232 6060 10284 6112
rect 12808 6060 12860 6112
rect 17408 6196 17460 6248
rect 19432 6128 19484 6180
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 15200 6060 15252 6112
rect 22192 6264 22244 6316
rect 21732 6196 21784 6248
rect 22836 6307 22888 6316
rect 22836 6273 22845 6307
rect 22845 6273 22879 6307
rect 22879 6273 22888 6307
rect 22836 6264 22888 6273
rect 21732 6060 21784 6112
rect 22560 6060 22612 6112
rect 22928 6196 22980 6248
rect 23572 6264 23624 6316
rect 24308 6332 24360 6384
rect 24584 6375 24636 6384
rect 24584 6341 24593 6375
rect 24593 6341 24627 6375
rect 24627 6341 24636 6375
rect 24584 6332 24636 6341
rect 24400 6307 24452 6316
rect 24400 6273 24409 6307
rect 24409 6273 24443 6307
rect 24443 6273 24452 6307
rect 24400 6264 24452 6273
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 25136 6239 25188 6248
rect 25136 6205 25145 6239
rect 25145 6205 25179 6239
rect 25179 6205 25188 6239
rect 25136 6196 25188 6205
rect 23020 6128 23072 6180
rect 26056 6307 26108 6316
rect 26056 6273 26065 6307
rect 26065 6273 26099 6307
rect 26099 6273 26108 6307
rect 26056 6264 26108 6273
rect 22928 6060 22980 6112
rect 23480 6103 23532 6112
rect 23480 6069 23489 6103
rect 23489 6069 23523 6103
rect 23523 6069 23532 6103
rect 23480 6060 23532 6069
rect 4124 5958 4176 6010
rect 4188 5958 4240 6010
rect 4252 5958 4304 6010
rect 4316 5958 4368 6010
rect 4380 5958 4432 6010
rect 10472 5958 10524 6010
rect 10536 5958 10588 6010
rect 10600 5958 10652 6010
rect 10664 5958 10716 6010
rect 10728 5958 10780 6010
rect 16820 5958 16872 6010
rect 16884 5958 16936 6010
rect 16948 5958 17000 6010
rect 17012 5958 17064 6010
rect 17076 5958 17128 6010
rect 23168 5958 23220 6010
rect 23232 5958 23284 6010
rect 23296 5958 23348 6010
rect 23360 5958 23412 6010
rect 23424 5958 23476 6010
rect 3148 5856 3200 5908
rect 3608 5856 3660 5908
rect 4436 5856 4488 5908
rect 4804 5856 4856 5908
rect 4896 5856 4948 5908
rect 5540 5856 5592 5908
rect 5632 5856 5684 5908
rect 6552 5856 6604 5908
rect 8668 5856 8720 5908
rect 9036 5856 9088 5908
rect 9220 5856 9272 5908
rect 11796 5856 11848 5908
rect 3240 5627 3292 5636
rect 3240 5593 3249 5627
rect 3249 5593 3283 5627
rect 3283 5593 3292 5627
rect 3240 5584 3292 5593
rect 3884 5652 3936 5704
rect 4804 5652 4856 5704
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 6920 5720 6972 5772
rect 8116 5720 8168 5772
rect 3608 5559 3660 5568
rect 3608 5525 3617 5559
rect 3617 5525 3651 5559
rect 3651 5525 3660 5559
rect 3608 5516 3660 5525
rect 3700 5516 3752 5568
rect 4068 5516 4120 5568
rect 6460 5584 6512 5636
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 10324 5652 10376 5704
rect 13360 5856 13412 5908
rect 14096 5856 14148 5908
rect 21732 5899 21784 5908
rect 21732 5865 21741 5899
rect 21741 5865 21775 5899
rect 21775 5865 21784 5899
rect 21732 5856 21784 5865
rect 22744 5899 22796 5908
rect 22744 5865 22753 5899
rect 22753 5865 22787 5899
rect 22787 5865 22796 5899
rect 22744 5856 22796 5865
rect 22836 5856 22888 5908
rect 22928 5856 22980 5908
rect 25228 5856 25280 5908
rect 12716 5788 12768 5840
rect 13084 5652 13136 5704
rect 14648 5831 14700 5840
rect 14648 5797 14657 5831
rect 14657 5797 14691 5831
rect 14691 5797 14700 5831
rect 14648 5788 14700 5797
rect 16580 5720 16632 5772
rect 19616 5763 19668 5772
rect 19616 5729 19625 5763
rect 19625 5729 19659 5763
rect 19659 5729 19668 5763
rect 19616 5720 19668 5729
rect 12348 5584 12400 5636
rect 17316 5652 17368 5704
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 21640 5788 21692 5840
rect 7104 5516 7156 5568
rect 13176 5516 13228 5568
rect 14464 5516 14516 5568
rect 15292 5516 15344 5568
rect 15568 5516 15620 5568
rect 16488 5584 16540 5636
rect 16948 5627 17000 5636
rect 16948 5593 16957 5627
rect 16957 5593 16991 5627
rect 16991 5593 17000 5627
rect 16948 5584 17000 5593
rect 19892 5627 19944 5636
rect 19892 5593 19901 5627
rect 19901 5593 19935 5627
rect 19935 5593 19944 5627
rect 19892 5584 19944 5593
rect 21180 5584 21232 5636
rect 17868 5516 17920 5568
rect 22836 5584 22888 5636
rect 23020 5652 23072 5704
rect 24952 5720 25004 5772
rect 25044 5695 25096 5704
rect 25044 5661 25053 5695
rect 25053 5661 25087 5695
rect 25087 5661 25096 5695
rect 25044 5652 25096 5661
rect 21916 5516 21968 5568
rect 22652 5516 22704 5568
rect 23204 5516 23256 5568
rect 7298 5414 7350 5466
rect 7362 5414 7414 5466
rect 7426 5414 7478 5466
rect 7490 5414 7542 5466
rect 7554 5414 7606 5466
rect 13646 5414 13698 5466
rect 13710 5414 13762 5466
rect 13774 5414 13826 5466
rect 13838 5414 13890 5466
rect 13902 5414 13954 5466
rect 19994 5414 20046 5466
rect 20058 5414 20110 5466
rect 20122 5414 20174 5466
rect 20186 5414 20238 5466
rect 20250 5414 20302 5466
rect 26342 5414 26394 5466
rect 26406 5414 26458 5466
rect 26470 5414 26522 5466
rect 26534 5414 26586 5466
rect 26598 5414 26650 5466
rect 3516 5312 3568 5364
rect 4896 5312 4948 5364
rect 5724 5312 5776 5364
rect 9496 5312 9548 5364
rect 9680 5312 9732 5364
rect 15108 5312 15160 5364
rect 3240 5244 3292 5296
rect 4068 5244 4120 5296
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 3700 5176 3752 5228
rect 2872 5108 2924 5160
rect 3976 5108 4028 5160
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 8392 5244 8444 5296
rect 11980 5244 12032 5296
rect 9680 5176 9732 5228
rect 5172 5108 5224 5160
rect 5908 5108 5960 5160
rect 4712 5040 4764 5092
rect 12808 5176 12860 5228
rect 13452 5040 13504 5092
rect 13544 5040 13596 5092
rect 14372 5176 14424 5228
rect 15384 5219 15436 5228
rect 15384 5185 15393 5219
rect 15393 5185 15427 5219
rect 15427 5185 15436 5219
rect 15384 5176 15436 5185
rect 16580 5312 16632 5364
rect 16948 5312 17000 5364
rect 19892 5312 19944 5364
rect 21548 5312 21600 5364
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 16396 5244 16448 5296
rect 17592 5287 17644 5296
rect 17592 5253 17601 5287
rect 17601 5253 17635 5287
rect 17635 5253 17644 5287
rect 17592 5244 17644 5253
rect 15844 5176 15896 5228
rect 17224 5176 17276 5228
rect 18696 5176 18748 5228
rect 22744 5312 22796 5364
rect 23204 5312 23256 5364
rect 23572 5312 23624 5364
rect 22468 5244 22520 5296
rect 22652 5244 22704 5296
rect 22008 5219 22060 5228
rect 22008 5185 22017 5219
rect 22017 5185 22051 5219
rect 22051 5185 22060 5219
rect 22008 5176 22060 5185
rect 22284 5219 22336 5228
rect 22284 5185 22319 5219
rect 22319 5185 22336 5219
rect 22284 5176 22336 5185
rect 22744 5219 22796 5228
rect 22744 5185 22753 5219
rect 22753 5185 22787 5219
rect 22787 5185 22796 5219
rect 22744 5176 22796 5185
rect 22928 5219 22980 5228
rect 22928 5185 22937 5219
rect 22937 5185 22971 5219
rect 22971 5185 22980 5219
rect 22928 5176 22980 5185
rect 24216 5287 24268 5296
rect 24216 5253 24225 5287
rect 24225 5253 24259 5287
rect 24259 5253 24268 5287
rect 25136 5312 25188 5364
rect 25412 5312 25464 5364
rect 24216 5244 24268 5253
rect 25228 5244 25280 5296
rect 23664 5176 23716 5228
rect 16396 5108 16448 5160
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 17316 5108 17368 5117
rect 3884 4972 3936 5024
rect 4804 4972 4856 5024
rect 5540 4972 5592 5024
rect 5908 4972 5960 5024
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 13360 4972 13412 5024
rect 14648 5040 14700 5092
rect 15108 5040 15160 5092
rect 15292 5040 15344 5092
rect 18144 5108 18196 5160
rect 22192 5108 22244 5160
rect 14188 4972 14240 5024
rect 16120 4972 16172 5024
rect 17684 4972 17736 5024
rect 18236 4972 18288 5024
rect 19248 4972 19300 5024
rect 21272 4972 21324 5024
rect 23848 4972 23900 5024
rect 23940 5015 23992 5024
rect 23940 4981 23949 5015
rect 23949 4981 23983 5015
rect 23983 4981 23992 5015
rect 23940 4972 23992 4981
rect 26516 4972 26568 5024
rect 4124 4870 4176 4922
rect 4188 4870 4240 4922
rect 4252 4870 4304 4922
rect 4316 4870 4368 4922
rect 4380 4870 4432 4922
rect 10472 4870 10524 4922
rect 10536 4870 10588 4922
rect 10600 4870 10652 4922
rect 10664 4870 10716 4922
rect 10728 4870 10780 4922
rect 16820 4870 16872 4922
rect 16884 4870 16936 4922
rect 16948 4870 17000 4922
rect 17012 4870 17064 4922
rect 17076 4870 17128 4922
rect 23168 4870 23220 4922
rect 23232 4870 23284 4922
rect 23296 4870 23348 4922
rect 23360 4870 23412 4922
rect 23424 4870 23476 4922
rect 3608 4768 3660 4820
rect 3700 4768 3752 4820
rect 4804 4768 4856 4820
rect 5080 4768 5132 4820
rect 5816 4768 5868 4820
rect 9680 4811 9732 4820
rect 9680 4777 9689 4811
rect 9689 4777 9723 4811
rect 9723 4777 9732 4811
rect 9680 4768 9732 4777
rect 10048 4811 10100 4820
rect 10048 4777 10057 4811
rect 10057 4777 10091 4811
rect 10091 4777 10100 4811
rect 10048 4768 10100 4777
rect 12624 4768 12676 4820
rect 13268 4768 13320 4820
rect 14372 4768 14424 4820
rect 15384 4768 15436 4820
rect 3240 4700 3292 4752
rect 4712 4700 4764 4752
rect 3056 4632 3108 4684
rect 3792 4675 3844 4684
rect 3792 4641 3801 4675
rect 3801 4641 3835 4675
rect 3835 4641 3844 4675
rect 3792 4632 3844 4641
rect 4528 4564 4580 4616
rect 3884 4496 3936 4548
rect 4712 4496 4764 4548
rect 4436 4471 4488 4480
rect 4436 4437 4463 4471
rect 4463 4437 4488 4471
rect 4436 4428 4488 4437
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 5172 4539 5224 4548
rect 5172 4505 5181 4539
rect 5181 4505 5215 4539
rect 5215 4505 5224 4539
rect 5172 4496 5224 4505
rect 5632 4496 5684 4548
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 8208 4700 8260 4752
rect 7196 4632 7248 4684
rect 8392 4632 8444 4684
rect 8668 4675 8720 4684
rect 8668 4641 8677 4675
rect 8677 4641 8711 4675
rect 8711 4641 8720 4675
rect 8668 4632 8720 4641
rect 8852 4564 8904 4616
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 8208 4496 8260 4548
rect 13176 4700 13228 4752
rect 12992 4675 13044 4684
rect 12992 4641 13001 4675
rect 13001 4641 13035 4675
rect 13035 4641 13044 4675
rect 12992 4632 13044 4641
rect 13452 4700 13504 4752
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 13544 4564 13596 4616
rect 14004 4564 14056 4616
rect 15476 4700 15528 4752
rect 15752 4768 15804 4820
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 16120 4811 16172 4820
rect 16120 4777 16129 4811
rect 16129 4777 16163 4811
rect 16163 4777 16172 4811
rect 16120 4768 16172 4777
rect 16764 4768 16816 4820
rect 17224 4768 17276 4820
rect 17592 4768 17644 4820
rect 22008 4768 22060 4820
rect 10324 4496 10376 4548
rect 12992 4496 13044 4548
rect 13360 4496 13412 4548
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14648 4564 14700 4616
rect 14924 4564 14976 4616
rect 15292 4564 15344 4616
rect 14740 4496 14792 4548
rect 5540 4428 5592 4480
rect 5724 4428 5776 4480
rect 7656 4428 7708 4480
rect 8300 4428 8352 4480
rect 11796 4428 11848 4480
rect 13084 4428 13136 4480
rect 14004 4428 14056 4480
rect 14096 4428 14148 4480
rect 15016 4471 15068 4480
rect 15016 4437 15025 4471
rect 15025 4437 15059 4471
rect 15059 4437 15068 4471
rect 15016 4428 15068 4437
rect 15476 4539 15528 4548
rect 15476 4505 15485 4539
rect 15485 4505 15519 4539
rect 15519 4505 15528 4539
rect 16028 4607 16080 4616
rect 16028 4573 16037 4607
rect 16037 4573 16071 4607
rect 16071 4573 16080 4607
rect 16028 4564 16080 4573
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 16488 4564 16540 4616
rect 15476 4496 15528 4505
rect 16120 4496 16172 4548
rect 16672 4496 16724 4548
rect 15660 4471 15712 4480
rect 15660 4437 15690 4471
rect 15690 4437 15712 4471
rect 15660 4428 15712 4437
rect 15844 4428 15896 4480
rect 17132 4607 17184 4616
rect 17132 4573 17141 4607
rect 17141 4573 17175 4607
rect 17175 4573 17184 4607
rect 17132 4564 17184 4573
rect 17408 4564 17460 4616
rect 17500 4564 17552 4616
rect 18144 4607 18196 4616
rect 18144 4573 18153 4607
rect 18153 4573 18187 4607
rect 18187 4573 18196 4607
rect 18144 4564 18196 4573
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 17224 4496 17276 4548
rect 17592 4428 17644 4480
rect 17868 4428 17920 4480
rect 18512 4539 18564 4548
rect 18512 4505 18521 4539
rect 18521 4505 18555 4539
rect 18555 4505 18564 4539
rect 18512 4496 18564 4505
rect 18972 4564 19024 4616
rect 19340 4564 19392 4616
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20628 4675 20680 4684
rect 20628 4641 20637 4675
rect 20637 4641 20671 4675
rect 20671 4641 20680 4675
rect 20628 4632 20680 4641
rect 19800 4607 19852 4616
rect 19800 4573 19809 4607
rect 19809 4573 19843 4607
rect 19843 4573 19852 4607
rect 19800 4564 19852 4573
rect 22744 4609 22796 4616
rect 22744 4575 22753 4609
rect 22753 4575 22787 4609
rect 22787 4575 22796 4609
rect 22744 4564 22796 4575
rect 22928 4607 22980 4616
rect 22928 4573 22937 4607
rect 22937 4573 22971 4607
rect 22971 4573 22980 4607
rect 23572 4700 23624 4752
rect 22928 4564 22980 4573
rect 25228 4675 25280 4684
rect 25228 4641 25237 4675
rect 25237 4641 25271 4675
rect 25271 4641 25280 4675
rect 25228 4632 25280 4641
rect 20904 4539 20956 4548
rect 20904 4505 20913 4539
rect 20913 4505 20947 4539
rect 20947 4505 20956 4539
rect 20904 4496 20956 4505
rect 21916 4496 21968 4548
rect 23940 4564 23992 4616
rect 24492 4564 24544 4616
rect 23664 4496 23716 4548
rect 24216 4496 24268 4548
rect 18880 4471 18932 4480
rect 18880 4437 18889 4471
rect 18889 4437 18923 4471
rect 18923 4437 18932 4471
rect 18880 4428 18932 4437
rect 18972 4428 19024 4480
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 22284 4428 22336 4480
rect 22928 4428 22980 4480
rect 23020 4428 23072 4480
rect 23296 4428 23348 4480
rect 24584 4471 24636 4480
rect 24584 4437 24593 4471
rect 24593 4437 24627 4471
rect 24627 4437 24636 4471
rect 24584 4428 24636 4437
rect 24860 4428 24912 4480
rect 7298 4326 7350 4378
rect 7362 4326 7414 4378
rect 7426 4326 7478 4378
rect 7490 4326 7542 4378
rect 7554 4326 7606 4378
rect 13646 4326 13698 4378
rect 13710 4326 13762 4378
rect 13774 4326 13826 4378
rect 13838 4326 13890 4378
rect 13902 4326 13954 4378
rect 19994 4326 20046 4378
rect 20058 4326 20110 4378
rect 20122 4326 20174 4378
rect 20186 4326 20238 4378
rect 20250 4326 20302 4378
rect 26342 4326 26394 4378
rect 26406 4326 26458 4378
rect 26470 4326 26522 4378
rect 26534 4326 26586 4378
rect 26598 4326 26650 4378
rect 3056 4267 3108 4276
rect 3056 4233 3065 4267
rect 3065 4233 3099 4267
rect 3099 4233 3108 4267
rect 3056 4224 3108 4233
rect 5448 4224 5500 4276
rect 5540 4224 5592 4276
rect 6000 4224 6052 4276
rect 3976 4199 4028 4208
rect 3976 4165 4011 4199
rect 4011 4165 4028 4199
rect 3976 4156 4028 4165
rect 5816 4156 5868 4208
rect 6368 4267 6420 4276
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 7196 4224 7248 4276
rect 8944 4224 8996 4276
rect 10048 4224 10100 4276
rect 10232 4224 10284 4276
rect 13544 4224 13596 4276
rect 3516 4088 3568 4140
rect 3792 4131 3844 4140
rect 3792 4097 3802 4131
rect 3802 4097 3836 4131
rect 3836 4097 3844 4131
rect 3792 4088 3844 4097
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5448 4131 5500 4140
rect 5448 4097 5483 4131
rect 5483 4097 5500 4131
rect 5448 4088 5500 4097
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 3332 3952 3384 4004
rect 2688 3927 2740 3936
rect 2688 3893 2697 3927
rect 2697 3893 2731 3927
rect 2731 3893 2740 3927
rect 2688 3884 2740 3893
rect 3240 3884 3292 3936
rect 4436 3884 4488 3936
rect 4620 3884 4672 3936
rect 5080 4020 5132 4072
rect 5724 4020 5776 4072
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 6644 4156 6696 4208
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 13176 4156 13228 4208
rect 6092 3952 6144 4004
rect 8576 4020 8628 4072
rect 10324 4131 10376 4140
rect 10324 4097 10333 4131
rect 10333 4097 10367 4131
rect 10367 4097 10376 4131
rect 10324 4088 10376 4097
rect 10416 4088 10468 4140
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 13176 4020 13228 4072
rect 7932 3884 7984 3936
rect 8760 3884 8812 3936
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 10324 3884 10376 3936
rect 11428 3884 11480 3936
rect 13912 4156 13964 4208
rect 14004 4156 14056 4208
rect 14372 4199 14424 4208
rect 14372 4165 14389 4199
rect 14389 4165 14424 4199
rect 14372 4156 14424 4165
rect 14372 4020 14424 4072
rect 15660 4224 15712 4276
rect 16580 4224 16632 4276
rect 15016 4088 15068 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 16764 4088 16816 4140
rect 15936 4063 15988 4072
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 17408 4088 17460 4140
rect 17592 4131 17644 4140
rect 17592 4097 17601 4131
rect 17601 4097 17635 4131
rect 17635 4097 17644 4131
rect 17592 4088 17644 4097
rect 17868 4088 17920 4140
rect 18604 4224 18656 4276
rect 19248 4224 19300 4276
rect 19800 4224 19852 4276
rect 22284 4267 22336 4276
rect 22284 4233 22293 4267
rect 22293 4233 22327 4267
rect 22327 4233 22336 4267
rect 22284 4224 22336 4233
rect 23848 4224 23900 4276
rect 25320 4224 25372 4276
rect 23020 4199 23072 4208
rect 23020 4165 23029 4199
rect 23029 4165 23063 4199
rect 23063 4165 23072 4199
rect 23020 4156 23072 4165
rect 23296 4156 23348 4208
rect 23572 4156 23624 4208
rect 24308 4156 24360 4208
rect 25688 4156 25740 4208
rect 18144 4088 18196 4140
rect 19616 4088 19668 4140
rect 16120 4020 16172 4029
rect 17132 4020 17184 4072
rect 18972 4020 19024 4072
rect 19340 4063 19392 4072
rect 19340 4029 19349 4063
rect 19349 4029 19383 4063
rect 19383 4029 19392 4063
rect 19340 4020 19392 4029
rect 13820 3952 13872 4004
rect 14464 3952 14516 4004
rect 15292 3952 15344 4004
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16120 3884 16172 3936
rect 17224 3952 17276 4004
rect 18420 3952 18472 4004
rect 18604 3952 18656 4004
rect 19984 4088 20036 4140
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 17960 3884 18012 3936
rect 18512 3927 18564 3936
rect 18512 3893 18521 3927
rect 18521 3893 18555 3927
rect 18555 3893 18564 3927
rect 18512 3884 18564 3893
rect 18788 3927 18840 3936
rect 18788 3893 18797 3927
rect 18797 3893 18831 3927
rect 18831 3893 18840 3927
rect 18788 3884 18840 3893
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 20352 3884 20404 3936
rect 21824 3927 21876 3936
rect 21824 3893 21833 3927
rect 21833 3893 21867 3927
rect 21867 3893 21876 3927
rect 21824 3884 21876 3893
rect 22652 3927 22704 3936
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 23388 4131 23440 4140
rect 23388 4097 23397 4131
rect 23397 4097 23431 4131
rect 23431 4097 23440 4131
rect 23388 4088 23440 4097
rect 23664 4131 23716 4140
rect 23664 4097 23673 4131
rect 23673 4097 23707 4131
rect 23707 4097 23716 4131
rect 23664 4088 23716 4097
rect 23756 4131 23808 4140
rect 23756 4097 23765 4131
rect 23765 4097 23799 4131
rect 23799 4097 23808 4131
rect 23756 4088 23808 4097
rect 23020 4020 23072 4072
rect 23572 4020 23624 4072
rect 24032 4063 24084 4072
rect 24032 4029 24041 4063
rect 24041 4029 24075 4063
rect 24075 4029 24084 4063
rect 24032 4020 24084 4029
rect 25228 3884 25280 3936
rect 4124 3782 4176 3834
rect 4188 3782 4240 3834
rect 4252 3782 4304 3834
rect 4316 3782 4368 3834
rect 4380 3782 4432 3834
rect 10472 3782 10524 3834
rect 10536 3782 10588 3834
rect 10600 3782 10652 3834
rect 10664 3782 10716 3834
rect 10728 3782 10780 3834
rect 16820 3782 16872 3834
rect 16884 3782 16936 3834
rect 16948 3782 17000 3834
rect 17012 3782 17064 3834
rect 17076 3782 17128 3834
rect 23168 3782 23220 3834
rect 23232 3782 23284 3834
rect 23296 3782 23348 3834
rect 23360 3782 23412 3834
rect 23424 3782 23476 3834
rect 3332 3680 3384 3732
rect 3792 3680 3844 3732
rect 4804 3680 4856 3732
rect 4988 3723 5040 3732
rect 4988 3689 5018 3723
rect 5018 3689 5040 3723
rect 4988 3680 5040 3689
rect 5632 3680 5684 3732
rect 6368 3680 6420 3732
rect 6644 3680 6696 3732
rect 8852 3680 8904 3732
rect 14924 3680 14976 3732
rect 15936 3680 15988 3732
rect 16212 3680 16264 3732
rect 7012 3587 7064 3596
rect 1400 3476 1452 3528
rect 2872 3476 2924 3528
rect 4068 3476 4120 3528
rect 4528 3476 4580 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 10324 3544 10376 3596
rect 11520 3544 11572 3596
rect 14280 3612 14332 3664
rect 1768 3451 1820 3460
rect 1768 3417 1777 3451
rect 1777 3417 1811 3451
rect 1811 3417 1820 3451
rect 1768 3408 1820 3417
rect 2780 3340 2832 3392
rect 6920 3408 6972 3460
rect 4712 3340 4764 3392
rect 6276 3340 6328 3392
rect 8576 3408 8628 3460
rect 8208 3340 8260 3392
rect 9220 3408 9272 3460
rect 9496 3340 9548 3392
rect 9772 3383 9824 3392
rect 9772 3349 9781 3383
rect 9781 3349 9815 3383
rect 9815 3349 9824 3383
rect 9772 3340 9824 3349
rect 10232 3476 10284 3528
rect 13084 3476 13136 3528
rect 13268 3519 13320 3528
rect 13268 3485 13277 3519
rect 13277 3485 13311 3519
rect 13311 3485 13320 3519
rect 13268 3476 13320 3485
rect 13820 3544 13872 3596
rect 14832 3544 14884 3596
rect 17776 3680 17828 3732
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 18880 3544 18932 3596
rect 19984 3723 20036 3732
rect 19984 3689 19993 3723
rect 19993 3689 20027 3723
rect 20027 3689 20036 3723
rect 19984 3680 20036 3689
rect 20076 3680 20128 3732
rect 22744 3680 22796 3732
rect 23572 3680 23624 3732
rect 24032 3680 24084 3732
rect 24308 3680 24360 3732
rect 10968 3451 11020 3460
rect 10968 3417 10977 3451
rect 10977 3417 11011 3451
rect 11011 3417 11020 3451
rect 10968 3408 11020 3417
rect 11428 3408 11480 3460
rect 17132 3476 17184 3528
rect 18696 3476 18748 3528
rect 19156 3476 19208 3528
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 21272 3544 21324 3596
rect 21916 3544 21968 3596
rect 12808 3383 12860 3392
rect 12808 3349 12817 3383
rect 12817 3349 12851 3383
rect 12851 3349 12860 3383
rect 12808 3340 12860 3349
rect 14004 3408 14056 3460
rect 14096 3451 14148 3460
rect 14096 3417 14105 3451
rect 14105 3417 14139 3451
rect 14139 3417 14148 3451
rect 14096 3408 14148 3417
rect 14372 3408 14424 3460
rect 13452 3340 13504 3392
rect 14464 3383 14516 3392
rect 14464 3349 14473 3383
rect 14473 3349 14507 3383
rect 14507 3349 14516 3383
rect 14464 3340 14516 3349
rect 14832 3451 14884 3460
rect 14832 3417 14841 3451
rect 14841 3417 14875 3451
rect 14875 3417 14884 3451
rect 14832 3408 14884 3417
rect 14924 3408 14976 3460
rect 16304 3408 16356 3460
rect 17592 3451 17644 3460
rect 17592 3417 17601 3451
rect 17601 3417 17635 3451
rect 17635 3417 17644 3451
rect 17592 3408 17644 3417
rect 24584 3544 24636 3596
rect 25320 3680 25372 3732
rect 23020 3476 23072 3528
rect 23848 3519 23900 3528
rect 23848 3485 23857 3519
rect 23857 3485 23891 3519
rect 23891 3485 23900 3519
rect 23848 3476 23900 3485
rect 24860 3476 24912 3528
rect 25320 3519 25372 3528
rect 25320 3485 25329 3519
rect 25329 3485 25363 3519
rect 25363 3485 25372 3519
rect 25320 3476 25372 3485
rect 25412 3519 25464 3528
rect 25412 3485 25421 3519
rect 25421 3485 25455 3519
rect 25455 3485 25464 3519
rect 25412 3476 25464 3485
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 17408 3340 17460 3392
rect 19340 3340 19392 3392
rect 23756 3340 23808 3392
rect 7298 3238 7350 3290
rect 7362 3238 7414 3290
rect 7426 3238 7478 3290
rect 7490 3238 7542 3290
rect 7554 3238 7606 3290
rect 13646 3238 13698 3290
rect 13710 3238 13762 3290
rect 13774 3238 13826 3290
rect 13838 3238 13890 3290
rect 13902 3238 13954 3290
rect 19994 3238 20046 3290
rect 20058 3238 20110 3290
rect 20122 3238 20174 3290
rect 20186 3238 20238 3290
rect 20250 3238 20302 3290
rect 26342 3238 26394 3290
rect 26406 3238 26458 3290
rect 26470 3238 26522 3290
rect 26534 3238 26586 3290
rect 26598 3238 26650 3290
rect 1768 3136 1820 3188
rect 2688 3136 2740 3188
rect 3240 3136 3292 3188
rect 4528 3179 4580 3188
rect 4528 3145 4537 3179
rect 4537 3145 4571 3179
rect 4571 3145 4580 3179
rect 4528 3136 4580 3145
rect 4620 3136 4672 3188
rect 4712 3136 4764 3188
rect 5172 3136 5224 3188
rect 6092 3136 6144 3188
rect 7012 3136 7064 3188
rect 8116 3136 8168 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 8300 3136 8352 3188
rect 8392 3136 8444 3188
rect 9220 3136 9272 3188
rect 9772 3136 9824 3188
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 4068 3000 4120 3052
rect 6276 3068 6328 3120
rect 7932 3068 7984 3120
rect 9496 3068 9548 3120
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 10876 3136 10928 3188
rect 10968 3136 11020 3188
rect 11796 3136 11848 3188
rect 12808 3136 12860 3188
rect 13360 3068 13412 3120
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 12900 3000 12952 3052
rect 13820 3136 13872 3188
rect 14556 3068 14608 3120
rect 15016 3111 15068 3120
rect 15016 3077 15025 3111
rect 15025 3077 15059 3111
rect 15059 3077 15068 3111
rect 15016 3068 15068 3077
rect 15108 3111 15160 3120
rect 15108 3077 15143 3111
rect 15143 3077 15160 3111
rect 15108 3068 15160 3077
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 10232 2932 10284 2984
rect 14280 3000 14332 3052
rect 15660 3136 15712 3188
rect 16396 3136 16448 3188
rect 16672 3179 16724 3188
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 17592 3136 17644 3188
rect 18696 3068 18748 3120
rect 20352 3136 20404 3188
rect 20904 3136 20956 3188
rect 21824 3136 21876 3188
rect 14188 2932 14240 2984
rect 13268 2907 13320 2916
rect 13268 2873 13277 2907
rect 13277 2873 13311 2907
rect 13311 2873 13320 2907
rect 13268 2864 13320 2873
rect 14004 2864 14056 2916
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 16120 3000 16172 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 20628 3000 20680 3052
rect 22652 3136 22704 3188
rect 23756 3136 23808 3188
rect 25688 3136 25740 3188
rect 24308 3068 24360 3120
rect 17408 2932 17460 2984
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 14832 2864 14884 2916
rect 3240 2796 3292 2848
rect 6184 2796 6236 2848
rect 16028 2839 16080 2848
rect 16028 2805 16037 2839
rect 16037 2805 16071 2839
rect 16071 2805 16080 2839
rect 16028 2796 16080 2805
rect 17776 2864 17828 2916
rect 18512 2796 18564 2848
rect 4124 2694 4176 2746
rect 4188 2694 4240 2746
rect 4252 2694 4304 2746
rect 4316 2694 4368 2746
rect 4380 2694 4432 2746
rect 10472 2694 10524 2746
rect 10536 2694 10588 2746
rect 10600 2694 10652 2746
rect 10664 2694 10716 2746
rect 10728 2694 10780 2746
rect 16820 2694 16872 2746
rect 16884 2694 16936 2746
rect 16948 2694 17000 2746
rect 17012 2694 17064 2746
rect 17076 2694 17128 2746
rect 23168 2694 23220 2746
rect 23232 2694 23284 2746
rect 23296 2694 23348 2746
rect 23360 2694 23412 2746
rect 23424 2694 23476 2746
rect 9036 2592 9088 2644
rect 14740 2592 14792 2644
rect 18328 2592 18380 2644
rect 14096 2524 14148 2576
rect 10048 2456 10100 2508
rect 14924 2456 14976 2508
rect 16028 2456 16080 2508
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 18788 2456 18840 2508
rect 18052 2431 18104 2440
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 18052 2388 18104 2397
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 19156 2388 19208 2440
rect 25780 2431 25832 2440
rect 25780 2397 25789 2431
rect 25789 2397 25823 2431
rect 25823 2397 25832 2431
rect 25780 2388 25832 2397
rect 18512 2320 18564 2372
rect 26148 2363 26200 2372
rect 26148 2329 26157 2363
rect 26157 2329 26191 2363
rect 26191 2329 26200 2363
rect 26148 2320 26200 2329
rect 18052 2252 18104 2304
rect 7298 2150 7350 2202
rect 7362 2150 7414 2202
rect 7426 2150 7478 2202
rect 7490 2150 7542 2202
rect 7554 2150 7606 2202
rect 13646 2150 13698 2202
rect 13710 2150 13762 2202
rect 13774 2150 13826 2202
rect 13838 2150 13890 2202
rect 13902 2150 13954 2202
rect 19994 2150 20046 2202
rect 20058 2150 20110 2202
rect 20122 2150 20174 2202
rect 20186 2150 20238 2202
rect 20250 2150 20302 2202
rect 26342 2150 26394 2202
rect 26406 2150 26458 2202
rect 26470 2150 26522 2202
rect 26534 2150 26586 2202
rect 26598 2150 26650 2202
<< metal2 >>
rect 18 28985 74 29785
rect 3882 28985 3938 29785
rect 7746 28985 7802 29785
rect 10966 28985 11022 29785
rect 14830 28985 14886 29785
rect 18050 28985 18106 29785
rect 21914 28985 21970 29785
rect 25778 28985 25834 29785
rect 3896 26994 3924 28985
rect 10980 27554 11008 28985
rect 10980 27526 11100 27554
rect 7298 27228 7606 27237
rect 7298 27226 7304 27228
rect 7360 27226 7384 27228
rect 7440 27226 7464 27228
rect 7520 27226 7544 27228
rect 7600 27226 7606 27228
rect 7360 27174 7362 27226
rect 7542 27174 7544 27226
rect 7298 27172 7304 27174
rect 7360 27172 7384 27174
rect 7440 27172 7464 27174
rect 7520 27172 7544 27174
rect 7600 27172 7606 27174
rect 7298 27163 7606 27172
rect 11072 26994 11100 27526
rect 13646 27228 13954 27237
rect 13646 27226 13652 27228
rect 13708 27226 13732 27228
rect 13788 27226 13812 27228
rect 13868 27226 13892 27228
rect 13948 27226 13954 27228
rect 13708 27174 13710 27226
rect 13890 27174 13892 27226
rect 13646 27172 13652 27174
rect 13708 27172 13732 27174
rect 13788 27172 13812 27174
rect 13868 27172 13892 27174
rect 13948 27172 13954 27174
rect 13646 27163 13954 27172
rect 14844 26994 14872 28985
rect 19994 27228 20302 27237
rect 19994 27226 20000 27228
rect 20056 27226 20080 27228
rect 20136 27226 20160 27228
rect 20216 27226 20240 27228
rect 20296 27226 20302 27228
rect 20056 27174 20058 27226
rect 20238 27174 20240 27226
rect 19994 27172 20000 27174
rect 20056 27172 20080 27174
rect 20136 27172 20160 27174
rect 20216 27172 20240 27174
rect 20296 27172 20302 27174
rect 19994 27163 20302 27172
rect 26342 27228 26650 27237
rect 26342 27226 26348 27228
rect 26404 27226 26428 27228
rect 26484 27226 26508 27228
rect 26564 27226 26588 27228
rect 26644 27226 26650 27228
rect 26404 27174 26406 27226
rect 26586 27174 26588 27226
rect 26342 27172 26348 27174
rect 26404 27172 26428 27174
rect 26484 27172 26508 27174
rect 26564 27172 26588 27174
rect 26644 27172 26650 27174
rect 26342 27163 26650 27172
rect 21180 27124 21232 27130
rect 21180 27066 21232 27072
rect 17500 27056 17552 27062
rect 17500 26998 17552 27004
rect 3884 26988 3936 26994
rect 3884 26930 3936 26936
rect 11060 26988 11112 26994
rect 11060 26930 11112 26936
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 16580 26988 16632 26994
rect 16580 26930 16632 26936
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 940 26920 992 26926
rect 940 26862 992 26868
rect 952 26625 980 26862
rect 4124 26684 4432 26693
rect 4124 26682 4130 26684
rect 4186 26682 4210 26684
rect 4266 26682 4290 26684
rect 4346 26682 4370 26684
rect 4426 26682 4432 26684
rect 4186 26630 4188 26682
rect 4368 26630 4370 26682
rect 4124 26628 4130 26630
rect 4186 26628 4210 26630
rect 4266 26628 4290 26630
rect 4346 26628 4370 26630
rect 4426 26628 4432 26630
rect 938 26616 994 26625
rect 4124 26619 4432 26628
rect 10472 26684 10780 26693
rect 10472 26682 10478 26684
rect 10534 26682 10558 26684
rect 10614 26682 10638 26684
rect 10694 26682 10718 26684
rect 10774 26682 10780 26684
rect 10534 26630 10536 26682
rect 10716 26630 10718 26682
rect 10472 26628 10478 26630
rect 10534 26628 10558 26630
rect 10614 26628 10638 26630
rect 10694 26628 10718 26630
rect 10774 26628 10780 26630
rect 10472 26619 10780 26628
rect 16592 26586 16620 26930
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 938 26551 994 26560
rect 16580 26580 16632 26586
rect 16580 26522 16632 26528
rect 16212 26444 16264 26450
rect 16212 26386 16264 26392
rect 16580 26444 16632 26450
rect 16580 26386 16632 26392
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 11428 26376 11480 26382
rect 11428 26318 11480 26324
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 7298 26140 7606 26149
rect 7298 26138 7304 26140
rect 7360 26138 7384 26140
rect 7440 26138 7464 26140
rect 7520 26138 7544 26140
rect 7600 26138 7606 26140
rect 7360 26086 7362 26138
rect 7542 26086 7544 26138
rect 7298 26084 7304 26086
rect 7360 26084 7384 26086
rect 7440 26084 7464 26086
rect 7520 26084 7544 26086
rect 7600 26084 7606 26086
rect 7298 26075 7606 26084
rect 9324 25906 9352 26182
rect 8116 25900 8168 25906
rect 8116 25842 8168 25848
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 4124 25596 4432 25605
rect 4124 25594 4130 25596
rect 4186 25594 4210 25596
rect 4266 25594 4290 25596
rect 4346 25594 4370 25596
rect 4426 25594 4432 25596
rect 4186 25542 4188 25594
rect 4368 25542 4370 25594
rect 4124 25540 4130 25542
rect 4186 25540 4210 25542
rect 4266 25540 4290 25542
rect 4346 25540 4370 25542
rect 4426 25540 4432 25542
rect 4124 25531 4432 25540
rect 7298 25052 7606 25061
rect 7298 25050 7304 25052
rect 7360 25050 7384 25052
rect 7440 25050 7464 25052
rect 7520 25050 7544 25052
rect 7600 25050 7606 25052
rect 7360 24998 7362 25050
rect 7542 24998 7544 25050
rect 7298 24996 7304 24998
rect 7360 24996 7384 24998
rect 7440 24996 7464 24998
rect 7520 24996 7544 24998
rect 7600 24996 7606 24998
rect 7298 24987 7606 24996
rect 4124 24508 4432 24517
rect 4124 24506 4130 24508
rect 4186 24506 4210 24508
rect 4266 24506 4290 24508
rect 4346 24506 4370 24508
rect 4426 24506 4432 24508
rect 4186 24454 4188 24506
rect 4368 24454 4370 24506
rect 4124 24452 4130 24454
rect 4186 24452 4210 24454
rect 4266 24452 4290 24454
rect 4346 24452 4370 24454
rect 4426 24452 4432 24454
rect 4124 24443 4432 24452
rect 8128 24206 8156 25842
rect 9508 25498 9536 26318
rect 10324 26240 10376 26246
rect 10324 26182 10376 26188
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9140 24410 9168 24754
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 9600 24342 9628 24754
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9692 24410 9720 24686
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9784 24342 9812 25434
rect 9876 25226 9904 25638
rect 9968 25498 9996 25842
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 10232 25288 10284 25294
rect 10232 25230 10284 25236
rect 9864 25220 9916 25226
rect 9864 25162 9916 25168
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 9876 24886 9904 25162
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 10048 24676 10100 24682
rect 10048 24618 10100 24624
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9588 24336 9640 24342
rect 9588 24278 9640 24284
rect 9772 24336 9824 24342
rect 9772 24278 9824 24284
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 9404 24200 9456 24206
rect 9404 24142 9456 24148
rect 7748 24132 7800 24138
rect 7748 24074 7800 24080
rect 7298 23964 7606 23973
rect 7298 23962 7304 23964
rect 7360 23962 7384 23964
rect 7440 23962 7464 23964
rect 7520 23962 7544 23964
rect 7600 23962 7606 23964
rect 7360 23910 7362 23962
rect 7542 23910 7544 23962
rect 7298 23908 7304 23910
rect 7360 23908 7384 23910
rect 7440 23908 7464 23910
rect 7520 23908 7544 23910
rect 7600 23908 7606 23910
rect 7298 23899 7606 23908
rect 7760 23866 7788 24074
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 8128 23730 8156 24142
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 4124 23420 4432 23429
rect 4124 23418 4130 23420
rect 4186 23418 4210 23420
rect 4266 23418 4290 23420
rect 4346 23418 4370 23420
rect 4426 23418 4432 23420
rect 4186 23366 4188 23418
rect 4368 23366 4370 23418
rect 4124 23364 4130 23366
rect 4186 23364 4210 23366
rect 4266 23364 4290 23366
rect 4346 23364 4370 23366
rect 4426 23364 4432 23366
rect 4124 23355 4432 23364
rect 7298 22876 7606 22885
rect 7298 22874 7304 22876
rect 7360 22874 7384 22876
rect 7440 22874 7464 22876
rect 7520 22874 7544 22876
rect 7600 22874 7606 22876
rect 7360 22822 7362 22874
rect 7542 22822 7544 22874
rect 7298 22820 7304 22822
rect 7360 22820 7384 22822
rect 7440 22820 7464 22822
rect 7520 22820 7544 22822
rect 7600 22820 7606 22822
rect 7298 22811 7606 22820
rect 8128 22642 8156 23666
rect 9416 23526 9444 24142
rect 9404 23520 9456 23526
rect 9404 23462 9456 23468
rect 9416 23186 9444 23462
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9600 23118 9628 24278
rect 9784 23866 9812 24278
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9968 23594 9996 24550
rect 10060 23866 10088 24618
rect 10152 24614 10180 25162
rect 10244 24886 10272 25230
rect 10336 25226 10364 26182
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 10472 25596 10780 25605
rect 10472 25594 10478 25596
rect 10534 25594 10558 25596
rect 10614 25594 10638 25596
rect 10694 25594 10718 25596
rect 10774 25594 10780 25596
rect 10534 25542 10536 25594
rect 10716 25542 10718 25594
rect 10472 25540 10478 25542
rect 10534 25540 10558 25542
rect 10614 25540 10638 25542
rect 10694 25540 10718 25542
rect 10774 25540 10780 25542
rect 10472 25531 10780 25540
rect 10416 25288 10468 25294
rect 10416 25230 10468 25236
rect 10324 25220 10376 25226
rect 10324 25162 10376 25168
rect 10232 24880 10284 24886
rect 10232 24822 10284 24828
rect 10232 24744 10284 24750
rect 10428 24698 10456 25230
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10784 25152 10836 25158
rect 10836 25100 10916 25106
rect 10784 25094 10916 25100
rect 10612 24954 10640 25094
rect 10796 25078 10916 25094
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10888 24750 10916 25078
rect 10232 24686 10284 24692
rect 10140 24608 10192 24614
rect 10140 24550 10192 24556
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 10152 23594 10180 24346
rect 10244 24206 10272 24686
rect 10336 24670 10456 24698
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 10140 23588 10192 23594
rect 10140 23530 10192 23536
rect 10048 23248 10100 23254
rect 10244 23202 10272 24142
rect 10336 23730 10364 24670
rect 10472 24508 10780 24517
rect 10472 24506 10478 24508
rect 10534 24506 10558 24508
rect 10614 24506 10638 24508
rect 10694 24506 10718 24508
rect 10774 24506 10780 24508
rect 10534 24454 10536 24506
rect 10716 24454 10718 24506
rect 10472 24452 10478 24454
rect 10534 24452 10558 24454
rect 10614 24452 10638 24454
rect 10694 24452 10718 24454
rect 10774 24452 10780 24454
rect 10472 24443 10780 24452
rect 10888 24342 10916 24686
rect 10980 24614 11008 25842
rect 11244 25832 11296 25838
rect 11244 25774 11296 25780
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 11164 25226 11192 25638
rect 11256 25294 11284 25774
rect 11244 25288 11296 25294
rect 11244 25230 11296 25236
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 10980 24342 11008 24550
rect 10876 24336 10928 24342
rect 10876 24278 10928 24284
rect 10968 24336 11020 24342
rect 10968 24278 11020 24284
rect 11164 24206 11192 24550
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10472 23420 10780 23429
rect 10472 23418 10478 23420
rect 10534 23418 10558 23420
rect 10614 23418 10638 23420
rect 10694 23418 10718 23420
rect 10774 23418 10780 23420
rect 10534 23366 10536 23418
rect 10716 23366 10718 23418
rect 10472 23364 10478 23366
rect 10534 23364 10558 23366
rect 10614 23364 10638 23366
rect 10694 23364 10718 23366
rect 10774 23364 10780 23366
rect 10472 23355 10780 23364
rect 11164 23254 11192 24142
rect 10100 23196 10272 23202
rect 10048 23190 10272 23196
rect 11152 23248 11204 23254
rect 11152 23190 11204 23196
rect 10060 23186 10272 23190
rect 10060 23180 10284 23186
rect 10060 23174 10232 23180
rect 10232 23122 10284 23128
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 9680 22976 9732 22982
rect 9680 22918 9732 22924
rect 9692 22778 9720 22918
rect 9968 22778 9996 22986
rect 11164 22778 11192 23054
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 11256 22642 11284 25230
rect 11348 24954 11376 25842
rect 11440 25770 11468 26318
rect 12438 25936 12494 25945
rect 12360 25906 12438 25922
rect 12348 25900 12438 25906
rect 12400 25894 12438 25900
rect 12438 25871 12494 25880
rect 12348 25842 12400 25848
rect 12256 25832 12308 25838
rect 12254 25800 12256 25809
rect 12308 25800 12310 25809
rect 11428 25764 11480 25770
rect 12254 25735 12310 25744
rect 12440 25764 12492 25770
rect 11428 25706 11480 25712
rect 12440 25706 12492 25712
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11808 24274 11836 25638
rect 11992 24818 12020 25638
rect 12268 25158 12296 25638
rect 12452 25498 12480 25706
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 12256 25152 12308 25158
rect 12256 25094 12308 25100
rect 12268 24818 12296 25094
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12544 24750 12572 26318
rect 12624 26240 12676 26246
rect 12624 26182 12676 26188
rect 12636 25294 12664 26182
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12636 24750 12664 24890
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12532 24336 12584 24342
rect 12532 24278 12584 24284
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 11716 22642 11744 23054
rect 11808 22778 11836 23054
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 11992 22778 12020 22918
rect 12176 22778 12204 23054
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12544 22710 12572 24278
rect 12636 24206 12664 24686
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12728 24138 12756 24686
rect 12912 24410 12940 26318
rect 15660 26240 15712 26246
rect 15660 26182 15712 26188
rect 13646 26140 13954 26149
rect 13646 26138 13652 26140
rect 13708 26138 13732 26140
rect 13788 26138 13812 26140
rect 13868 26138 13892 26140
rect 13948 26138 13954 26140
rect 13708 26086 13710 26138
rect 13890 26086 13892 26138
rect 13646 26084 13652 26086
rect 13708 26084 13732 26086
rect 13788 26084 13812 26086
rect 13868 26084 13892 26086
rect 13948 26084 13954 26086
rect 13646 26075 13954 26084
rect 13544 25968 13596 25974
rect 14556 25968 14608 25974
rect 13544 25910 13596 25916
rect 13634 25936 13690 25945
rect 13360 25900 13412 25906
rect 13360 25842 13412 25848
rect 13372 24954 13400 25842
rect 13556 25770 13584 25910
rect 14556 25910 14608 25916
rect 13634 25871 13690 25880
rect 13544 25764 13596 25770
rect 13544 25706 13596 25712
rect 13452 25152 13504 25158
rect 13556 25140 13584 25706
rect 13648 25702 13676 25871
rect 14464 25832 14516 25838
rect 14462 25800 14464 25809
rect 14516 25800 14518 25809
rect 14462 25735 14518 25744
rect 13636 25696 13688 25702
rect 13636 25638 13688 25644
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 14292 25498 14320 25638
rect 14280 25492 14332 25498
rect 14280 25434 14332 25440
rect 14188 25356 14240 25362
rect 14188 25298 14240 25304
rect 13504 25112 13584 25140
rect 14004 25152 14056 25158
rect 13452 25094 13504 25100
rect 14004 25094 14056 25100
rect 13360 24948 13412 24954
rect 13360 24890 13412 24896
rect 13084 24880 13136 24886
rect 13084 24822 13136 24828
rect 13096 24410 13124 24822
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13372 24410 13400 24686
rect 13464 24682 13492 25094
rect 13646 25052 13954 25061
rect 13646 25050 13652 25052
rect 13708 25050 13732 25052
rect 13788 25050 13812 25052
rect 13868 25050 13892 25052
rect 13948 25050 13954 25052
rect 13708 24998 13710 25050
rect 13890 24998 13892 25050
rect 13646 24996 13652 24998
rect 13708 24996 13732 24998
rect 13788 24996 13812 24998
rect 13868 24996 13892 24998
rect 13948 24996 13954 24998
rect 13646 24987 13954 24996
rect 13452 24676 13504 24682
rect 13452 24618 13504 24624
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 13084 23248 13136 23254
rect 13084 23190 13136 23196
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 9312 22636 9364 22642
rect 9312 22578 9364 22584
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 4124 22332 4432 22341
rect 4124 22330 4130 22332
rect 4186 22330 4210 22332
rect 4266 22330 4290 22332
rect 4346 22330 4370 22332
rect 4426 22330 4432 22332
rect 4186 22278 4188 22330
rect 4368 22278 4370 22330
rect 4124 22276 4130 22278
rect 4186 22276 4210 22278
rect 4266 22276 4290 22278
rect 4346 22276 4370 22278
rect 4426 22276 4432 22278
rect 4124 22267 4432 22276
rect 7298 21788 7606 21797
rect 7298 21786 7304 21788
rect 7360 21786 7384 21788
rect 7440 21786 7464 21788
rect 7520 21786 7544 21788
rect 7600 21786 7606 21788
rect 7360 21734 7362 21786
rect 7542 21734 7544 21786
rect 7298 21732 7304 21734
rect 7360 21732 7384 21734
rect 7440 21732 7464 21734
rect 7520 21732 7544 21734
rect 7600 21732 7606 21734
rect 7298 21723 7606 21732
rect 8128 21690 8156 22578
rect 9324 22234 9352 22578
rect 9312 22228 9364 22234
rect 9312 22170 9364 22176
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 4124 21244 4432 21253
rect 4124 21242 4130 21244
rect 4186 21242 4210 21244
rect 4266 21242 4290 21244
rect 4346 21242 4370 21244
rect 4426 21242 4432 21244
rect 4186 21190 4188 21242
rect 4368 21190 4370 21242
rect 4124 21188 4130 21190
rect 4186 21188 4210 21190
rect 4266 21188 4290 21190
rect 4346 21188 4370 21190
rect 4426 21188 4432 21190
rect 4124 21179 4432 21188
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7298 20700 7606 20709
rect 7298 20698 7304 20700
rect 7360 20698 7384 20700
rect 7440 20698 7464 20700
rect 7520 20698 7544 20700
rect 7600 20698 7606 20700
rect 7360 20646 7362 20698
rect 7542 20646 7544 20698
rect 7298 20644 7304 20646
rect 7360 20644 7384 20646
rect 7440 20644 7464 20646
rect 7520 20644 7544 20646
rect 7600 20644 7606 20646
rect 7298 20635 7606 20644
rect 7852 20466 7880 20742
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 4124 20156 4432 20165
rect 4124 20154 4130 20156
rect 4186 20154 4210 20156
rect 4266 20154 4290 20156
rect 4346 20154 4370 20156
rect 4426 20154 4432 20156
rect 4186 20102 4188 20154
rect 4368 20102 4370 20154
rect 4124 20100 4130 20102
rect 4186 20100 4210 20102
rect 4266 20100 4290 20102
rect 4346 20100 4370 20102
rect 4426 20100 4432 20102
rect 4124 20091 4432 20100
rect 7576 20058 7604 20402
rect 7944 20058 7972 21422
rect 8024 20460 8076 20466
rect 8128 20448 8156 21626
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8076 20420 8156 20448
rect 8024 20402 8076 20408
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8312 19922 8340 20742
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8404 19854 8432 20810
rect 8588 20505 8616 20878
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8680 20602 8708 20742
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8574 20496 8630 20505
rect 8574 20431 8630 20440
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 940 19168 992 19174
rect 938 19136 940 19145
rect 992 19136 994 19145
rect 938 19071 994 19080
rect 1780 18426 1808 19314
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 4124 19068 4432 19077
rect 4124 19066 4130 19068
rect 4186 19066 4210 19068
rect 4266 19066 4290 19068
rect 4346 19066 4370 19068
rect 4426 19066 4432 19068
rect 4186 19014 4188 19066
rect 4368 19014 4370 19066
rect 4124 19012 4130 19014
rect 4186 19012 4210 19014
rect 4266 19012 4290 19014
rect 4346 19012 4370 19014
rect 4426 19012 4432 19014
rect 4124 19003 4432 19012
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 6380 18222 6408 18770
rect 6564 18358 6592 19110
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 4124 17980 4432 17989
rect 4124 17978 4130 17980
rect 4186 17978 4210 17980
rect 4266 17978 4290 17980
rect 4346 17978 4370 17980
rect 4426 17978 4432 17980
rect 4186 17926 4188 17978
rect 4368 17926 4370 17978
rect 4124 17924 4130 17926
rect 4186 17924 4210 17926
rect 4266 17924 4290 17926
rect 4346 17924 4370 17926
rect 4426 17924 4432 17926
rect 4124 17915 4432 17924
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 2424 16794 2452 17070
rect 3252 16794 3280 17070
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3988 16250 4016 17138
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4124 16892 4432 16901
rect 4124 16890 4130 16892
rect 4186 16890 4210 16892
rect 4266 16890 4290 16892
rect 4346 16890 4370 16892
rect 4426 16890 4432 16892
rect 4186 16838 4188 16890
rect 4368 16838 4370 16890
rect 4124 16836 4130 16838
rect 4186 16836 4210 16838
rect 4266 16836 4290 16838
rect 4346 16836 4370 16838
rect 4426 16836 4432 16838
rect 4124 16827 4432 16836
rect 4540 16590 4568 16934
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3148 16176 3200 16182
rect 3148 16118 3200 16124
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15201 1440 15438
rect 1398 15192 1454 15201
rect 1398 15127 1454 15136
rect 1688 14822 1716 15846
rect 1872 15706 1900 15982
rect 3160 15706 3188 16118
rect 4264 16046 4292 16458
rect 4448 16436 4476 16526
rect 4632 16436 4660 17478
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 4448 16408 4660 16436
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 13394 1716 14758
rect 2332 14618 2360 15438
rect 3160 15094 3188 15642
rect 3148 15088 3200 15094
rect 2976 15048 3148 15076
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1964 14074 1992 14282
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 14074 2268 14214
rect 2424 14074 2452 14894
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2700 13938 2728 14214
rect 2884 13938 2912 14214
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2700 13530 2728 13874
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1688 12986 1716 13194
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 2700 12850 2728 13466
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2792 12782 2820 13670
rect 2884 12918 2912 13874
rect 2976 13258 3004 15048
rect 3148 15030 3200 15036
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3252 14414 3280 14894
rect 3436 14414 3464 15982
rect 4124 15804 4432 15813
rect 4124 15802 4130 15804
rect 4186 15802 4210 15804
rect 4266 15802 4290 15804
rect 4346 15802 4370 15804
rect 4426 15802 4432 15804
rect 4186 15750 4188 15802
rect 4368 15750 4370 15802
rect 4124 15748 4130 15750
rect 4186 15748 4210 15750
rect 4266 15748 4290 15750
rect 4346 15748 4370 15750
rect 4426 15748 4432 15750
rect 4124 15739 4432 15748
rect 4908 15502 4936 17070
rect 5552 15910 5580 17070
rect 5828 16250 5856 17614
rect 6012 16454 6040 17682
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15570 5580 15846
rect 5736 15706 5764 16050
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4124 14716 4432 14725
rect 4124 14714 4130 14716
rect 4186 14714 4210 14716
rect 4266 14714 4290 14716
rect 4346 14714 4370 14716
rect 4426 14714 4432 14716
rect 4186 14662 4188 14714
rect 4368 14662 4370 14714
rect 4124 14660 4130 14662
rect 4186 14660 4210 14662
rect 4266 14660 4290 14662
rect 4346 14660 4370 14662
rect 4426 14660 4432 14662
rect 4124 14651 4432 14660
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2792 11812 2820 12718
rect 3068 12714 3096 14282
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3160 14074 3188 14214
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3252 13938 3280 14350
rect 3436 14074 3464 14350
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3252 13734 3280 13874
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12782 3188 13126
rect 3252 12782 3280 13670
rect 3436 13410 3464 14010
rect 3620 14006 3648 14214
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 4724 13870 4752 14418
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3344 13382 3464 13410
rect 3344 12782 3372 13382
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 3436 12102 3464 13262
rect 3528 13258 3556 13466
rect 3620 13462 3648 13806
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4124 13628 4432 13637
rect 4124 13626 4130 13628
rect 4186 13626 4210 13628
rect 4266 13626 4290 13628
rect 4346 13626 4370 13628
rect 4426 13626 4432 13628
rect 4186 13574 4188 13626
rect 4368 13574 4370 13626
rect 4124 13572 4130 13574
rect 4186 13572 4210 13574
rect 4266 13572 4290 13574
rect 4346 13572 4370 13574
rect 4426 13572 4432 13574
rect 4124 13563 4432 13572
rect 3608 13456 3660 13462
rect 3608 13398 3660 13404
rect 4436 13456 4488 13462
rect 4436 13398 4488 13404
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3516 12776 3568 12782
rect 3620 12764 3648 13398
rect 4448 13326 4476 13398
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 3568 12736 3648 12764
rect 3516 12718 3568 12724
rect 4448 12714 4476 13262
rect 4632 13190 4660 13670
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4436 12708 4488 12714
rect 4436 12650 4488 12656
rect 4124 12540 4432 12549
rect 4124 12538 4130 12540
rect 4186 12538 4210 12540
rect 4266 12538 4290 12540
rect 4346 12538 4370 12540
rect 4426 12538 4432 12540
rect 4186 12486 4188 12538
rect 4368 12486 4370 12538
rect 4124 12484 4130 12486
rect 4186 12484 4210 12486
rect 4266 12484 4290 12486
rect 4346 12484 4370 12486
rect 4426 12484 4432 12486
rect 4124 12475 4432 12484
rect 4632 12306 4660 12718
rect 4724 12434 4752 13194
rect 4816 12832 4844 14282
rect 4908 12986 4936 15302
rect 5460 14482 5488 15506
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 6012 14414 6040 16390
rect 6288 16182 6316 17138
rect 6380 16658 6408 18158
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 6380 15502 6408 16458
rect 6472 16250 6500 17070
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6472 15502 6500 15982
rect 6656 15502 6684 17478
rect 6932 16590 6960 18634
rect 7024 18630 7052 19654
rect 7298 19612 7606 19621
rect 7298 19610 7304 19612
rect 7360 19610 7384 19612
rect 7440 19610 7464 19612
rect 7520 19610 7544 19612
rect 7600 19610 7606 19612
rect 7360 19558 7362 19610
rect 7542 19558 7544 19610
rect 7298 19556 7304 19558
rect 7360 19556 7384 19558
rect 7440 19556 7464 19558
rect 7520 19556 7544 19558
rect 7600 19556 7606 19558
rect 7298 19547 7606 19556
rect 7668 19514 7696 19790
rect 8024 19780 8076 19786
rect 8076 19740 8340 19768
rect 8024 19722 8076 19728
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7944 19514 7972 19654
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7116 18970 7144 19314
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 8312 18834 8340 19740
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8588 19258 8616 20431
rect 8772 20058 8800 20878
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8772 19514 8800 19994
rect 8864 19854 8892 20742
rect 8956 20262 8984 20742
rect 9048 20534 9076 21490
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9600 20942 9628 21286
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9036 20528 9088 20534
rect 9036 20470 9088 20476
rect 9048 20398 9076 20470
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9416 20262 9444 20742
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 9232 19836 9260 19994
rect 9416 19854 9444 20198
rect 9312 19848 9364 19854
rect 9232 19808 9312 19836
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8404 18970 8432 19246
rect 8588 19230 8708 19258
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8300 18828 8352 18834
rect 8352 18788 8432 18816
rect 8300 18770 8352 18776
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 7298 18524 7606 18533
rect 7298 18522 7304 18524
rect 7360 18522 7384 18524
rect 7440 18522 7464 18524
rect 7520 18522 7544 18524
rect 7600 18522 7606 18524
rect 7360 18470 7362 18522
rect 7542 18470 7544 18522
rect 7298 18468 7304 18470
rect 7360 18468 7384 18470
rect 7440 18468 7464 18470
rect 7520 18468 7544 18470
rect 7600 18468 7606 18470
rect 7298 18459 7606 18468
rect 8128 18426 8156 18566
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6932 16182 6960 16526
rect 7024 16182 7052 16594
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 7116 15994 7144 18022
rect 7944 17542 7972 18226
rect 8220 17882 8248 18634
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18426 8340 18566
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8404 17882 8432 18788
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8496 17678 8524 19110
rect 8588 18358 8616 19110
rect 8680 18766 8708 19230
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8588 17882 8616 18294
rect 8864 18204 8892 19790
rect 8956 19514 8984 19790
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9048 19242 9076 19314
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 18358 9076 18566
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8944 18216 8996 18222
rect 8864 18176 8944 18204
rect 8944 18158 8996 18164
rect 9140 17882 9168 19450
rect 9232 18766 9260 19808
rect 9312 19790 9364 19796
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9416 19446 9444 19790
rect 9508 19514 9536 19790
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9508 18970 9536 19314
rect 9600 19174 9628 20878
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 19854 9720 20742
rect 9968 20482 9996 22578
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 10060 22030 10088 22374
rect 10472 22332 10780 22341
rect 10472 22330 10478 22332
rect 10534 22330 10558 22332
rect 10614 22330 10638 22332
rect 10694 22330 10718 22332
rect 10774 22330 10780 22332
rect 10534 22278 10536 22330
rect 10716 22278 10718 22330
rect 10472 22276 10478 22278
rect 10534 22276 10558 22278
rect 10614 22276 10638 22278
rect 10694 22276 10718 22278
rect 10774 22276 10780 22278
rect 10472 22267 10780 22276
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10472 21244 10780 21253
rect 10472 21242 10478 21244
rect 10534 21242 10558 21244
rect 10614 21242 10638 21244
rect 10694 21242 10718 21244
rect 10774 21242 10780 21244
rect 10534 21190 10536 21242
rect 10716 21190 10718 21242
rect 10472 21188 10478 21190
rect 10534 21188 10558 21190
rect 10614 21188 10638 21190
rect 10694 21188 10718 21190
rect 10774 21188 10780 21190
rect 10472 21179 10780 21188
rect 11256 20874 11284 22578
rect 11716 21894 11744 22578
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 12176 21554 12204 22578
rect 12544 22438 12572 22646
rect 13004 22574 13032 22986
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12360 21690 12388 21898
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 13096 21554 13124 23190
rect 13372 22778 13400 24346
rect 14016 24274 14044 25094
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 13646 23964 13954 23973
rect 13646 23962 13652 23964
rect 13708 23962 13732 23964
rect 13788 23962 13812 23964
rect 13868 23962 13892 23964
rect 13948 23962 13954 23964
rect 13708 23910 13710 23962
rect 13890 23910 13892 23962
rect 13646 23908 13652 23910
rect 13708 23908 13732 23910
rect 13788 23908 13812 23910
rect 13868 23908 13892 23910
rect 13948 23908 13954 23910
rect 13646 23899 13954 23908
rect 14200 23118 14228 25298
rect 14476 25294 14504 25735
rect 14568 25430 14596 25910
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14556 25424 14608 25430
rect 14556 25366 14608 25372
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14740 25288 14792 25294
rect 14740 25230 14792 25236
rect 14292 24818 14320 25230
rect 14476 24954 14504 25230
rect 14464 24948 14516 24954
rect 14464 24890 14516 24896
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14660 24410 14688 24754
rect 14752 24614 14780 25230
rect 14844 25226 14872 25638
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14936 24954 14964 25638
rect 15028 25498 15056 25842
rect 15016 25492 15068 25498
rect 15016 25434 15068 25440
rect 15672 25226 15700 26182
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 15752 25968 15804 25974
rect 15752 25910 15804 25916
rect 15660 25220 15712 25226
rect 15660 25162 15712 25168
rect 15764 24954 15792 25910
rect 15948 24954 15976 25978
rect 16040 25906 16068 26318
rect 16132 25974 16160 26318
rect 16120 25968 16172 25974
rect 16120 25910 16172 25916
rect 16224 25906 16252 26386
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16028 25900 16080 25906
rect 16028 25842 16080 25848
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16040 25430 16068 25842
rect 16028 25424 16080 25430
rect 16028 25366 16080 25372
rect 16040 24954 16068 25366
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 16132 24614 16160 25230
rect 16224 25158 16252 25842
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24954 16252 25094
rect 16212 24948 16264 24954
rect 16212 24890 16264 24896
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14280 23316 14332 23322
rect 14280 23258 14332 23264
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13452 22704 13504 22710
rect 13452 22646 13504 22652
rect 13464 22094 13492 22646
rect 13556 22234 13584 23054
rect 13646 22876 13954 22885
rect 13646 22874 13652 22876
rect 13708 22874 13732 22876
rect 13788 22874 13812 22876
rect 13868 22874 13892 22876
rect 13948 22874 13954 22876
rect 13708 22822 13710 22874
rect 13890 22822 13892 22874
rect 13646 22820 13652 22822
rect 13708 22820 13732 22822
rect 13788 22820 13812 22822
rect 13868 22820 13892 22822
rect 13948 22820 13954 22822
rect 13646 22811 13954 22820
rect 14004 22636 14056 22642
rect 14004 22578 14056 22584
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13740 22098 13768 22510
rect 14016 22234 14044 22578
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 13464 22066 13676 22094
rect 13648 22030 13676 22066
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 14292 22030 14320 23258
rect 14568 22030 14596 23598
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14660 21962 14688 23462
rect 14752 22098 14780 24550
rect 16132 24410 16160 24550
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 16224 24274 16252 24890
rect 16316 24342 16344 25230
rect 16408 24954 16436 25638
rect 16396 24948 16448 24954
rect 16396 24890 16448 24896
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 16500 24274 16528 26250
rect 16592 24818 16620 26386
rect 16684 25226 16712 26726
rect 16820 26684 17128 26693
rect 16820 26682 16826 26684
rect 16882 26682 16906 26684
rect 16962 26682 16986 26684
rect 17042 26682 17066 26684
rect 17122 26682 17128 26684
rect 16882 26630 16884 26682
rect 17064 26630 17066 26682
rect 16820 26628 16826 26630
rect 16882 26628 16906 26630
rect 16962 26628 16986 26630
rect 17042 26628 17066 26630
rect 17122 26628 17128 26630
rect 16820 26619 17128 26628
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16776 26042 16804 26318
rect 16764 26036 16816 26042
rect 16764 25978 16816 25984
rect 16820 25596 17128 25605
rect 16820 25594 16826 25596
rect 16882 25594 16906 25596
rect 16962 25594 16986 25596
rect 17042 25594 17066 25596
rect 17122 25594 17128 25596
rect 16882 25542 16884 25594
rect 17064 25542 17066 25594
rect 16820 25540 16826 25542
rect 16882 25540 16906 25542
rect 16962 25540 16986 25542
rect 17042 25540 17066 25542
rect 17122 25540 17128 25542
rect 16820 25531 17128 25540
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 17236 24886 17264 26930
rect 17512 26586 17540 26998
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 21008 26586 21036 26862
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 17316 25288 17368 25294
rect 17420 25242 17448 26522
rect 17512 26058 17540 26522
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 17512 26030 17632 26058
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17368 25236 17448 25242
rect 17316 25230 17448 25236
rect 17328 25214 17448 25230
rect 17224 24880 17276 24886
rect 17224 24822 17276 24828
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 17420 24682 17448 25214
rect 17512 24954 17540 25842
rect 17500 24948 17552 24954
rect 17500 24890 17552 24896
rect 17604 24818 17632 26030
rect 18064 25498 18092 26318
rect 19248 26240 19300 26246
rect 19248 26182 19300 26188
rect 19260 25974 19288 26182
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 19168 25294 19196 25842
rect 19156 25288 19208 25294
rect 19156 25230 19208 25236
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18064 24818 18092 25094
rect 18616 24886 18644 25094
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 19168 24818 19196 25230
rect 19352 24954 19380 25230
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 17592 24812 17644 24818
rect 17592 24754 17644 24760
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 18328 24744 18380 24750
rect 18328 24686 18380 24692
rect 17408 24676 17460 24682
rect 17408 24618 17460 24624
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 16820 24508 17128 24517
rect 16820 24506 16826 24508
rect 16882 24506 16906 24508
rect 16962 24506 16986 24508
rect 17042 24506 17066 24508
rect 17122 24506 17128 24508
rect 16882 24454 16884 24506
rect 17064 24454 17066 24506
rect 16820 24452 16826 24454
rect 16882 24452 16906 24454
rect 16962 24452 16986 24454
rect 17042 24452 17066 24454
rect 17122 24452 17128 24454
rect 16820 24443 17128 24452
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 16488 24268 16540 24274
rect 16488 24210 16540 24216
rect 16028 23724 16080 23730
rect 16080 23684 16160 23712
rect 16028 23666 16080 23672
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 15120 23322 15148 23462
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 14924 23112 14976 23118
rect 14924 23054 14976 23060
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 13646 21788 13954 21797
rect 13646 21786 13652 21788
rect 13708 21786 13732 21788
rect 13788 21786 13812 21788
rect 13868 21786 13892 21788
rect 13948 21786 13954 21788
rect 13708 21734 13710 21786
rect 13890 21734 13892 21786
rect 13646 21732 13652 21734
rect 13708 21732 13732 21734
rect 13788 21732 13812 21734
rect 13868 21732 13892 21734
rect 13948 21732 13954 21734
rect 13646 21723 13954 21732
rect 14752 21690 14780 22034
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 14752 21010 14780 21626
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 11256 20534 11284 20810
rect 11348 20602 11376 20946
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11244 20528 11296 20534
rect 9864 20460 9916 20466
rect 9968 20454 10180 20482
rect 11612 20528 11664 20534
rect 11244 20470 11296 20476
rect 11610 20496 11612 20505
rect 11664 20496 11666 20505
rect 9864 20402 9916 20408
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9416 18222 9444 18702
rect 9876 18698 9904 20402
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 10060 20058 10088 20334
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 7932 17536 7984 17542
rect 9140 17524 9168 17614
rect 9312 17536 9364 17542
rect 9140 17496 9312 17524
rect 7932 17478 7984 17484
rect 9312 17478 9364 17484
rect 7298 17436 7606 17445
rect 7298 17434 7304 17436
rect 7360 17434 7384 17436
rect 7440 17434 7464 17436
rect 7520 17434 7544 17436
rect 7600 17434 7606 17436
rect 7360 17382 7362 17434
rect 7542 17382 7544 17434
rect 7298 17380 7304 17382
rect 7360 17380 7384 17382
rect 7440 17380 7464 17382
rect 7520 17380 7544 17382
rect 7600 17380 7606 17382
rect 7298 17371 7606 17380
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 16794 7604 16934
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7298 16348 7606 16357
rect 7298 16346 7304 16348
rect 7360 16346 7384 16348
rect 7440 16346 7464 16348
rect 7520 16346 7544 16348
rect 7600 16346 7606 16348
rect 7360 16294 7362 16346
rect 7542 16294 7544 16346
rect 7298 16292 7304 16294
rect 7360 16292 7384 16294
rect 7440 16292 7464 16294
rect 7520 16292 7544 16294
rect 7600 16292 7606 16294
rect 7298 16283 7606 16292
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 6932 15966 7144 15994
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6472 15162 6500 15438
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6656 14618 6684 15438
rect 6748 15026 6776 15506
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5368 14074 5396 14214
rect 5552 14074 5580 14214
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5552 13938 5580 14010
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 5000 13394 5028 13670
rect 5184 13530 5212 13874
rect 5368 13734 5396 13874
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5092 13258 5120 13466
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 5000 12850 5028 13126
rect 4896 12844 4948 12850
rect 4816 12804 4896 12832
rect 4896 12786 4948 12792
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5000 12442 5028 12786
rect 4988 12436 5040 12442
rect 4724 12406 4844 12434
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 2872 11824 2924 11830
rect 2792 11784 2872 11812
rect 2872 11766 2924 11772
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 11354 2176 11494
rect 2884 11354 2912 11766
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10130 1440 11154
rect 3068 10742 3096 11562
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3160 11082 3188 11494
rect 3436 11286 3464 12038
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 3056 10736 3108 10742
rect 3056 10678 3108 10684
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 10266 2176 10406
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1872 9586 1900 10066
rect 3160 9994 3188 11018
rect 3528 10742 3556 11834
rect 3896 11762 3924 12174
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 3896 11354 3924 11698
rect 4448 11626 4476 11698
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4124 11452 4432 11461
rect 4124 11450 4130 11452
rect 4186 11450 4210 11452
rect 4266 11450 4290 11452
rect 4346 11450 4370 11452
rect 4426 11450 4432 11452
rect 4186 11398 4188 11450
rect 4368 11398 4370 11450
rect 4124 11396 4130 11398
rect 4186 11396 4210 11398
rect 4266 11396 4290 11398
rect 4346 11396 4370 11398
rect 4426 11396 4432 11398
rect 4124 11387 4432 11396
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3516 10736 3568 10742
rect 3516 10678 3568 10684
rect 3712 10674 3740 11018
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10810 3832 10950
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3896 10674 3924 11154
rect 4540 11082 4568 12174
rect 4816 11898 4844 12406
rect 5368 12434 5396 13670
rect 5552 13394 5580 13874
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5644 12918 5672 13670
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 4988 12378 5040 12384
rect 5276 12406 5396 12434
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10742 4384 10950
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4436 10692 4488 10698
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3884 10668 3936 10674
rect 4436 10634 4488 10640
rect 3884 10610 3936 10616
rect 4448 10554 4476 10634
rect 4540 10554 4568 11018
rect 4632 10826 4660 11290
rect 4724 11286 4752 11698
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4816 11218 4844 11834
rect 5276 11762 5304 12406
rect 5552 12238 5580 12650
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5644 12170 5672 12582
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5736 11762 5764 14350
rect 6656 13954 6684 14554
rect 6748 14074 6776 14962
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6656 13926 6776 13954
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5920 13190 5948 13806
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6012 12170 6040 12650
rect 6288 12442 6316 12854
rect 6380 12646 6408 13466
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6656 12442 6684 12786
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5000 11354 5028 11698
rect 5276 11558 5304 11698
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4632 10810 4752 10826
rect 4632 10804 4764 10810
rect 4632 10798 4712 10804
rect 4712 10746 4764 10752
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4448 10538 4568 10554
rect 4632 10538 4660 10678
rect 5092 10606 5120 11494
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5184 10742 5212 10950
rect 5276 10810 5304 11494
rect 6012 11354 6040 12106
rect 6564 11762 6592 12174
rect 6748 12102 6776 13926
rect 6840 13258 6868 14282
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12238 6868 12582
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 4436 10532 4568 10538
rect 4488 10526 4568 10532
rect 4620 10532 4672 10538
rect 4436 10474 4488 10480
rect 4620 10474 4672 10480
rect 3620 10266 3648 10474
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4124 10364 4432 10373
rect 4124 10362 4130 10364
rect 4186 10362 4210 10364
rect 4266 10362 4290 10364
rect 4346 10362 4370 10364
rect 4426 10362 4432 10364
rect 4186 10310 4188 10362
rect 4368 10310 4370 10362
rect 4124 10308 4130 10310
rect 4186 10308 4210 10310
rect 4266 10308 4290 10310
rect 4346 10308 4370 10310
rect 4426 10308 4432 10310
rect 4124 10299 4432 10308
rect 4540 10266 4568 10406
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 7546 1716 8366
rect 1872 8294 1900 9522
rect 3804 9330 3832 9930
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9518 3924 9862
rect 5184 9586 5212 10678
rect 5460 10538 5488 11086
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5552 10266 5580 11222
rect 6380 11150 6408 11630
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 5736 10810 5764 11086
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 6196 10606 6224 11018
rect 6840 10742 6868 11630
rect 6932 10810 6960 15966
rect 7484 15434 7512 16050
rect 7748 15700 7800 15706
rect 7944 15688 7972 17478
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 16250 8984 16390
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 9784 16130 9812 17614
rect 9876 17202 9904 18634
rect 9968 18290 9996 19450
rect 10060 18290 10088 19994
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9968 17746 9996 18226
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10060 17542 10088 18226
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 10152 16454 10180 20454
rect 11610 20431 11666 20440
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 10472 20156 10780 20165
rect 10472 20154 10478 20156
rect 10534 20154 10558 20156
rect 10614 20154 10638 20156
rect 10694 20154 10718 20156
rect 10774 20154 10780 20156
rect 10534 20102 10536 20154
rect 10716 20102 10718 20154
rect 10472 20100 10478 20102
rect 10534 20100 10558 20102
rect 10614 20100 10638 20102
rect 10694 20100 10718 20102
rect 10774 20100 10780 20102
rect 10472 20091 10780 20100
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 10520 19378 10548 19858
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10244 18884 10272 19178
rect 10336 18952 10364 19314
rect 10876 19304 10928 19310
rect 10414 19272 10470 19281
rect 10876 19246 10928 19252
rect 10414 19207 10416 19216
rect 10468 19207 10470 19216
rect 10416 19178 10468 19184
rect 10472 19068 10780 19077
rect 10472 19066 10478 19068
rect 10534 19066 10558 19068
rect 10614 19066 10638 19068
rect 10694 19066 10718 19068
rect 10774 19066 10780 19068
rect 10534 19014 10536 19066
rect 10716 19014 10718 19066
rect 10472 19012 10478 19014
rect 10534 19012 10558 19014
rect 10614 19012 10638 19014
rect 10694 19012 10718 19014
rect 10774 19012 10780 19014
rect 10472 19003 10780 19012
rect 10888 18952 10916 19246
rect 10336 18924 10456 18952
rect 10244 18856 10364 18884
rect 10336 18290 10364 18856
rect 10428 18766 10456 18924
rect 10704 18924 10916 18952
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10428 18154 10456 18702
rect 10704 18290 10732 18924
rect 11072 18290 11100 19314
rect 11164 18970 11192 19314
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10472 17980 10780 17989
rect 10472 17978 10478 17980
rect 10534 17978 10558 17980
rect 10614 17978 10638 17980
rect 10694 17978 10718 17980
rect 10774 17978 10780 17980
rect 10534 17926 10536 17978
rect 10716 17926 10718 17978
rect 10472 17924 10478 17926
rect 10534 17924 10558 17926
rect 10614 17924 10638 17926
rect 10694 17924 10718 17926
rect 10774 17924 10780 17926
rect 10472 17915 10780 17924
rect 10980 17134 11008 18158
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 17746 11100 18022
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11164 17610 11192 18702
rect 11256 18698 11284 19722
rect 11624 19446 11652 19722
rect 11900 19446 11928 20402
rect 11612 19440 11664 19446
rect 11888 19440 11940 19446
rect 11612 19382 11664 19388
rect 11716 19400 11888 19428
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11348 19242 11376 19314
rect 11336 19236 11388 19242
rect 11336 19178 11388 19184
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11256 18426 11284 18634
rect 11440 18426 11468 19314
rect 11716 18902 11744 19400
rect 11888 19382 11940 19388
rect 11992 19378 12020 20538
rect 12636 20058 12664 20810
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12820 20534 12848 20742
rect 13646 20700 13954 20709
rect 13646 20698 13652 20700
rect 13708 20698 13732 20700
rect 13788 20698 13812 20700
rect 13868 20698 13892 20700
rect 13948 20698 13954 20700
rect 13708 20646 13710 20698
rect 13890 20646 13892 20698
rect 13646 20644 13652 20646
rect 13708 20644 13732 20646
rect 13788 20644 13812 20646
rect 13868 20644 13892 20646
rect 13948 20644 13954 20646
rect 13646 20635 13954 20644
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12452 19378 12480 19926
rect 12636 19786 12664 19994
rect 12820 19854 12848 20334
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12624 19780 12676 19786
rect 12624 19722 12676 19728
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 11888 19304 11940 19310
rect 12268 19258 12296 19314
rect 11888 19246 11940 19252
rect 11900 18902 11928 19246
rect 11992 19230 12296 19258
rect 12360 19242 12388 19314
rect 12348 19236 12400 19242
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 16130 10180 16390
rect 10244 16250 10272 17070
rect 10472 16892 10780 16901
rect 10472 16890 10478 16892
rect 10534 16890 10558 16892
rect 10614 16890 10638 16892
rect 10694 16890 10718 16892
rect 10774 16890 10780 16892
rect 10534 16838 10536 16890
rect 10716 16838 10718 16890
rect 10472 16836 10478 16838
rect 10534 16836 10558 16838
rect 10614 16836 10638 16838
rect 10694 16836 10718 16838
rect 10774 16836 10780 16838
rect 10472 16827 10780 16836
rect 11256 16658 11284 18362
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11348 18154 11376 18226
rect 11336 18148 11388 18154
rect 11336 18090 11388 18096
rect 11348 17678 11376 18090
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11440 17542 11468 18362
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11532 17678 11560 18022
rect 11992 17882 12020 19230
rect 12348 19178 12400 19184
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12084 18290 12112 19110
rect 12176 18698 12204 19110
rect 12360 18850 12388 19178
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12268 18822 12388 18850
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12268 18290 12296 18822
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12084 18154 12296 18170
rect 12072 18148 12308 18154
rect 12124 18142 12256 18148
rect 12072 18090 12124 18096
rect 12256 18090 12308 18096
rect 12360 17882 12388 18702
rect 12452 18358 12480 18906
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12544 17814 12572 19450
rect 12636 19378 12664 19722
rect 12820 19718 12848 19790
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12820 19530 12848 19654
rect 12728 19502 12848 19530
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12622 19272 12678 19281
rect 12622 19207 12678 19216
rect 12636 18834 12664 19207
rect 12728 18902 12756 19502
rect 12912 19310 12940 19654
rect 13188 19514 13216 20402
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 13188 18766 13216 19450
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13372 18970 13400 19246
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 13096 18290 13124 18634
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13188 18086 13216 18702
rect 13464 18630 13492 20266
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 18970 13584 20198
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 13646 19612 13954 19621
rect 13646 19610 13652 19612
rect 13708 19610 13732 19612
rect 13788 19610 13812 19612
rect 13868 19610 13892 19612
rect 13948 19610 13954 19612
rect 13708 19558 13710 19610
rect 13890 19558 13892 19610
rect 13646 19556 13652 19558
rect 13708 19556 13732 19558
rect 13788 19556 13812 19558
rect 13868 19556 13892 19558
rect 13948 19556 13954 19558
rect 13646 19547 13954 19556
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13648 18850 13676 19110
rect 13556 18822 13676 18850
rect 13556 18766 13584 18822
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 18290 13492 18566
rect 13556 18290 13584 18702
rect 13646 18524 13954 18533
rect 13646 18522 13652 18524
rect 13708 18522 13732 18524
rect 13788 18522 13812 18524
rect 13868 18522 13892 18524
rect 13948 18522 13954 18524
rect 13708 18470 13710 18522
rect 13890 18470 13892 18522
rect 13646 18468 13652 18470
rect 13708 18468 13732 18470
rect 13788 18468 13812 18470
rect 13868 18468 13892 18470
rect 13948 18468 13954 18470
rect 13646 18459 13954 18468
rect 14016 18290 14044 19654
rect 14108 19174 14136 20402
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 14280 18896 14332 18902
rect 14280 18838 14332 18844
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18426 14136 18566
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11624 17338 11652 17546
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11440 16794 11468 16934
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 12084 16726 12112 17614
rect 12176 17066 12204 17614
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12268 17202 12296 17478
rect 12728 17338 12756 17546
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 9784 16102 9904 16130
rect 10060 16114 10180 16130
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 7800 15660 7972 15688
rect 7748 15642 7800 15648
rect 9692 15570 9720 15914
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7298 15260 7606 15269
rect 7298 15258 7304 15260
rect 7360 15258 7384 15260
rect 7440 15258 7464 15260
rect 7520 15258 7544 15260
rect 7600 15258 7606 15260
rect 7360 15206 7362 15258
rect 7542 15206 7544 15258
rect 7298 15204 7304 15206
rect 7360 15204 7384 15206
rect 7440 15204 7464 15206
rect 7520 15204 7544 15206
rect 7600 15204 7606 15206
rect 7298 15195 7606 15204
rect 9692 15162 9720 15506
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 7668 14618 7696 14894
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7380 14272 7432 14278
rect 7208 14232 7380 14260
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7024 13394 7052 13670
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7024 12986 7052 13330
rect 7116 12986 7144 13942
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7208 12434 7236 14232
rect 7380 14214 7432 14220
rect 7298 14172 7606 14181
rect 7298 14170 7304 14172
rect 7360 14170 7384 14172
rect 7440 14170 7464 14172
rect 7520 14170 7544 14172
rect 7600 14170 7606 14172
rect 7360 14118 7362 14170
rect 7542 14118 7544 14170
rect 7298 14116 7304 14118
rect 7360 14116 7384 14118
rect 7440 14116 7464 14118
rect 7520 14116 7544 14118
rect 7600 14116 7606 14118
rect 7298 14107 7606 14116
rect 8208 13524 8260 13530
rect 8312 13512 8340 14350
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8484 14272 8536 14278
rect 8680 14260 8708 14758
rect 8772 14482 8800 14826
rect 9600 14618 9628 14894
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8772 14362 8800 14418
rect 9692 14414 9720 15098
rect 9784 14550 9812 15982
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9680 14408 9732 14414
rect 8772 14334 8892 14362
rect 9680 14350 9732 14356
rect 9876 14346 9904 16102
rect 10048 16108 10180 16114
rect 10100 16102 10180 16108
rect 10048 16050 10100 16056
rect 10152 15706 10180 16102
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10152 15450 10180 15642
rect 10336 15586 10364 16594
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10796 15994 10824 16458
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10796 15966 10916 15994
rect 10472 15804 10780 15813
rect 10472 15802 10478 15804
rect 10534 15802 10558 15804
rect 10614 15802 10638 15804
rect 10694 15802 10718 15804
rect 10774 15802 10780 15804
rect 10534 15750 10536 15802
rect 10716 15750 10718 15802
rect 10472 15748 10478 15750
rect 10534 15748 10558 15750
rect 10614 15748 10638 15750
rect 10694 15748 10718 15750
rect 10774 15748 10780 15750
rect 10472 15739 10780 15748
rect 10336 15558 10456 15586
rect 10060 15422 10180 15450
rect 10060 15026 10088 15422
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10152 15026 10180 15302
rect 10336 15162 10364 15302
rect 10428 15162 10456 15558
rect 10888 15162 10916 15966
rect 10980 15434 11008 16390
rect 11256 16250 11284 16594
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11256 15570 11284 16186
rect 12084 16114 12112 16662
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 8536 14232 8708 14260
rect 8760 14272 8812 14278
rect 8484 14214 8536 14220
rect 8760 14214 8812 14220
rect 8404 13530 8432 14214
rect 8260 13484 8340 13512
rect 8392 13524 8444 13530
rect 8208 13466 8260 13472
rect 8392 13466 8444 13472
rect 8496 13410 8524 14214
rect 8772 14006 8800 14214
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8404 13394 8524 13410
rect 8392 13388 8524 13394
rect 8444 13382 8524 13388
rect 8392 13330 8444 13336
rect 7298 13084 7606 13093
rect 7298 13082 7304 13084
rect 7360 13082 7384 13084
rect 7440 13082 7464 13084
rect 7520 13082 7544 13084
rect 7600 13082 7606 13084
rect 7360 13030 7362 13082
rect 7542 13030 7544 13082
rect 7298 13028 7304 13030
rect 7360 13028 7384 13030
rect 7440 13028 7464 13030
rect 7520 13028 7544 13030
rect 7600 13028 7606 13030
rect 7298 13019 7606 13028
rect 8864 12850 8892 14334
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8956 12850 8984 13262
rect 9140 12986 9168 13670
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 12986 9812 13330
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 7116 12406 7236 12434
rect 7116 12238 7144 12406
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11762 7052 12038
rect 7298 11996 7606 12005
rect 7298 11994 7304 11996
rect 7360 11994 7384 11996
rect 7440 11994 7464 11996
rect 7520 11994 7544 11996
rect 7600 11994 7606 11996
rect 7360 11942 7362 11994
rect 7542 11942 7544 11994
rect 7298 11940 7304 11942
rect 7360 11940 7384 11942
rect 7440 11940 7464 11942
rect 7520 11940 7544 11942
rect 7600 11940 7606 11942
rect 7298 11931 7606 11940
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7116 11642 7144 11834
rect 7024 11614 7144 11642
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6656 10266 6684 10542
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6840 10130 6868 10678
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 5552 9722 5580 10066
rect 7024 9994 7052 11614
rect 7298 10908 7606 10917
rect 7298 10906 7304 10908
rect 7360 10906 7384 10908
rect 7440 10906 7464 10908
rect 7520 10906 7544 10908
rect 7600 10906 7606 10908
rect 7360 10854 7362 10906
rect 7542 10854 7544 10906
rect 7298 10852 7304 10854
rect 7360 10852 7384 10854
rect 7440 10852 7464 10854
rect 7520 10852 7544 10854
rect 7600 10852 7606 10854
rect 7298 10843 7606 10852
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7208 10062 7236 10610
rect 7760 10062 7788 12310
rect 8128 12238 8156 12718
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8128 11694 8156 12174
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8128 11354 8156 11630
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8496 11150 8524 11698
rect 8588 11218 8616 12038
rect 8772 11642 8800 12038
rect 8864 11830 8892 12786
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8956 11762 8984 12582
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8772 11614 8892 11642
rect 9232 11626 9260 12854
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9692 12434 9720 12786
rect 9324 12406 9720 12434
rect 9324 12170 9352 12406
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9324 11898 9352 12106
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 8864 11558 8892 11614
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8864 11150 8892 11494
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 9232 11082 9260 11562
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8312 10742 8340 10950
rect 8956 10810 8984 10950
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 9324 10674 9352 11834
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 8116 10464 8168 10470
rect 8168 10412 8248 10418
rect 8116 10406 8248 10412
rect 8128 10390 8248 10406
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3884 9376 3936 9382
rect 3804 9324 3884 9330
rect 3804 9318 3936 9324
rect 3804 9302 3924 9318
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 7886 1900 8230
rect 2884 7954 2912 8774
rect 3528 8498 3556 8910
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 2792 7206 2820 7754
rect 3344 7342 3372 8230
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6322 2820 7142
rect 3436 6866 3464 8434
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3528 6866 3556 7346
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 6458 3188 6734
rect 3528 6458 3556 6802
rect 3620 6730 3648 8434
rect 3712 8362 3740 8774
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5234 1440 6190
rect 2792 5522 2820 6258
rect 3160 5914 3188 6394
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3620 5914 3648 6258
rect 3712 6186 3740 8298
rect 3804 7546 3832 8774
rect 3896 8634 3924 9302
rect 4124 9276 4432 9285
rect 4124 9274 4130 9276
rect 4186 9274 4210 9276
rect 4266 9274 4290 9276
rect 4346 9274 4370 9276
rect 4426 9274 4432 9276
rect 4186 9222 4188 9274
rect 4368 9222 4370 9274
rect 4124 9220 4130 9222
rect 4186 9220 4210 9222
rect 4266 9220 4290 9222
rect 4346 9220 4370 9222
rect 4426 9220 4432 9222
rect 4124 9211 4432 9220
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3896 7478 3924 8570
rect 4080 8566 4108 8910
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4172 8276 4200 8978
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4540 8634 4568 8910
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4528 8628 4580 8634
rect 4580 8588 4660 8616
rect 4528 8570 4580 8576
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 3988 8248 4200 8276
rect 3988 8090 4016 8248
rect 4124 8188 4432 8197
rect 4124 8186 4130 8188
rect 4186 8186 4210 8188
rect 4266 8186 4290 8188
rect 4346 8186 4370 8188
rect 4426 8186 4432 8188
rect 4186 8134 4188 8186
rect 4368 8134 4370 8186
rect 4124 8132 4130 8134
rect 4186 8132 4210 8134
rect 4266 8132 4290 8134
rect 4346 8132 4370 8134
rect 4426 8132 4432 8134
rect 4124 8123 4432 8132
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3804 6458 3832 6870
rect 3988 6730 4016 7822
rect 4080 7585 4108 8026
rect 4540 8022 4568 8366
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4528 7880 4580 7886
rect 4632 7834 4660 8588
rect 4580 7828 4660 7834
rect 4528 7822 4660 7828
rect 4540 7806 4660 7822
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 4124 7100 4432 7109
rect 4124 7098 4130 7100
rect 4186 7098 4210 7100
rect 4266 7098 4290 7100
rect 4346 7098 4370 7100
rect 4426 7098 4432 7100
rect 4186 7046 4188 7098
rect 4368 7046 4370 7098
rect 4124 7044 4130 7046
rect 4186 7044 4210 7046
rect 4266 7044 4290 7046
rect 4346 7044 4370 7046
rect 4426 7044 4432 7046
rect 4124 7035 4432 7044
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3896 6458 3924 6666
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3988 6390 4016 6666
rect 4356 6662 4384 6938
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3712 5794 3740 6122
rect 4080 6100 4108 6598
rect 4632 6390 4660 7686
rect 4724 7478 4752 8774
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4528 6248 4580 6254
rect 4724 6236 4752 6734
rect 4816 6458 4844 8910
rect 5552 8566 5580 9658
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 4988 8424 5040 8430
rect 5552 8378 5580 8502
rect 5920 8498 5948 9114
rect 6932 8974 6960 9862
rect 7024 9722 7052 9930
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7024 9042 7052 9522
rect 7208 9518 7236 9998
rect 7298 9820 7606 9829
rect 7298 9818 7304 9820
rect 7360 9818 7384 9820
rect 7440 9818 7464 9820
rect 7520 9818 7544 9820
rect 7600 9818 7606 9820
rect 7360 9766 7362 9818
rect 7542 9766 7544 9818
rect 7298 9764 7304 9766
rect 7360 9764 7384 9766
rect 7440 9764 7464 9766
rect 7520 9764 7544 9766
rect 7600 9764 7606 9766
rect 7298 9755 7606 9764
rect 7668 9722 7696 9998
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7576 9602 7604 9658
rect 7576 9574 7696 9602
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 4988 8366 5040 8372
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4908 6390 4936 7278
rect 5000 7206 5028 8366
rect 5460 8350 5580 8378
rect 5460 7954 5488 8350
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5184 7342 5212 7822
rect 5920 7410 5948 8434
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6390 5028 7142
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 4580 6208 4752 6236
rect 4528 6190 4580 6196
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 3620 5766 3740 5794
rect 3988 6072 4108 6100
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 2792 5494 2912 5522
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 3534 1440 5170
rect 2884 5166 2912 5494
rect 3252 5302 3280 5578
rect 3620 5574 3648 5766
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1780 3194 1808 3402
rect 2700 3194 2728 3878
rect 2884 3534 2912 5102
rect 3252 4758 3280 5238
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 3068 4282 3096 4626
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3528 4146 3556 5306
rect 3712 5234 3740 5510
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3620 4826 3648 5170
rect 3712 4826 3740 5170
rect 3896 5030 3924 5646
rect 3988 5166 4016 6072
rect 4124 6012 4432 6021
rect 4124 6010 4130 6012
rect 4186 6010 4210 6012
rect 4266 6010 4290 6012
rect 4346 6010 4370 6012
rect 4426 6010 4432 6012
rect 4186 5958 4188 6010
rect 4368 5958 4370 6010
rect 4124 5956 4130 5958
rect 4186 5956 4210 5958
rect 4266 5956 4290 5958
rect 4346 5956 4370 5958
rect 4426 5956 4432 5958
rect 4124 5947 4432 5956
rect 4816 5914 4844 6122
rect 4908 5914 4936 6326
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5302 4108 5510
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3804 4298 3832 4626
rect 3896 4554 3924 4966
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 3804 4270 3924 4298
rect 3896 4146 3924 4270
rect 3988 4214 4016 5102
rect 4448 5012 4476 5850
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4448 4984 4568 5012
rect 4124 4924 4432 4933
rect 4124 4922 4130 4924
rect 4186 4922 4210 4924
rect 4266 4922 4290 4924
rect 4346 4922 4370 4924
rect 4426 4922 4432 4924
rect 4186 4870 4188 4922
rect 4368 4870 4370 4922
rect 4124 4868 4130 4870
rect 4186 4868 4210 4870
rect 4266 4868 4290 4870
rect 4346 4868 4370 4870
rect 4426 4868 4432 4870
rect 4124 4859 4432 4868
rect 4540 4622 4568 4984
rect 4724 4758 4752 5034
rect 4816 5030 4844 5646
rect 4908 5370 4936 5850
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 5092 4826 5120 5646
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 3058 2820 3334
rect 3252 3194 3280 3878
rect 3344 3738 3372 3946
rect 3804 3738 3832 4082
rect 4448 3942 4476 4422
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4124 3836 4432 3845
rect 4124 3834 4130 3836
rect 4186 3834 4210 3836
rect 4266 3834 4290 3836
rect 4346 3834 4370 3836
rect 4426 3834 4432 3836
rect 4186 3782 4188 3834
rect 4368 3782 4370 3834
rect 4124 3780 4130 3782
rect 4186 3780 4210 3782
rect 4266 3780 4290 3782
rect 4346 3780 4370 3782
rect 4426 3780 4432 3782
rect 4124 3771 4432 3780
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 4632 3618 4660 3878
rect 4540 3590 4660 3618
rect 4540 3534 4568 3590
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 4080 3058 4108 3470
rect 4540 3194 4568 3470
rect 4632 3194 4660 3470
rect 4724 3398 4752 4490
rect 4816 3738 4844 4762
rect 5184 4554 5212 5102
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5184 4298 5212 4490
rect 5092 4270 5212 4298
rect 5092 4078 5120 4270
rect 5368 4146 5396 6122
rect 5552 5914 5580 6190
rect 5644 5914 5672 6258
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5736 5370 5764 6258
rect 5920 6118 5948 7346
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 6012 6458 6040 6666
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4622 5580 4966
rect 5828 4826 5856 6054
rect 5920 5166 5948 6054
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4282 5580 4422
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5460 4146 5488 4218
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5000 3738 5028 3878
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3194 4752 3334
rect 5184 3194 5212 4082
rect 5644 3738 5672 4490
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5736 4078 5764 4422
rect 5828 4214 5856 4762
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5920 4146 5948 4966
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 4282 6040 4558
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 6104 3194 6132 3946
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 6196 2854 6224 8842
rect 6564 8514 6592 8910
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6472 8486 6592 8514
rect 6840 8498 6868 8774
rect 6828 8492 6880 8498
rect 6472 5642 6500 8486
rect 6828 8434 6880 8440
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6564 7954 6592 8366
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7478 6960 7754
rect 7116 7546 7144 7890
rect 7208 7750 7236 9454
rect 7298 8732 7606 8741
rect 7298 8730 7304 8732
rect 7360 8730 7384 8732
rect 7440 8730 7464 8732
rect 7520 8730 7544 8732
rect 7600 8730 7606 8732
rect 7360 8678 7362 8730
rect 7542 8678 7544 8730
rect 7298 8676 7304 8678
rect 7360 8676 7384 8678
rect 7440 8676 7464 8678
rect 7520 8676 7544 8678
rect 7600 8676 7606 8678
rect 7298 8667 7606 8676
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 7818 7328 8230
rect 7668 7818 7696 9574
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 8498 7788 9318
rect 7852 8974 7880 9658
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7944 8498 7972 9862
rect 8128 9722 8156 9998
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8220 9518 8248 10390
rect 9324 9908 9352 10610
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9416 10266 9444 10474
rect 9508 10266 9536 12242
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9600 11898 9628 12174
rect 9876 12050 9904 13398
rect 9968 13326 9996 14758
rect 10472 14716 10780 14725
rect 10472 14714 10478 14716
rect 10534 14714 10558 14716
rect 10614 14714 10638 14716
rect 10694 14714 10718 14716
rect 10774 14714 10780 14716
rect 10534 14662 10536 14714
rect 10716 14662 10718 14714
rect 10472 14660 10478 14662
rect 10534 14660 10558 14662
rect 10614 14660 10638 14662
rect 10694 14660 10718 14662
rect 10774 14660 10780 14662
rect 10472 14651 10780 14660
rect 11256 14482 11284 15506
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 13870 10088 14214
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9692 12022 9904 12050
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9692 11830 9720 12022
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 11354 9812 11698
rect 10060 11694 10088 12718
rect 10152 12646 10180 14282
rect 10336 13394 10364 14350
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10472 13628 10780 13637
rect 10472 13626 10478 13628
rect 10534 13626 10558 13628
rect 10614 13626 10638 13628
rect 10694 13626 10718 13628
rect 10774 13626 10780 13628
rect 10534 13574 10536 13626
rect 10716 13574 10718 13626
rect 10472 13572 10478 13574
rect 10534 13572 10558 13574
rect 10614 13572 10638 13574
rect 10694 13572 10718 13574
rect 10774 13572 10780 13574
rect 10472 13563 10780 13572
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10888 13326 10916 13738
rect 11256 13394 11284 14418
rect 11532 13938 11560 14894
rect 11992 14006 12020 15846
rect 12084 14958 12112 16050
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 15162 12296 15302
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12544 15026 12572 16526
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12636 16153 12664 16390
rect 12728 16182 12756 16390
rect 12912 16250 12940 17138
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 12716 16176 12768 16182
rect 12622 16144 12678 16153
rect 12716 16118 12768 16124
rect 12622 16079 12678 16088
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12912 15706 12940 15982
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12360 14618 12388 14758
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12636 14346 12664 15438
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9692 10810 9720 11290
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9324 9880 9444 9908
rect 9416 9722 9444 9880
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8036 8634 8064 8910
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7298 7644 7606 7653
rect 7298 7642 7304 7644
rect 7360 7642 7384 7644
rect 7440 7642 7464 7644
rect 7520 7642 7544 7644
rect 7600 7642 7606 7644
rect 7360 7590 7362 7642
rect 7542 7590 7544 7642
rect 7298 7588 7304 7590
rect 7360 7588 7384 7590
rect 7440 7588 7464 7590
rect 7520 7588 7544 7590
rect 7600 7588 7606 7590
rect 7298 7579 7606 7588
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6564 5914 6592 6054
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6932 5778 6960 7414
rect 7116 6254 7144 7482
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7944 6866 7972 7142
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7298 6556 7606 6565
rect 7298 6554 7304 6556
rect 7360 6554 7384 6556
rect 7440 6554 7464 6556
rect 7520 6554 7544 6556
rect 7600 6554 7606 6556
rect 7360 6502 7362 6554
rect 7542 6502 7544 6554
rect 7298 6500 7304 6502
rect 7360 6500 7384 6502
rect 7440 6500 7464 6502
rect 7520 6500 7544 6502
rect 7600 6500 7606 6502
rect 7298 6491 7606 6500
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 8036 6202 8064 8570
rect 8128 8566 8156 9318
rect 8220 9178 8248 9454
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8220 9042 8248 9114
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8312 8906 8340 9318
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8772 8294 8800 9454
rect 9416 8566 9444 9658
rect 9508 8634 9536 10202
rect 10152 9994 10180 12582
rect 10472 12540 10780 12549
rect 10472 12538 10478 12540
rect 10534 12538 10558 12540
rect 10614 12538 10638 12540
rect 10694 12538 10718 12540
rect 10774 12538 10780 12540
rect 10534 12486 10536 12538
rect 10716 12486 10718 12538
rect 10472 12484 10478 12486
rect 10534 12484 10558 12486
rect 10614 12484 10638 12486
rect 10694 12484 10718 12486
rect 10774 12484 10780 12486
rect 10472 12475 10780 12484
rect 11072 12306 11100 12718
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11898 10548 12038
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10472 11452 10780 11461
rect 10472 11450 10478 11452
rect 10534 11450 10558 11452
rect 10614 11450 10638 11452
rect 10694 11450 10718 11452
rect 10774 11450 10780 11452
rect 10534 11398 10536 11450
rect 10716 11398 10718 11450
rect 10472 11396 10478 11398
rect 10534 11396 10558 11398
rect 10614 11396 10638 11398
rect 10694 11396 10718 11398
rect 10774 11396 10780 11398
rect 10472 11387 10780 11396
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10472 10364 10780 10373
rect 10472 10362 10478 10364
rect 10534 10362 10558 10364
rect 10614 10362 10638 10364
rect 10694 10362 10718 10364
rect 10774 10362 10780 10364
rect 10534 10310 10536 10362
rect 10716 10310 10718 10362
rect 10472 10308 10478 10310
rect 10534 10308 10558 10310
rect 10614 10308 10638 10310
rect 10694 10308 10718 10310
rect 10774 10308 10780 10310
rect 10472 10299 10780 10308
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 9178 9720 9454
rect 10472 9276 10780 9285
rect 10472 9274 10478 9276
rect 10534 9274 10558 9276
rect 10614 9274 10638 9276
rect 10694 9274 10718 9276
rect 10774 9274 10780 9276
rect 10534 9222 10536 9274
rect 10716 9222 10718 9274
rect 10472 9220 10478 9222
rect 10534 9220 10558 9222
rect 10614 9220 10638 9222
rect 10694 9220 10718 9222
rect 10774 9220 10780 9222
rect 10472 9211 10780 9220
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9404 8560 9456 8566
rect 9456 8508 9812 8514
rect 9404 8502 9812 8508
rect 9416 8486 9812 8502
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8772 7954 8800 8230
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6458 8248 6734
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8128 6338 8156 6394
rect 8312 6338 8340 7890
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 6866 9536 7142
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9692 6662 9720 7482
rect 9784 7478 9812 8486
rect 10060 8022 10088 8842
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8634 10272 8774
rect 10888 8634 10916 10610
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10266 11008 10406
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11072 10130 11100 12242
rect 11164 11762 11192 13126
rect 11532 12374 11560 13874
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13394 11652 13670
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 12452 12918 12480 14214
rect 12636 13870 12664 14282
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12636 13258 12664 13806
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 13394 12940 13670
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11900 12442 11928 12718
rect 13004 12646 13032 17138
rect 13556 16538 13584 18022
rect 13646 17436 13954 17445
rect 13646 17434 13652 17436
rect 13708 17434 13732 17436
rect 13788 17434 13812 17436
rect 13868 17434 13892 17436
rect 13948 17434 13954 17436
rect 13708 17382 13710 17434
rect 13890 17382 13892 17434
rect 13646 17380 13652 17382
rect 13708 17380 13732 17382
rect 13788 17380 13812 17382
rect 13868 17380 13892 17382
rect 13948 17380 13954 17382
rect 13646 17371 13954 17380
rect 13372 16510 13584 16538
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 15706 13308 16390
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 13004 12238 13032 12582
rect 13188 12238 13216 13126
rect 13372 12238 13400 16510
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13464 15502 13492 16186
rect 13556 16046 13584 16390
rect 13646 16348 13954 16357
rect 13646 16346 13652 16348
rect 13708 16346 13732 16348
rect 13788 16346 13812 16348
rect 13868 16346 13892 16348
rect 13948 16346 13954 16348
rect 13708 16294 13710 16346
rect 13890 16294 13892 16346
rect 13646 16292 13652 16294
rect 13708 16292 13732 16294
rect 13788 16292 13812 16294
rect 13868 16292 13892 16294
rect 13948 16292 13954 16294
rect 13646 16283 13954 16292
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13556 15706 13584 15982
rect 13832 15706 13860 15982
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13924 15706 13952 15846
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14016 15502 14044 15846
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 14004 15496 14056 15502
rect 14200 15484 14228 18634
rect 14292 17270 14320 18838
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14384 18426 14412 18702
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14476 18086 14504 19858
rect 14568 18748 14596 20402
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14660 18970 14688 19790
rect 14936 19378 14964 23054
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 15028 21622 15056 22918
rect 15396 22710 15424 23598
rect 15476 23588 15528 23594
rect 15476 23530 15528 23536
rect 15384 22704 15436 22710
rect 15384 22646 15436 22652
rect 15396 21962 15424 22646
rect 15488 22642 15516 23530
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15580 22778 15608 23054
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15396 21690 15424 21898
rect 15948 21690 15976 23054
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 16040 21690 16068 22714
rect 16132 22522 16160 23684
rect 18156 23526 18184 24550
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 16820 23420 17128 23429
rect 16820 23418 16826 23420
rect 16882 23418 16906 23420
rect 16962 23418 16986 23420
rect 17042 23418 17066 23420
rect 17122 23418 17128 23420
rect 16882 23366 16884 23418
rect 17064 23366 17066 23418
rect 16820 23364 16826 23366
rect 16882 23364 16906 23366
rect 16962 23364 16986 23366
rect 17042 23364 17066 23366
rect 17122 23364 17128 23366
rect 16820 23355 17128 23364
rect 18156 23118 18184 23462
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 16488 23044 16540 23050
rect 16488 22986 16540 22992
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16224 22642 16252 22918
rect 16212 22636 16264 22642
rect 16264 22596 16436 22624
rect 16212 22578 16264 22584
rect 16132 22494 16252 22522
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16132 22234 16160 22374
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 15016 21616 15068 21622
rect 15016 21558 15068 21564
rect 16132 21536 16160 22170
rect 16224 22098 16252 22494
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 16408 21962 16436 22596
rect 16500 22234 16528 22986
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 16684 22642 16712 22918
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16580 22568 16632 22574
rect 16764 22568 16816 22574
rect 16580 22510 16632 22516
rect 16684 22516 16764 22522
rect 16684 22510 16816 22516
rect 16488 22228 16540 22234
rect 16488 22170 16540 22176
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16592 21622 16620 22510
rect 16684 22494 16804 22510
rect 16684 22030 16712 22494
rect 16820 22332 17128 22341
rect 16820 22330 16826 22332
rect 16882 22330 16906 22332
rect 16962 22330 16986 22332
rect 17042 22330 17066 22332
rect 17122 22330 17128 22332
rect 16882 22278 16884 22330
rect 17064 22278 17066 22330
rect 16820 22276 16826 22278
rect 16882 22276 16906 22278
rect 16962 22276 16986 22278
rect 17042 22276 17066 22278
rect 17122 22276 17128 22278
rect 16820 22267 17128 22276
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17328 21690 17356 21830
rect 17420 21690 17448 22918
rect 17696 21690 17724 22986
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 16580 21616 16632 21622
rect 17696 21593 17724 21626
rect 16580 21558 16632 21564
rect 16762 21584 16818 21593
rect 16212 21548 16264 21554
rect 16132 21508 16212 21536
rect 16212 21490 16264 21496
rect 16488 21072 16540 21078
rect 16488 21014 16540 21020
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15120 19854 15148 20538
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15304 20058 15332 20402
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14648 18760 14700 18766
rect 14568 18720 14648 18748
rect 14648 18702 14700 18708
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14568 17338 14596 17614
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16794 14412 16934
rect 14568 16794 14596 17002
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14660 16153 14688 18702
rect 14936 18630 14964 19314
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 17066 14872 17478
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14844 16522 14872 17002
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14844 16182 14872 16458
rect 14832 16176 14884 16182
rect 14646 16144 14702 16153
rect 14832 16118 14884 16124
rect 14646 16079 14702 16088
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14200 15456 14320 15484
rect 14004 15438 14056 15444
rect 13464 15094 13492 15438
rect 13646 15260 13954 15269
rect 13646 15258 13652 15260
rect 13708 15258 13732 15260
rect 13788 15258 13812 15260
rect 13868 15258 13892 15260
rect 13948 15258 13954 15260
rect 13708 15206 13710 15258
rect 13890 15206 13892 15258
rect 13646 15204 13652 15206
rect 13708 15204 13732 15206
rect 13788 15204 13812 15206
rect 13868 15204 13892 15206
rect 13948 15204 13954 15206
rect 13646 15195 13954 15204
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14328 13860 14962
rect 13832 14300 14044 14328
rect 13646 14172 13954 14181
rect 13646 14170 13652 14172
rect 13708 14170 13732 14172
rect 13788 14170 13812 14172
rect 13868 14170 13892 14172
rect 13948 14170 13954 14172
rect 13708 14118 13710 14170
rect 13890 14118 13892 14170
rect 13646 14116 13652 14118
rect 13708 14116 13732 14118
rect 13788 14116 13812 14118
rect 13868 14116 13892 14118
rect 13948 14116 13954 14118
rect 13646 14107 13954 14116
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 13924 13394 13952 13738
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13646 13084 13954 13093
rect 13646 13082 13652 13084
rect 13708 13082 13732 13084
rect 13788 13082 13812 13084
rect 13868 13082 13892 13084
rect 13948 13082 13954 13084
rect 13708 13030 13710 13082
rect 13890 13030 13892 13082
rect 13646 13028 13652 13030
rect 13708 13028 13732 13030
rect 13788 13028 13812 13030
rect 13868 13028 13892 13030
rect 13948 13028 13954 13030
rect 13646 13019 13954 13028
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11256 11898 11284 12106
rect 12728 11898 12756 12174
rect 13004 11898 13032 12174
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13188 11762 13216 12174
rect 13646 11996 13954 12005
rect 13646 11994 13652 11996
rect 13708 11994 13732 11996
rect 13788 11994 13812 11996
rect 13868 11994 13892 11996
rect 13948 11994 13954 11996
rect 13708 11942 13710 11994
rect 13890 11942 13892 11994
rect 13646 11940 13652 11942
rect 13708 11940 13732 11942
rect 13788 11940 13812 11942
rect 13868 11940 13892 11942
rect 13948 11940 13954 11942
rect 13646 11931 13954 11940
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13556 11082 13584 11698
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13646 10908 13954 10917
rect 13646 10906 13652 10908
rect 13708 10906 13732 10908
rect 13788 10906 13812 10908
rect 13868 10906 13892 10908
rect 13948 10906 13954 10908
rect 13708 10854 13710 10906
rect 13890 10854 13892 10906
rect 13646 10852 13652 10854
rect 13708 10852 13732 10854
rect 13788 10852 13812 10854
rect 13868 10852 13892 10854
rect 13948 10852 13954 10854
rect 13646 10843 13954 10852
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11072 9654 11100 10066
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10980 8974 11008 9386
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 9042 11376 9318
rect 11428 9104 11480 9110
rect 11428 9046 11480 9052
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 11072 8430 11100 8910
rect 11150 8800 11206 8809
rect 11150 8735 11206 8744
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11164 8362 11192 8735
rect 11440 8634 11468 9046
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11532 8430 11560 9930
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 8974 11744 9862
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11624 8566 11652 8774
rect 11808 8634 11836 9454
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10472 8188 10780 8197
rect 10472 8186 10478 8188
rect 10534 8186 10558 8188
rect 10614 8186 10638 8188
rect 10694 8186 10718 8188
rect 10774 8186 10780 8188
rect 10534 8134 10536 8186
rect 10716 8134 10718 8186
rect 10472 8132 10478 8134
rect 10534 8132 10558 8134
rect 10614 8132 10638 8134
rect 10694 8132 10718 8134
rect 10774 8132 10780 8134
rect 10472 8123 10780 8132
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10060 6798 10088 7278
rect 10472 7100 10780 7109
rect 10472 7098 10478 7100
rect 10534 7098 10558 7100
rect 10614 7098 10638 7100
rect 10694 7098 10718 7100
rect 10774 7098 10780 7100
rect 10534 7046 10536 7098
rect 10716 7046 10718 7098
rect 10472 7044 10478 7046
rect 10534 7044 10558 7046
rect 10614 7044 10638 7046
rect 10694 7044 10718 7046
rect 10774 7044 10780 7046
rect 10472 7035 10780 7044
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 8128 6310 8340 6338
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6380 3738 6408 4218
rect 6656 4214 6684 4558
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6656 3738 6684 4150
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6932 3466 6960 5714
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 5234 7144 5510
rect 7298 5468 7606 5477
rect 7298 5466 7304 5468
rect 7360 5466 7384 5468
rect 7440 5466 7464 5468
rect 7520 5466 7544 5468
rect 7600 5466 7606 5468
rect 7360 5414 7362 5466
rect 7542 5414 7544 5466
rect 7298 5412 7304 5414
rect 7360 5412 7384 5414
rect 7440 5412 7464 5414
rect 7520 5412 7544 5414
rect 7600 5412 7606 5414
rect 7298 5403 7606 5412
rect 7944 5234 7972 6190
rect 8036 6174 8248 6202
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5778 8156 6054
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7208 4282 7236 4626
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7298 4380 7606 4389
rect 7298 4378 7304 4380
rect 7360 4378 7384 4380
rect 7440 4378 7464 4380
rect 7520 4378 7544 4380
rect 7600 4378 7606 4380
rect 7360 4326 7362 4378
rect 7542 4326 7544 4378
rect 7298 4324 7304 4326
rect 7360 4324 7384 4326
rect 7440 4324 7464 4326
rect 7520 4324 7544 4326
rect 7600 4324 7606 4326
rect 7298 4315 7606 4324
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7668 4146 7696 4422
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6288 3126 6316 3334
rect 7024 3194 7052 3538
rect 7298 3292 7606 3301
rect 7298 3290 7304 3292
rect 7360 3290 7384 3292
rect 7440 3290 7464 3292
rect 7520 3290 7544 3292
rect 7600 3290 7606 3292
rect 7360 3238 7362 3290
rect 7542 3238 7544 3290
rect 7298 3236 7304 3238
rect 7360 3236 7384 3238
rect 7440 3236 7464 3238
rect 7520 3236 7544 3238
rect 7600 3236 7606 3238
rect 7298 3227 7606 3236
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7944 3126 7972 3878
rect 8128 3194 8156 5714
rect 8220 4758 8248 6174
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8220 4554 8248 4694
rect 8404 4690 8432 5238
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8220 3194 8248 3334
rect 8312 3194 8340 4422
rect 8404 3194 8432 4626
rect 8588 4078 8616 6054
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8680 4690 8708 5850
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8588 3466 8616 4014
rect 8772 3942 8800 6054
rect 9048 5914 9076 6598
rect 9692 6390 9720 6598
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 5914 9260 6190
rect 10244 6118 10272 6802
rect 10888 6458 10916 7890
rect 11900 7886 11928 8978
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8430 12020 8774
rect 12084 8498 12112 10406
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12176 8022 12204 8842
rect 12268 8362 12296 9454
rect 12256 8356 12308 8362
rect 12360 8344 12388 9862
rect 12438 9072 12494 9081
rect 12438 9007 12494 9016
rect 12452 8498 12480 9007
rect 12544 8838 12572 10610
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 9874 12756 10542
rect 12820 10130 12848 10678
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13188 10130 13216 10610
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12808 9920 12860 9926
rect 12728 9868 12808 9874
rect 12728 9862 12860 9868
rect 12728 9846 12848 9862
rect 12820 9178 12848 9846
rect 12912 9586 12940 9930
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12820 8974 12848 9114
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12912 8922 12940 9522
rect 13096 9450 13124 9998
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13096 9110 13124 9386
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 8566 12756 8774
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12716 8356 12768 8362
rect 12360 8316 12716 8344
rect 12256 8298 12308 8304
rect 12716 8298 12768 8304
rect 12820 8294 12848 8910
rect 12912 8894 13032 8922
rect 13096 8906 13124 9046
rect 12900 8832 12952 8838
rect 12898 8800 12900 8809
rect 12952 8800 12954 8809
rect 12898 8735 12954 8744
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11532 7274 11560 7754
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11164 6458 11192 6938
rect 11532 6866 11560 7210
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11532 6322 11560 6802
rect 11624 6458 11652 7142
rect 11992 7002 12020 7822
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12084 7546 12112 7686
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12268 7342 12296 7686
rect 12820 7546 12848 8230
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6458 11836 6598
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10472 6012 10780 6021
rect 10472 6010 10478 6012
rect 10534 6010 10558 6012
rect 10614 6010 10638 6012
rect 10694 6010 10718 6012
rect 10774 6010 10780 6012
rect 10534 5958 10536 6010
rect 10716 5958 10718 6010
rect 10472 5956 10478 5958
rect 10534 5956 10558 5958
rect 10614 5956 10638 5958
rect 10694 5956 10718 5958
rect 10774 5956 10780 5958
rect 10472 5947 10780 5956
rect 11808 5914 11836 6190
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 9508 5370 9536 5646
rect 9692 5370 9720 5646
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9692 4826 9720 5170
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 8772 3058 8800 3878
rect 8864 3738 8892 4558
rect 8956 4282 8984 4558
rect 10060 4282 10088 4762
rect 10336 4706 10364 5646
rect 11992 5302 12020 6938
rect 12268 6882 12296 7278
rect 12268 6854 12388 6882
rect 12452 6866 12480 7278
rect 12360 6730 12388 6854
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12360 5642 12388 6666
rect 12728 5846 12756 7414
rect 13004 7290 13032 8894
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8498 13124 8842
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13188 8022 13216 10066
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13280 8634 13308 9658
rect 13372 9081 13400 9862
rect 13646 9820 13954 9829
rect 13646 9818 13652 9820
rect 13708 9818 13732 9820
rect 13788 9818 13812 9820
rect 13868 9818 13892 9820
rect 13948 9818 13954 9820
rect 13708 9766 13710 9818
rect 13890 9766 13892 9818
rect 13646 9764 13652 9766
rect 13708 9764 13732 9766
rect 13788 9764 13812 9766
rect 13868 9764 13892 9766
rect 13948 9764 13954 9766
rect 13646 9755 13954 9764
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13358 9072 13414 9081
rect 13358 9007 13414 9016
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 13464 7954 13492 9454
rect 13646 8732 13954 8741
rect 13646 8730 13652 8732
rect 13708 8730 13732 8732
rect 13788 8730 13812 8732
rect 13868 8730 13892 8732
rect 13948 8730 13954 8732
rect 13708 8678 13710 8730
rect 13890 8678 13892 8730
rect 13646 8676 13652 8678
rect 13708 8676 13732 8678
rect 13788 8676 13812 8678
rect 13868 8676 13892 8678
rect 13948 8676 13954 8678
rect 13646 8667 13954 8676
rect 14016 8090 14044 14300
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14108 13870 14136 14214
rect 14200 13938 14228 14214
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14108 13546 14136 13806
rect 14108 13518 14228 13546
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14108 12850 14136 13126
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14200 12434 14228 13518
rect 14292 12442 14320 15456
rect 14568 15366 14596 15642
rect 14844 15570 14872 16118
rect 15028 15706 15056 17070
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14844 15434 14872 15506
rect 14832 15428 14884 15434
rect 14832 15370 14884 15376
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 15028 14618 15056 15642
rect 15120 14822 15148 19790
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15212 19174 15240 19654
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15212 18290 15240 19110
rect 15488 18426 15516 19246
rect 15948 18834 15976 20198
rect 16316 19854 16344 20878
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16500 19514 16528 21014
rect 16592 20890 16620 21558
rect 17682 21584 17738 21593
rect 16762 21519 16764 21528
rect 16816 21519 16818 21528
rect 17408 21548 17460 21554
rect 16764 21490 16816 21496
rect 17408 21490 17460 21496
rect 17592 21548 17644 21554
rect 17682 21519 17738 21528
rect 17592 21490 17644 21496
rect 17222 21448 17278 21457
rect 17222 21383 17224 21392
rect 17276 21383 17278 21392
rect 17224 21354 17276 21360
rect 17420 21332 17448 21490
rect 17500 21344 17552 21350
rect 17420 21304 17500 21332
rect 17500 21286 17552 21292
rect 16820 21244 17128 21253
rect 16820 21242 16826 21244
rect 16882 21242 16906 21244
rect 16962 21242 16986 21244
rect 17042 21242 17066 21244
rect 17122 21242 17128 21244
rect 16882 21190 16884 21242
rect 17064 21190 17066 21242
rect 16820 21188 16826 21190
rect 16882 21188 16906 21190
rect 16962 21188 16986 21190
rect 17042 21188 17066 21190
rect 17122 21188 17128 21190
rect 16820 21179 17128 21188
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17052 20942 17080 21014
rect 17040 20936 17092 20942
rect 16592 20862 16804 20890
rect 17040 20878 17092 20884
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16592 20534 16620 20742
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16592 20058 16620 20470
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16592 19310 16620 19722
rect 16684 19718 16712 20742
rect 16776 20534 16804 20862
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 16960 20641 16988 20810
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16946 20632 17002 20641
rect 16946 20567 17002 20576
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 17052 20244 17080 20742
rect 17144 20466 17172 21014
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17316 20256 17368 20262
rect 17052 20216 17264 20244
rect 16820 20156 17128 20165
rect 16820 20154 16826 20156
rect 16882 20154 16906 20156
rect 16962 20154 16986 20156
rect 17042 20154 17066 20156
rect 17122 20154 17128 20156
rect 16882 20102 16884 20154
rect 17064 20102 17066 20154
rect 16820 20100 16826 20102
rect 16882 20100 16906 20102
rect 16962 20100 16986 20102
rect 17042 20100 17066 20102
rect 17122 20100 17128 20102
rect 16820 20091 17128 20100
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 17236 19446 17264 20216
rect 17316 20198 17368 20204
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 16592 18766 16620 19246
rect 16820 19068 17128 19077
rect 16820 19066 16826 19068
rect 16882 19066 16906 19068
rect 16962 19066 16986 19068
rect 17042 19066 17066 19068
rect 17122 19066 17128 19068
rect 16882 19014 16884 19066
rect 17064 19014 17066 19066
rect 16820 19012 16826 19014
rect 16882 19012 16906 19014
rect 16962 19012 16986 19014
rect 17042 19012 17066 19014
rect 17122 19012 17128 19014
rect 16820 19003 17128 19012
rect 17328 18766 17356 20198
rect 17420 20058 17448 20402
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17512 19718 17540 21286
rect 17604 19718 17632 21490
rect 17788 20398 17816 21830
rect 17868 21548 17920 21554
rect 17972 21536 18000 22918
rect 18064 22438 18092 23054
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18064 21690 18092 22374
rect 18156 22234 18184 23054
rect 18248 22506 18276 23054
rect 18340 22710 18368 24686
rect 19536 24410 19564 25162
rect 19628 24410 19656 26318
rect 19720 25702 19748 26318
rect 19892 26240 19944 26246
rect 19892 26182 19944 26188
rect 19904 25702 19932 26182
rect 19994 26140 20302 26149
rect 19994 26138 20000 26140
rect 20056 26138 20080 26140
rect 20136 26138 20160 26140
rect 20216 26138 20240 26140
rect 20296 26138 20302 26140
rect 20056 26086 20058 26138
rect 20238 26086 20240 26138
rect 19994 26084 20000 26086
rect 20056 26084 20080 26086
rect 20136 26084 20160 26086
rect 20216 26084 20240 26086
rect 20296 26084 20302 26086
rect 19994 26075 20302 26084
rect 21100 25906 21128 26930
rect 21192 25906 21220 27066
rect 21456 26920 21508 26926
rect 21456 26862 21508 26868
rect 21640 26920 21692 26926
rect 21640 26862 21692 26868
rect 21824 26920 21876 26926
rect 21824 26862 21876 26868
rect 21468 26586 21496 26862
rect 21456 26580 21508 26586
rect 21456 26522 21508 26528
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 21284 25906 21312 26318
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 19708 25696 19760 25702
rect 19708 25638 19760 25644
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 19524 24404 19576 24410
rect 19524 24346 19576 24352
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 19720 24342 19748 25638
rect 19800 25220 19852 25226
rect 19800 25162 19852 25168
rect 19708 24336 19760 24342
rect 19708 24278 19760 24284
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 19076 23118 19104 23462
rect 19536 23254 19564 24210
rect 19812 24206 19840 25162
rect 19904 24886 19932 25638
rect 20364 25158 20392 25842
rect 20812 25832 20864 25838
rect 20732 25780 20812 25786
rect 21100 25786 21128 25842
rect 20864 25780 20944 25786
rect 20732 25758 20944 25780
rect 20732 25498 20760 25758
rect 20812 25696 20864 25702
rect 20812 25638 20864 25644
rect 20824 25498 20852 25638
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20916 25294 20944 25758
rect 21008 25758 21128 25786
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 19994 25052 20302 25061
rect 19994 25050 20000 25052
rect 20056 25050 20080 25052
rect 20136 25050 20160 25052
rect 20216 25050 20240 25052
rect 20296 25050 20302 25052
rect 20056 24998 20058 25050
rect 20238 24998 20240 25050
rect 19994 24996 20000 24998
rect 20056 24996 20080 24998
rect 20136 24996 20160 24998
rect 20216 24996 20240 24998
rect 20296 24996 20302 24998
rect 19994 24987 20302 24996
rect 19892 24880 19944 24886
rect 19892 24822 19944 24828
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 19904 24138 19932 24822
rect 20364 24698 20392 25094
rect 20536 24744 20588 24750
rect 20364 24692 20536 24698
rect 20364 24686 20588 24692
rect 20364 24670 20576 24686
rect 20076 24200 20128 24206
rect 20364 24188 20392 24670
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20548 24410 20576 24550
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20640 24274 20668 25230
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20128 24160 20392 24188
rect 20076 24142 20128 24148
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19800 24064 19852 24070
rect 19800 24006 19852 24012
rect 19524 23248 19576 23254
rect 19524 23190 19576 23196
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 18328 22704 18380 22710
rect 18328 22646 18380 22652
rect 19260 22642 19288 22918
rect 19812 22760 19840 24006
rect 19994 23964 20302 23973
rect 19994 23962 20000 23964
rect 20056 23962 20080 23964
rect 20136 23962 20160 23964
rect 20216 23962 20240 23964
rect 20296 23962 20302 23964
rect 20056 23910 20058 23962
rect 20238 23910 20240 23962
rect 19994 23908 20000 23910
rect 20056 23908 20080 23910
rect 20136 23908 20160 23910
rect 20216 23908 20240 23910
rect 20296 23908 20302 23910
rect 19994 23899 20302 23908
rect 20352 23656 20404 23662
rect 20352 23598 20404 23604
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19720 22732 19840 22760
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 18236 22500 18288 22506
rect 18236 22442 18288 22448
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 18052 21548 18104 21554
rect 17972 21508 18052 21536
rect 17868 21490 17920 21496
rect 18052 21490 18104 21496
rect 17880 21146 17908 21490
rect 18156 21434 18184 22034
rect 18248 21690 18276 22442
rect 19720 22094 19748 22732
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19812 22234 19840 22578
rect 19904 22234 19932 23122
rect 20364 23118 20392 23598
rect 20916 23322 20944 25230
rect 21008 25158 21036 25758
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 21100 25294 21128 25638
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 21100 24954 21128 25230
rect 21088 24948 21140 24954
rect 21088 24890 21140 24896
rect 21192 24750 21220 25842
rect 21468 25770 21496 26522
rect 21456 25764 21508 25770
rect 21456 25706 21508 25712
rect 21180 24744 21232 24750
rect 21180 24686 21232 24692
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 21652 23118 21680 26862
rect 21732 26240 21784 26246
rect 21732 26182 21784 26188
rect 21744 26042 21772 26182
rect 21836 26042 21864 26862
rect 22560 26852 22612 26858
rect 22560 26794 22612 26800
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 21732 26036 21784 26042
rect 21732 25978 21784 25984
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 21836 25906 21864 25978
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 21836 24596 21864 25842
rect 22008 24608 22060 24614
rect 21836 24568 22008 24596
rect 22008 24550 22060 24556
rect 21916 23248 21968 23254
rect 22112 23202 22140 26386
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22388 25498 22416 26318
rect 22468 26240 22520 26246
rect 22468 26182 22520 26188
rect 22480 25974 22508 26182
rect 22572 25974 22600 26794
rect 23168 26684 23476 26693
rect 23168 26682 23174 26684
rect 23230 26682 23254 26684
rect 23310 26682 23334 26684
rect 23390 26682 23414 26684
rect 23470 26682 23476 26684
rect 23230 26630 23232 26682
rect 23412 26630 23414 26682
rect 23168 26628 23174 26630
rect 23230 26628 23254 26630
rect 23310 26628 23334 26630
rect 23390 26628 23414 26630
rect 23470 26628 23476 26630
rect 23168 26619 23476 26628
rect 26342 26140 26650 26149
rect 26342 26138 26348 26140
rect 26404 26138 26428 26140
rect 26484 26138 26508 26140
rect 26564 26138 26588 26140
rect 26644 26138 26650 26140
rect 26404 26086 26406 26138
rect 26586 26086 26588 26138
rect 26342 26084 26348 26086
rect 26404 26084 26428 26086
rect 26484 26084 26508 26086
rect 26564 26084 26588 26086
rect 26644 26084 26650 26086
rect 26342 26075 26650 26084
rect 22468 25968 22520 25974
rect 22468 25910 22520 25916
rect 22560 25968 22612 25974
rect 22560 25910 22612 25916
rect 22744 25968 22796 25974
rect 22744 25910 22796 25916
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22388 24954 22416 25434
rect 22756 25294 22784 25910
rect 23168 25596 23476 25605
rect 23168 25594 23174 25596
rect 23230 25594 23254 25596
rect 23310 25594 23334 25596
rect 23390 25594 23414 25596
rect 23470 25594 23476 25596
rect 23230 25542 23232 25594
rect 23412 25542 23414 25594
rect 23168 25540 23174 25542
rect 23230 25540 23254 25542
rect 23310 25540 23334 25542
rect 23390 25540 23414 25542
rect 23470 25540 23476 25542
rect 23168 25531 23476 25540
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22296 23730 22324 24618
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 22388 23730 22416 24142
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22480 23798 22508 24006
rect 22468 23792 22520 23798
rect 22468 23734 22520 23740
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22296 23254 22324 23666
rect 21968 23196 22140 23202
rect 21916 23190 22140 23196
rect 22284 23248 22336 23254
rect 22284 23190 22336 23196
rect 21928 23174 22140 23190
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 19994 22876 20302 22885
rect 19994 22874 20000 22876
rect 20056 22874 20080 22876
rect 20136 22874 20160 22876
rect 20216 22874 20240 22876
rect 20296 22874 20302 22876
rect 20056 22822 20058 22874
rect 20238 22822 20240 22874
rect 19994 22820 20000 22822
rect 20056 22820 20080 22822
rect 20136 22820 20160 22822
rect 20216 22820 20240 22822
rect 20296 22820 20302 22822
rect 19994 22811 20302 22820
rect 20456 22778 20484 22918
rect 20444 22772 20496 22778
rect 20444 22714 20496 22720
rect 20824 22506 20852 23054
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 20812 22500 20864 22506
rect 20812 22442 20864 22448
rect 20996 22500 21048 22506
rect 20996 22442 21048 22448
rect 19800 22228 19852 22234
rect 19800 22170 19852 22176
rect 19892 22228 19944 22234
rect 19892 22170 19944 22176
rect 19720 22066 19932 22094
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18984 21690 19012 21830
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18972 21684 19024 21690
rect 18972 21626 19024 21632
rect 19904 21622 19932 22066
rect 19994 21788 20302 21797
rect 19994 21786 20000 21788
rect 20056 21786 20080 21788
rect 20136 21786 20160 21788
rect 20216 21786 20240 21788
rect 20296 21786 20302 21788
rect 20056 21734 20058 21786
rect 20238 21734 20240 21786
rect 19994 21732 20000 21734
rect 20056 21732 20080 21734
rect 20136 21732 20160 21734
rect 20216 21732 20240 21734
rect 20296 21732 20302 21734
rect 19994 21723 20302 21732
rect 19892 21616 19944 21622
rect 18326 21584 18382 21593
rect 18236 21548 18288 21554
rect 19892 21558 19944 21564
rect 20824 21554 20852 22442
rect 21008 22030 21036 22442
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21192 21962 21220 22374
rect 21284 22098 21312 22510
rect 21456 22500 21508 22506
rect 21456 22442 21508 22448
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 18326 21519 18328 21528
rect 18236 21490 18288 21496
rect 18380 21519 18382 21528
rect 20628 21548 20680 21554
rect 18328 21490 18380 21496
rect 20628 21490 20680 21496
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 18064 21418 18184 21434
rect 18052 21412 18184 21418
rect 18104 21406 18184 21412
rect 18052 21354 18104 21360
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 18156 20942 18184 21406
rect 18248 21146 18276 21490
rect 18602 21448 18658 21457
rect 18602 21383 18604 21392
rect 18656 21383 18658 21392
rect 18604 21354 18656 21360
rect 18236 21140 18288 21146
rect 18236 21082 18288 21088
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 17696 19854 17724 20198
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17512 19174 17540 19654
rect 18248 19258 18276 20742
rect 18340 20466 18368 20742
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18340 19378 18368 20402
rect 18432 19786 18460 20742
rect 18510 20632 18566 20641
rect 18510 20567 18512 20576
rect 18564 20567 18566 20576
rect 18512 20538 18564 20544
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18432 19378 18460 19722
rect 18524 19514 18552 20538
rect 18616 20466 18644 20878
rect 19994 20700 20302 20709
rect 19994 20698 20000 20700
rect 20056 20698 20080 20700
rect 20136 20698 20160 20700
rect 20216 20698 20240 20700
rect 20296 20698 20302 20700
rect 20056 20646 20058 20698
rect 20238 20646 20240 20698
rect 19994 20644 20000 20646
rect 20056 20644 20080 20646
rect 20136 20644 20160 20646
rect 20216 20644 20240 20646
rect 20296 20644 20302 20646
rect 19994 20635 20302 20644
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 18616 20058 18644 20402
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18984 19446 19012 19790
rect 18972 19440 19024 19446
rect 18972 19382 19024 19388
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18248 19242 18368 19258
rect 18248 19236 18380 19242
rect 18248 19230 18328 19236
rect 18328 19178 18380 19184
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 18432 18970 18460 19314
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 15660 18692 15712 18698
rect 15660 18634 15712 18640
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15672 17678 15700 18634
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15212 15366 15240 17138
rect 16592 17134 16620 18702
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 16820 17980 17128 17989
rect 16820 17978 16826 17980
rect 16882 17978 16906 17980
rect 16962 17978 16986 17980
rect 17042 17978 17066 17980
rect 17122 17978 17128 17980
rect 16882 17926 16884 17978
rect 17064 17926 17066 17978
rect 16820 17924 16826 17926
rect 16882 17924 16906 17926
rect 16962 17924 16986 17926
rect 17042 17924 17066 17926
rect 17122 17924 17128 17926
rect 16820 17915 17128 17924
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17236 17338 17264 17478
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 15292 17128 15344 17134
rect 16580 17128 16632 17134
rect 15292 17070 15344 17076
rect 15750 17096 15806 17105
rect 15304 15910 15332 17070
rect 16580 17070 16632 17076
rect 15750 17031 15806 17040
rect 15764 16998 15792 17031
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 13530 14504 13806
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14568 12986 14596 13670
rect 14660 13394 14688 14282
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14108 12406 14228 12434
rect 14280 12436 14332 12442
rect 14108 11762 14136 12406
rect 14280 12378 14332 12384
rect 14568 12306 14596 12922
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 11830 14228 12106
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11830 14504 12038
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14660 11762 14688 13330
rect 15120 11801 15148 14758
rect 15304 14482 15332 15846
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15488 14278 15516 16050
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15396 13530 15424 14010
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15212 12442 15240 13262
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15304 12322 15332 13262
rect 15212 12294 15332 12322
rect 15212 12170 15240 12294
rect 15488 12238 15516 14214
rect 15580 13938 15608 15506
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15580 13258 15608 13874
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15580 12918 15608 13194
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15106 11792 15162 11801
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14924 11756 14976 11762
rect 15106 11727 15162 11736
rect 15292 11756 15344 11762
rect 14924 11698 14976 11704
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14108 9450 14136 11562
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14200 11257 14228 11494
rect 14186 11248 14242 11257
rect 14186 11183 14242 11192
rect 14200 10606 14228 11183
rect 14464 11144 14516 11150
rect 14568 11121 14596 11494
rect 14464 11086 14516 11092
rect 14554 11112 14610 11121
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14096 9444 14148 9450
rect 14096 9386 14148 9392
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 9042 14228 9318
rect 14292 9042 14320 10406
rect 14476 9994 14504 11086
rect 14554 11047 14610 11056
rect 14660 10538 14688 11494
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14752 10674 14780 11086
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 13646 7644 13954 7653
rect 13646 7642 13652 7644
rect 13708 7642 13732 7644
rect 13788 7642 13812 7644
rect 13868 7642 13892 7644
rect 13948 7642 13954 7644
rect 13708 7590 13710 7642
rect 13890 7590 13892 7642
rect 13646 7588 13652 7590
rect 13708 7588 13732 7590
rect 13788 7588 13812 7590
rect 13868 7588 13892 7590
rect 13948 7588 13954 7590
rect 13646 7579 13954 7588
rect 14568 7546 14596 7686
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 12912 7262 13032 7290
rect 12912 7206 12940 7262
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 12912 6730 12940 7142
rect 14200 6866 14228 7142
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 12820 5234 12848 6054
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 10472 4924 10780 4933
rect 10472 4922 10478 4924
rect 10534 4922 10558 4924
rect 10614 4922 10638 4924
rect 10694 4922 10718 4924
rect 10774 4922 10780 4924
rect 10534 4870 10536 4922
rect 10716 4870 10718 4922
rect 10472 4868 10478 4870
rect 10534 4868 10558 4870
rect 10614 4868 10638 4870
rect 10694 4868 10718 4870
rect 10774 4868 10780 4870
rect 10472 4859 10780 4868
rect 12636 4826 12664 4966
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 10336 4678 10456 4706
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9232 3194 9260 3402
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9508 3126 9536 3334
rect 9784 3194 9812 3334
rect 9772 3188 9824 3194
rect 10152 3176 10180 3878
rect 10244 3534 10272 4218
rect 10336 4146 10364 4490
rect 10428 4146 10456 4678
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3602 10364 3878
rect 10472 3836 10780 3845
rect 10472 3834 10478 3836
rect 10534 3834 10558 3836
rect 10614 3834 10638 3836
rect 10694 3834 10718 3836
rect 10774 3834 10780 3836
rect 10534 3782 10536 3834
rect 10716 3782 10718 3834
rect 10472 3780 10478 3782
rect 10534 3780 10558 3782
rect 10614 3780 10638 3782
rect 10694 3780 10718 3782
rect 10774 3780 10780 3782
rect 10472 3771 10780 3780
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9772 3130 9824 3136
rect 10060 3148 10180 3176
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 3252 800 3280 2790
rect 4124 2748 4432 2757
rect 4124 2746 4130 2748
rect 4186 2746 4210 2748
rect 4266 2746 4290 2748
rect 4346 2746 4370 2748
rect 4426 2746 4432 2748
rect 4186 2694 4188 2746
rect 4368 2694 4370 2746
rect 4124 2692 4130 2694
rect 4186 2692 4210 2694
rect 4266 2692 4290 2694
rect 4346 2692 4370 2694
rect 4426 2692 4432 2694
rect 4124 2683 4432 2692
rect 9048 2650 9076 2926
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 10060 2514 10088 3148
rect 10244 2990 10272 3470
rect 10888 3194 10916 4082
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3466 11468 3878
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 10980 3194 11008 3402
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11532 3058 11560 3538
rect 11808 3194 11836 4422
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 3194 12848 3334
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12912 3058 12940 6666
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 13646 6556 13954 6565
rect 13646 6554 13652 6556
rect 13708 6554 13732 6556
rect 13788 6554 13812 6556
rect 13868 6554 13892 6556
rect 13948 6554 13954 6556
rect 13708 6502 13710 6554
rect 13890 6502 13892 6554
rect 13646 6500 13652 6502
rect 13708 6500 13732 6502
rect 13788 6500 13812 6502
rect 13868 6500 13892 6502
rect 13948 6500 13954 6502
rect 13646 6491 13954 6500
rect 14016 6458 14044 6598
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5914 13400 6054
rect 14108 5914 14136 6598
rect 14476 6458 14504 6598
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14660 5846 14688 6802
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4690 13032 4966
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13096 4570 13124 5646
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 13188 4758 13216 5510
rect 13646 5468 13954 5477
rect 13646 5466 13652 5468
rect 13708 5466 13732 5468
rect 13788 5466 13812 5468
rect 13868 5466 13892 5468
rect 13948 5466 13954 5468
rect 13708 5414 13710 5466
rect 13890 5414 13892 5466
rect 13646 5412 13652 5414
rect 13708 5412 13732 5414
rect 13788 5412 13812 5414
rect 13868 5412 13892 5414
rect 13948 5412 13954 5414
rect 13646 5403 13954 5412
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13280 4826 13308 4966
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13176 4752 13228 4758
rect 13372 4706 13400 4966
rect 13464 4758 13492 5034
rect 13176 4694 13228 4700
rect 13004 4554 13124 4570
rect 12992 4548 13124 4554
rect 13044 4542 13124 4548
rect 13280 4678 13400 4706
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 12992 4490 13044 4496
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 3534 13124 4422
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13188 4078 13216 4150
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13280 3534 13308 4678
rect 13556 4622 13584 5034
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 14004 4616 14056 4622
rect 14200 4604 14228 4966
rect 14384 4826 14412 5170
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14280 4616 14332 4622
rect 14056 4576 14136 4604
rect 14004 4558 14056 4564
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 13280 2922 13308 3470
rect 13372 3126 13400 4490
rect 13464 3398 13492 4558
rect 13556 4282 13584 4558
rect 14108 4486 14136 4576
rect 14200 4576 14280 4604
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13646 4380 13954 4389
rect 13646 4378 13652 4380
rect 13708 4378 13732 4380
rect 13788 4378 13812 4380
rect 13868 4378 13892 4380
rect 13948 4378 13954 4380
rect 13708 4326 13710 4378
rect 13890 4326 13892 4378
rect 13646 4324 13652 4326
rect 13708 4324 13732 4326
rect 13788 4324 13812 4326
rect 13868 4324 13892 4326
rect 13948 4324 13954 4326
rect 13646 4315 13954 4324
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 14016 4214 14044 4422
rect 13912 4208 13964 4214
rect 13910 4176 13912 4185
rect 14004 4208 14056 4214
rect 13964 4176 13966 4185
rect 14004 4150 14056 4156
rect 13910 4111 13966 4120
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13832 3602 13860 3946
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 14108 3466 14136 4422
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13360 3120 13412 3126
rect 13358 3088 13360 3097
rect 13412 3088 13414 3097
rect 13358 3023 13414 3032
rect 13464 2972 13492 3334
rect 13646 3292 13954 3301
rect 13646 3290 13652 3292
rect 13708 3290 13732 3292
rect 13788 3290 13812 3292
rect 13868 3290 13892 3292
rect 13948 3290 13954 3292
rect 13708 3238 13710 3290
rect 13890 3238 13892 3290
rect 13646 3236 13652 3238
rect 13708 3236 13732 3238
rect 13788 3236 13812 3238
rect 13868 3236 13892 3238
rect 13948 3236 13954 3238
rect 13646 3227 13954 3236
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13832 2972 13860 3130
rect 13464 2944 13860 2972
rect 14016 2922 14044 3402
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 14004 2916 14056 2922
rect 14004 2858 14056 2864
rect 10472 2748 10780 2757
rect 10472 2746 10478 2748
rect 10534 2746 10558 2748
rect 10614 2746 10638 2748
rect 10694 2746 10718 2748
rect 10774 2746 10780 2748
rect 10534 2694 10536 2746
rect 10716 2694 10718 2746
rect 10472 2692 10478 2694
rect 10534 2692 10558 2694
rect 10614 2692 10638 2694
rect 10694 2692 10718 2694
rect 10774 2692 10780 2694
rect 10472 2683 10780 2692
rect 14108 2582 14136 3402
rect 14200 2990 14228 4576
rect 14280 4558 14332 4564
rect 14372 4208 14424 4214
rect 14476 4196 14504 5510
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14660 4622 14688 5034
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14424 4168 14596 4196
rect 14372 4150 14424 4156
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14280 3664 14332 3670
rect 14280 3606 14332 3612
rect 14292 3058 14320 3606
rect 14384 3466 14412 4014
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14476 3398 14504 3946
rect 14464 3392 14516 3398
rect 14462 3360 14464 3369
rect 14516 3360 14518 3369
rect 14462 3295 14518 3304
rect 14568 3126 14596 4168
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14752 2650 14780 4490
rect 14844 3602 14872 8774
rect 14936 8634 14964 11698
rect 15120 9110 15148 11727
rect 15292 11698 15344 11704
rect 15304 11642 15332 11698
rect 15212 11614 15332 11642
rect 15212 11354 15240 11614
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15304 11014 15332 11494
rect 15488 11234 15516 11834
rect 15580 11762 15608 12038
rect 15672 11898 15700 12310
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15396 11206 15516 11234
rect 15580 11218 15608 11494
rect 15568 11212 15620 11218
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15212 9518 15240 10950
rect 15396 10742 15424 11206
rect 15568 11154 15620 11160
rect 15476 11076 15528 11082
rect 15528 11036 15608 11064
rect 15476 11018 15528 11024
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15580 10674 15608 11036
rect 15672 10810 15700 11494
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15384 10532 15436 10538
rect 15384 10474 15436 10480
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15304 9382 15332 9862
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15396 8634 15424 10474
rect 15488 9178 15516 10610
rect 15580 10538 15608 10610
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10266 15608 10474
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15764 9602 15792 16934
rect 16592 16658 16620 17070
rect 16820 16892 17128 16901
rect 16820 16890 16826 16892
rect 16882 16890 16906 16892
rect 16962 16890 16986 16892
rect 17042 16890 17066 16892
rect 17122 16890 17128 16892
rect 16882 16838 16884 16890
rect 17064 16838 17066 16890
rect 16820 16836 16826 16838
rect 16882 16836 16906 16838
rect 16962 16836 16986 16838
rect 17042 16836 17066 16838
rect 17122 16836 17128 16838
rect 16820 16827 17128 16836
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16210 16144 16266 16153
rect 16592 16114 16620 16594
rect 17512 16522 17540 18634
rect 18984 18290 19012 19382
rect 19352 19310 19380 20402
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20272 19718 20300 20198
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 19994 19612 20302 19621
rect 19994 19610 20000 19612
rect 20056 19610 20080 19612
rect 20136 19610 20160 19612
rect 20216 19610 20240 19612
rect 20296 19610 20302 19612
rect 20056 19558 20058 19610
rect 20238 19558 20240 19610
rect 19994 19556 20000 19558
rect 20056 19556 20080 19558
rect 20136 19556 20160 19558
rect 20216 19556 20240 19558
rect 20296 19556 20302 19558
rect 19994 19547 20302 19556
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19812 19242 19932 19258
rect 19800 19236 19932 19242
rect 19852 19230 19932 19236
rect 19800 19178 19852 19184
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17338 18460 17478
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17512 16182 17540 16458
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 16210 16079 16266 16088
rect 16396 16108 16448 16114
rect 16224 15978 16252 16079
rect 16396 16050 16448 16056
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16408 14618 16436 16050
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16684 15706 16712 15914
rect 16820 15804 17128 15813
rect 16820 15802 16826 15804
rect 16882 15802 16906 15804
rect 16962 15802 16986 15804
rect 17042 15802 17066 15804
rect 17122 15802 17128 15804
rect 16882 15750 16884 15802
rect 17064 15750 17066 15802
rect 16820 15748 16826 15750
rect 16882 15748 16906 15750
rect 16962 15748 16986 15750
rect 17042 15748 17066 15750
rect 17122 15748 17128 15750
rect 16820 15739 17128 15748
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 18340 15570 18368 16526
rect 18432 16114 18460 17274
rect 18616 16726 18644 17614
rect 18694 17232 18750 17241
rect 18694 17167 18696 17176
rect 18748 17167 18750 17176
rect 18696 17138 18748 17144
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18708 16658 18736 16934
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18800 16590 18828 17614
rect 18892 17338 18920 17614
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18984 17134 19012 18226
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 19076 17338 19104 17478
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19062 17232 19118 17241
rect 19352 17218 19380 18838
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19720 18426 19748 18566
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19118 17190 19380 17218
rect 19062 17167 19118 17176
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18972 17128 19024 17134
rect 19248 17128 19300 17134
rect 18972 17070 19024 17076
rect 19246 17096 19248 17105
rect 19300 17096 19302 17105
rect 18892 16998 18920 17070
rect 19246 17031 19302 17040
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16658 19380 16934
rect 19904 16674 19932 19230
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 19994 18524 20302 18533
rect 19994 18522 20000 18524
rect 20056 18522 20080 18524
rect 20136 18522 20160 18524
rect 20216 18522 20240 18524
rect 20296 18522 20302 18524
rect 20056 18470 20058 18522
rect 20238 18470 20240 18522
rect 19994 18468 20000 18470
rect 20056 18468 20080 18470
rect 20136 18468 20160 18470
rect 20216 18468 20240 18470
rect 20296 18468 20302 18470
rect 19994 18459 20302 18468
rect 19994 17436 20302 17445
rect 19994 17434 20000 17436
rect 20056 17434 20080 17436
rect 20136 17434 20160 17436
rect 20216 17434 20240 17436
rect 20296 17434 20302 17436
rect 20056 17382 20058 17434
rect 20238 17382 20240 17434
rect 19994 17380 20000 17382
rect 20056 17380 20080 17382
rect 20136 17380 20160 17382
rect 20216 17380 20240 17382
rect 20296 17380 20302 17382
rect 19994 17371 20302 17380
rect 20364 17354 20392 18702
rect 20548 18290 20576 20402
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20548 17678 20576 18226
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20364 17326 20484 17354
rect 20456 16794 20484 17326
rect 20548 17270 20576 17614
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20640 17134 20668 21490
rect 21376 20942 21404 21898
rect 21468 21554 21496 22442
rect 21652 22030 21680 23054
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20824 20058 20852 20198
rect 20916 20058 20944 20402
rect 21652 20330 21680 21966
rect 21928 21690 21956 22986
rect 22020 22710 22048 23174
rect 22296 23118 22324 23190
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 22112 21554 22140 23054
rect 22192 23044 22244 23050
rect 22192 22986 22244 22992
rect 22204 22438 22232 22986
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22296 22778 22324 22918
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22282 22672 22338 22681
rect 22388 22658 22416 23666
rect 22756 23662 22784 25230
rect 26342 25052 26650 25061
rect 26342 25050 26348 25052
rect 26404 25050 26428 25052
rect 26484 25050 26508 25052
rect 26564 25050 26588 25052
rect 26644 25050 26650 25052
rect 26404 24998 26406 25050
rect 26586 24998 26588 25050
rect 26342 24996 26348 24998
rect 26404 24996 26428 24998
rect 26484 24996 26508 24998
rect 26564 24996 26588 24998
rect 26644 24996 26650 24998
rect 26342 24987 26650 24996
rect 23020 24676 23072 24682
rect 23020 24618 23072 24624
rect 23032 24290 23060 24618
rect 23168 24508 23476 24517
rect 23168 24506 23174 24508
rect 23230 24506 23254 24508
rect 23310 24506 23334 24508
rect 23390 24506 23414 24508
rect 23470 24506 23476 24508
rect 23230 24454 23232 24506
rect 23412 24454 23414 24506
rect 23168 24452 23174 24454
rect 23230 24452 23254 24454
rect 23310 24452 23334 24454
rect 23390 24452 23414 24454
rect 23470 24452 23476 24454
rect 23168 24443 23476 24452
rect 23032 24262 23152 24290
rect 23124 24206 23152 24262
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22652 23248 22704 23254
rect 22652 23190 22704 23196
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22480 22778 22508 22918
rect 22572 22778 22600 23054
rect 22468 22772 22520 22778
rect 22468 22714 22520 22720
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22338 22630 22416 22658
rect 22282 22607 22284 22616
rect 22336 22607 22338 22616
rect 22284 22578 22336 22584
rect 22664 22574 22692 23190
rect 22756 23118 22784 23598
rect 22744 23112 22796 23118
rect 22744 23054 22796 23060
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22664 21690 22692 22510
rect 22756 22234 22784 23054
rect 22928 23044 22980 23050
rect 22928 22986 22980 22992
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 22848 22642 22876 22918
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22940 22234 22968 22986
rect 22744 22228 22796 22234
rect 22744 22170 22796 22176
rect 22928 22228 22980 22234
rect 22928 22170 22980 22176
rect 23032 22094 23060 24142
rect 23308 23866 23336 24142
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23168 23420 23476 23429
rect 23168 23418 23174 23420
rect 23230 23418 23254 23420
rect 23310 23418 23334 23420
rect 23390 23418 23414 23420
rect 23470 23418 23476 23420
rect 23230 23366 23232 23418
rect 23412 23366 23414 23418
rect 23168 23364 23174 23366
rect 23230 23364 23254 23366
rect 23310 23364 23334 23366
rect 23390 23364 23414 23366
rect 23470 23364 23476 23366
rect 23168 23355 23476 23364
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23110 22672 23166 22681
rect 23110 22607 23166 22616
rect 23124 22574 23152 22607
rect 23308 22574 23336 23258
rect 23584 22778 23612 23802
rect 26160 23769 26188 24142
rect 26342 23964 26650 23973
rect 26342 23962 26348 23964
rect 26404 23962 26428 23964
rect 26484 23962 26508 23964
rect 26564 23962 26588 23964
rect 26644 23962 26650 23964
rect 26404 23910 26406 23962
rect 26586 23910 26588 23962
rect 26342 23908 26348 23910
rect 26404 23908 26428 23910
rect 26484 23908 26508 23910
rect 26564 23908 26588 23910
rect 26644 23908 26650 23910
rect 26342 23899 26650 23908
rect 26146 23760 26202 23769
rect 24768 23724 24820 23730
rect 26146 23695 26202 23704
rect 24768 23666 24820 23672
rect 24780 23202 24808 23666
rect 24596 23186 24808 23202
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 24596 23180 24820 23186
rect 24596 23174 24768 23180
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23676 22778 23704 22918
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 24044 22710 24072 23122
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24032 22704 24084 22710
rect 24032 22646 24084 22652
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23112 22568 23164 22574
rect 23112 22510 23164 22516
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 23168 22332 23476 22341
rect 23168 22330 23174 22332
rect 23230 22330 23254 22332
rect 23310 22330 23334 22332
rect 23390 22330 23414 22332
rect 23470 22330 23476 22332
rect 23230 22278 23232 22330
rect 23412 22278 23414 22330
rect 23168 22276 23174 22278
rect 23230 22276 23254 22278
rect 23310 22276 23334 22278
rect 23390 22276 23414 22278
rect 23470 22276 23476 22278
rect 23168 22267 23476 22276
rect 22940 22066 23060 22094
rect 22940 21894 22968 22066
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22020 21146 22048 21490
rect 22560 21412 22612 21418
rect 22560 21354 22612 21360
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22112 20534 22140 21286
rect 22572 20942 22600 21354
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20916 19446 20944 19994
rect 21652 19514 21680 20266
rect 22204 20262 22232 20810
rect 22572 20466 22600 20878
rect 22756 20806 22784 20878
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22756 20602 22784 20742
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22204 19922 22232 20198
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 22204 19378 22232 19858
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22756 19514 22784 19722
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20732 17338 20760 18702
rect 22204 18290 22232 19314
rect 22848 19310 22876 21286
rect 22940 20942 22968 21830
rect 23676 21690 23704 21898
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23168 21244 23476 21253
rect 23168 21242 23174 21244
rect 23230 21242 23254 21244
rect 23310 21242 23334 21244
rect 23390 21242 23414 21244
rect 23470 21242 23476 21244
rect 23230 21190 23232 21242
rect 23412 21190 23414 21242
rect 23168 21188 23174 21190
rect 23230 21188 23254 21190
rect 23310 21188 23334 21190
rect 23390 21188 23414 21190
rect 23470 21188 23476 21190
rect 23168 21179 23476 21188
rect 23204 21140 23256 21146
rect 23584 21128 23612 21422
rect 23204 21082 23256 21088
rect 23400 21100 23612 21128
rect 23216 20942 23244 21082
rect 23400 20942 23428 21100
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 22940 20398 22968 20878
rect 23216 20466 23244 20878
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 23400 20330 23428 20878
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 23492 20262 23520 20470
rect 23584 20398 23612 20878
rect 23676 20602 23704 21490
rect 23768 20806 23796 22578
rect 24136 22098 24164 22918
rect 24228 22778 24532 22794
rect 24216 22772 24544 22778
rect 24268 22766 24492 22772
rect 24216 22714 24268 22720
rect 24492 22714 24544 22720
rect 24400 22704 24452 22710
rect 24596 22658 24624 23174
rect 24768 23122 24820 23128
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 25320 23112 25372 23118
rect 25320 23054 25372 23060
rect 24452 22652 24624 22658
rect 24400 22646 24624 22652
rect 24412 22630 24624 22646
rect 24688 22522 24716 23054
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24964 22710 24992 22986
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 24952 22704 25004 22710
rect 24952 22646 25004 22652
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24504 22506 24716 22522
rect 24492 22500 24716 22506
rect 24544 22494 24716 22500
rect 24492 22442 24544 22448
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 24780 22030 24808 22374
rect 24872 22234 24900 22578
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 25148 22098 25176 22918
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23664 20460 23716 20466
rect 23768 20448 23796 20742
rect 23952 20602 23980 21490
rect 24044 21418 24072 21966
rect 24780 21690 24808 21966
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24032 21412 24084 21418
rect 24032 21354 24084 21360
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 23716 20420 23796 20448
rect 23664 20402 23716 20408
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23168 20156 23476 20165
rect 23168 20154 23174 20156
rect 23230 20154 23254 20156
rect 23310 20154 23334 20156
rect 23390 20154 23414 20156
rect 23470 20154 23476 20156
rect 23230 20102 23232 20154
rect 23412 20102 23414 20154
rect 23168 20100 23174 20102
rect 23230 20100 23254 20102
rect 23310 20100 23334 20102
rect 23390 20100 23414 20102
rect 23470 20100 23476 20102
rect 23168 20091 23476 20100
rect 23584 20058 23612 20334
rect 24136 20262 24164 21490
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24228 20942 24256 21286
rect 24216 20936 24268 20942
rect 24216 20878 24268 20884
rect 25148 20714 25176 22034
rect 25332 21690 25360 23054
rect 26342 22876 26650 22885
rect 26342 22874 26348 22876
rect 26404 22874 26428 22876
rect 26484 22874 26508 22876
rect 26564 22874 26588 22876
rect 26644 22874 26650 22876
rect 26404 22822 26406 22874
rect 26586 22822 26588 22874
rect 26342 22820 26348 22822
rect 26404 22820 26428 22822
rect 26484 22820 26508 22822
rect 26564 22820 26588 22822
rect 26644 22820 26650 22822
rect 26342 22811 26650 22820
rect 25780 22772 25832 22778
rect 25780 22714 25832 22720
rect 25792 22098 25820 22714
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25320 21684 25372 21690
rect 25320 21626 25372 21632
rect 25792 21554 25820 22034
rect 26342 21788 26650 21797
rect 26342 21786 26348 21788
rect 26404 21786 26428 21788
rect 26484 21786 26508 21788
rect 26564 21786 26588 21788
rect 26644 21786 26650 21788
rect 26404 21734 26406 21786
rect 26586 21734 26588 21786
rect 26342 21732 26348 21734
rect 26404 21732 26428 21734
rect 26484 21732 26508 21734
rect 26564 21732 26588 21734
rect 26644 21732 26650 21734
rect 26342 21723 26650 21732
rect 25780 21548 25832 21554
rect 25780 21490 25832 21496
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25332 21146 25360 21422
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 24964 20686 25176 20714
rect 26342 20700 26650 20709
rect 26342 20698 26348 20700
rect 26404 20698 26428 20700
rect 26484 20698 26508 20700
rect 26564 20698 26588 20700
rect 26644 20698 26650 20700
rect 24964 20602 24992 20686
rect 26404 20646 26406 20698
rect 26586 20646 26588 20698
rect 26342 20644 26348 20646
rect 26404 20644 26428 20646
rect 26484 20644 26508 20646
rect 26564 20644 26588 20646
rect 26644 20644 26650 20646
rect 26342 20635 26650 20644
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23676 19378 23704 20198
rect 26342 19612 26650 19621
rect 26342 19610 26348 19612
rect 26404 19610 26428 19612
rect 26484 19610 26508 19612
rect 26564 19610 26588 19612
rect 26644 19610 26650 19612
rect 26404 19558 26406 19610
rect 26586 19558 26588 19610
rect 26342 19556 26348 19558
rect 26404 19556 26428 19558
rect 26484 19556 26508 19558
rect 26564 19556 26588 19558
rect 26644 19556 26650 19558
rect 26342 19547 26650 19556
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 23168 19068 23476 19077
rect 23168 19066 23174 19068
rect 23230 19066 23254 19068
rect 23310 19066 23334 19068
rect 23390 19066 23414 19068
rect 23470 19066 23476 19068
rect 23230 19014 23232 19066
rect 23412 19014 23414 19066
rect 23168 19012 23174 19014
rect 23230 19012 23254 19014
rect 23310 19012 23334 19014
rect 23390 19012 23414 19014
rect 23470 19012 23476 19014
rect 23168 19003 23476 19012
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22008 18216 22060 18222
rect 22008 18158 22060 18164
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20732 16794 20760 17274
rect 20916 17202 20944 18022
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21100 17542 21128 17682
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20824 16726 20852 16934
rect 20812 16720 20864 16726
rect 19340 16652 19392 16658
rect 19904 16646 20392 16674
rect 20812 16662 20864 16668
rect 19340 16594 19392 16600
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19260 16250 19288 16526
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18524 15706 18552 15846
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18616 15502 18644 16186
rect 19536 16114 19564 16390
rect 19812 16250 19840 16526
rect 19904 16250 19932 16526
rect 19994 16348 20302 16357
rect 19994 16346 20000 16348
rect 20056 16346 20080 16348
rect 20136 16346 20160 16348
rect 20216 16346 20240 16348
rect 20296 16346 20302 16348
rect 20056 16294 20058 16346
rect 20238 16294 20240 16346
rect 19994 16292 20000 16294
rect 20056 16292 20080 16294
rect 20136 16292 20160 16294
rect 20216 16292 20240 16294
rect 20296 16292 20302 16294
rect 19994 16283 20302 16292
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 16820 14716 17128 14725
rect 16820 14714 16826 14716
rect 16882 14714 16906 14716
rect 16962 14714 16986 14716
rect 17042 14714 17066 14716
rect 17122 14714 17128 14716
rect 16882 14662 16884 14714
rect 17064 14662 17066 14714
rect 16820 14660 16826 14662
rect 16882 14660 16906 14662
rect 16962 14660 16986 14662
rect 17042 14660 17066 14662
rect 17122 14660 17128 14662
rect 16820 14651 17128 14660
rect 17420 14618 17448 14894
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 14074 15976 14350
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16684 14074 16712 14214
rect 16868 14074 16896 14214
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 16820 13628 17128 13637
rect 16820 13626 16826 13628
rect 16882 13626 16906 13628
rect 16962 13626 16986 13628
rect 17042 13626 17066 13628
rect 17122 13626 17128 13628
rect 16882 13574 16884 13626
rect 17064 13574 17066 13626
rect 16820 13572 16826 13574
rect 16882 13572 16906 13574
rect 16962 13572 16986 13574
rect 17042 13572 17066 13574
rect 17122 13572 17128 13574
rect 16820 13563 17128 13572
rect 17328 13394 17356 13670
rect 17512 13394 17540 15098
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17604 13734 17632 14350
rect 17972 13938 18000 15030
rect 18432 14550 18460 15370
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17604 13462 17632 13670
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17316 13388 17368 13394
rect 17500 13388 17552 13394
rect 17316 13330 17368 13336
rect 17420 13348 17500 13376
rect 17420 12918 17448 13348
rect 17500 13330 17552 13336
rect 17972 12986 18000 13874
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13530 18092 13806
rect 18432 13530 18460 14486
rect 18800 14414 18828 15302
rect 19260 15162 19288 15438
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18892 14618 18920 14894
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 19260 14074 19288 15098
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19352 14618 19380 14962
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19352 13802 19380 14214
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19248 13728 19300 13734
rect 19300 13676 19380 13682
rect 19248 13670 19380 13676
rect 19260 13654 19380 13670
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19260 12986 19288 13126
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 16820 12540 17128 12549
rect 16820 12538 16826 12540
rect 16882 12538 16906 12540
rect 16962 12538 16986 12540
rect 17042 12538 17066 12540
rect 17122 12538 17128 12540
rect 16882 12486 16884 12538
rect 17064 12486 17066 12538
rect 16820 12484 16826 12486
rect 16882 12484 16906 12486
rect 16962 12484 16986 12486
rect 17042 12484 17066 12486
rect 17122 12484 17128 12486
rect 16820 12475 17128 12484
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15856 11257 15884 11290
rect 15842 11248 15898 11257
rect 15842 11183 15898 11192
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 10266 15884 10406
rect 15948 10266 15976 11698
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16040 11286 16068 11494
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16316 11082 16344 12038
rect 16408 11830 16436 12174
rect 17420 11830 17448 12854
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19260 12238 19288 12378
rect 19352 12306 19380 13654
rect 19444 13376 19472 15846
rect 19536 14346 19564 16050
rect 19904 15570 19932 16186
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19628 14414 19656 15370
rect 19994 15260 20302 15269
rect 19994 15258 20000 15260
rect 20056 15258 20080 15260
rect 20136 15258 20160 15260
rect 20216 15258 20240 15260
rect 20296 15258 20302 15260
rect 20056 15206 20058 15258
rect 20238 15206 20240 15258
rect 19994 15204 20000 15206
rect 20056 15204 20080 15206
rect 20136 15204 20160 15206
rect 20216 15204 20240 15206
rect 20296 15204 20302 15206
rect 19994 15195 20302 15204
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19904 13870 19932 14758
rect 19994 14172 20302 14181
rect 19994 14170 20000 14172
rect 20056 14170 20080 14172
rect 20136 14170 20160 14172
rect 20216 14170 20240 14172
rect 20296 14170 20302 14172
rect 20056 14118 20058 14170
rect 20238 14118 20240 14170
rect 19994 14116 20000 14118
rect 20056 14116 20080 14118
rect 20136 14116 20160 14118
rect 20216 14116 20240 14118
rect 20296 14116 20302 14118
rect 19994 14107 20302 14116
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19524 13388 19576 13394
rect 19444 13348 19524 13376
rect 19444 12782 19472 13348
rect 19524 13330 19576 13336
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19812 12238 19840 13126
rect 19904 12306 19932 13806
rect 19994 13084 20302 13093
rect 19994 13082 20000 13084
rect 20056 13082 20080 13084
rect 20136 13082 20160 13084
rect 20216 13082 20240 13084
rect 20296 13082 20302 13084
rect 20056 13030 20058 13082
rect 20238 13030 20240 13082
rect 19994 13028 20000 13030
rect 20056 13028 20080 13030
rect 20136 13028 20160 13030
rect 20216 13028 20240 13030
rect 20296 13028 20302 13030
rect 19994 13019 20302 13028
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 16396 11824 16448 11830
rect 16396 11766 16448 11772
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17958 11792 18014 11801
rect 16408 11354 16436 11766
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16500 11082 16528 11630
rect 16820 11452 17128 11461
rect 16820 11450 16826 11452
rect 16882 11450 16906 11452
rect 16962 11450 16986 11452
rect 17042 11450 17066 11452
rect 17122 11450 17128 11452
rect 16882 11398 16884 11450
rect 17064 11398 17066 11450
rect 16820 11396 16826 11398
rect 16882 11396 16906 11398
rect 16962 11396 16986 11398
rect 17042 11396 17066 11398
rect 17122 11396 17128 11398
rect 16820 11387 17128 11396
rect 17236 11082 17264 11698
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 16316 10606 16344 11018
rect 16500 10810 16528 11018
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 15764 9574 15884 9602
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15120 5370 15148 8434
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15212 6934 15240 7890
rect 15304 7886 15332 8230
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14936 3738 14964 4558
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 15028 4146 15056 4422
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14936 3466 14964 3674
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 14844 2922 14872 3402
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14936 2514 14964 3402
rect 15120 3126 15148 5034
rect 15212 4185 15240 6054
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15304 5098 15332 5510
rect 15580 5234 15608 5510
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15396 4826 15424 5170
rect 15672 4842 15700 7754
rect 15856 6730 15884 9574
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15948 8634 15976 8774
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16040 8566 16068 9522
rect 16132 9518 16160 9998
rect 16316 9994 16344 10542
rect 16408 10266 16436 10610
rect 16500 10470 16528 10746
rect 16684 10674 16712 11018
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 17236 10470 17264 11018
rect 17420 10674 17448 11766
rect 17958 11727 17960 11736
rect 18012 11727 18014 11736
rect 17960 11698 18012 11704
rect 17972 11354 18000 11698
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17880 10742 17908 11154
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16500 10130 16528 10406
rect 16820 10364 17128 10373
rect 16820 10362 16826 10364
rect 16882 10362 16906 10364
rect 16962 10362 16986 10364
rect 17042 10362 17066 10364
rect 17122 10362 17128 10364
rect 16882 10310 16884 10362
rect 17064 10310 17066 10362
rect 16820 10308 16826 10310
rect 16882 10308 16906 10310
rect 16962 10308 16986 10310
rect 17042 10308 17066 10310
rect 17122 10308 17128 10310
rect 16820 10299 17128 10308
rect 17236 10130 17264 10406
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16132 9042 16160 9454
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 16820 9276 17128 9285
rect 16820 9274 16826 9276
rect 16882 9274 16906 9276
rect 16962 9274 16986 9276
rect 17042 9274 17066 9276
rect 17122 9274 17128 9276
rect 16882 9222 16884 9274
rect 17064 9222 17066 9274
rect 16820 9220 16826 9222
rect 16882 9220 16906 9222
rect 16962 9220 16986 9222
rect 17042 9220 17066 9222
rect 17122 9220 17128 9222
rect 16820 9211 17128 9220
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 16040 7546 16068 8502
rect 16132 8362 16160 8978
rect 17880 8906 17908 9318
rect 17972 8974 18000 11290
rect 18064 10470 18092 11630
rect 18156 11218 18184 11834
rect 18696 11824 18748 11830
rect 18696 11766 18748 11772
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18248 11286 18276 11494
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10062 18092 10406
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18156 9926 18184 11154
rect 18524 11150 18552 11630
rect 18708 11286 18736 11766
rect 18696 11280 18748 11286
rect 19352 11234 19380 12038
rect 19536 11898 19564 12174
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19628 11762 19656 12174
rect 19720 12102 19748 12174
rect 20272 12102 20300 12582
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 19616 11756 19668 11762
rect 19536 11716 19616 11744
rect 18696 11222 18748 11228
rect 19168 11206 19472 11234
rect 19168 11150 19196 11206
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19338 11112 19394 11121
rect 18524 10810 18552 11086
rect 19338 11047 19394 11056
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18340 10606 18368 10678
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18340 9654 18368 10542
rect 18708 10062 18736 10950
rect 19352 10674 19380 11047
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19260 10198 19288 10406
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16132 7410 16160 8298
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16224 8090 16252 8230
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16040 7002 16068 7278
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 16408 6934 16436 8230
rect 16820 8188 17128 8197
rect 16820 8186 16826 8188
rect 16882 8186 16906 8188
rect 16962 8186 16986 8188
rect 17042 8186 17066 8188
rect 17122 8186 17128 8188
rect 16882 8134 16884 8186
rect 17064 8134 17066 8186
rect 16820 8132 16826 8134
rect 16882 8132 16906 8134
rect 16962 8132 16986 8134
rect 17042 8132 17066 8134
rect 17122 8132 17128 8134
rect 16820 8123 17128 8132
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7478 16528 7686
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 16500 5642 16528 7414
rect 17328 7342 17356 7822
rect 17420 7750 17448 8774
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 16820 7100 17128 7109
rect 16820 7098 16826 7100
rect 16882 7098 16906 7100
rect 16962 7098 16986 7100
rect 17042 7098 17066 7100
rect 17122 7098 17128 7100
rect 16882 7046 16884 7098
rect 17064 7046 17066 7098
rect 16820 7044 16826 7046
rect 16882 7044 16906 7046
rect 16962 7044 16986 7046
rect 17042 7044 17066 7046
rect 17122 7044 17128 7046
rect 16820 7035 17128 7044
rect 17328 6798 17356 7278
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 16592 5778 16620 6734
rect 16820 6012 17128 6021
rect 16820 6010 16826 6012
rect 16882 6010 16906 6012
rect 16962 6010 16986 6012
rect 17042 6010 17066 6012
rect 17122 6010 17128 6012
rect 16882 5958 16884 6010
rect 17064 5958 17066 6010
rect 16820 5956 16826 5958
rect 16882 5956 16906 5958
rect 16962 5956 16986 5958
rect 17042 5956 17066 5958
rect 17122 5956 17128 5958
rect 16820 5947 17128 5956
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 17328 5710 17356 6734
rect 17420 6254 17448 7686
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17604 7002 17632 7142
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17696 6730 17724 7686
rect 17788 7274 17816 8366
rect 17880 7342 17908 8842
rect 18340 8294 18368 9590
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18432 9178 18460 9454
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18892 8974 18920 10134
rect 19444 10044 19472 11206
rect 19536 11014 19564 11716
rect 19616 11698 19668 11704
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19628 11218 19656 11494
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19536 10742 19564 10950
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19628 10606 19656 10950
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19720 10266 19748 11698
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19812 10742 19840 11018
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19812 10198 19840 10678
rect 19904 10674 19932 12038
rect 19994 11996 20302 12005
rect 19994 11994 20000 11996
rect 20056 11994 20080 11996
rect 20136 11994 20160 11996
rect 20216 11994 20240 11996
rect 20296 11994 20302 11996
rect 20056 11942 20058 11994
rect 20238 11942 20240 11994
rect 19994 11940 20000 11942
rect 20056 11940 20080 11942
rect 20136 11940 20160 11942
rect 20216 11940 20240 11942
rect 20296 11940 20302 11942
rect 19994 11931 20302 11940
rect 20364 11898 20392 16646
rect 20916 16590 20944 17138
rect 21008 16590 21036 17478
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20916 16250 20944 16390
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 21100 15706 21128 17478
rect 21638 17232 21694 17241
rect 21638 17167 21694 17176
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20916 15094 20944 15506
rect 21192 15502 21220 17070
rect 21652 16794 21680 17167
rect 22020 17134 22048 18158
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22112 17610 22140 17818
rect 22204 17746 22232 18226
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22284 17536 22336 17542
rect 22112 17484 22284 17490
rect 22112 17478 22336 17484
rect 22112 17462 22324 17478
rect 22112 17202 22140 17462
rect 22284 17332 22336 17338
rect 22388 17320 22416 17614
rect 22336 17292 22416 17320
rect 22284 17274 22336 17280
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 20904 15088 20956 15094
rect 20824 15036 20904 15042
rect 20824 15030 20956 15036
rect 20824 15014 20944 15030
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20640 13870 20668 14350
rect 20824 14006 20852 15014
rect 21100 14414 21128 15302
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 14482 21404 14758
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20456 13530 20484 13806
rect 20640 13530 20668 13806
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20916 13326 20944 14214
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13394 21404 13670
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20456 12850 20484 13194
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20904 12844 20956 12850
rect 21376 12832 21404 13330
rect 21456 12844 21508 12850
rect 21376 12804 21456 12832
rect 20904 12786 20956 12792
rect 21456 12786 21508 12792
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12434 20760 12582
rect 20456 12406 20760 12434
rect 20456 12374 20484 12406
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20824 12170 20852 12718
rect 20916 12442 20944 12786
rect 21560 12782 21588 16662
rect 21732 16652 21784 16658
rect 21916 16652 21968 16658
rect 21784 16612 21916 16640
rect 21732 16594 21784 16600
rect 21916 16594 21968 16600
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 22020 16046 22048 16526
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 22296 15094 22324 17138
rect 22480 17105 22508 17206
rect 22466 17096 22522 17105
rect 22466 17031 22522 17040
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16522 22416 16934
rect 22572 16658 22600 18022
rect 22756 17762 22784 18226
rect 22848 17882 22876 18702
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 23308 18358 23336 18566
rect 26342 18524 26650 18533
rect 26342 18522 26348 18524
rect 26404 18522 26428 18524
rect 26484 18522 26508 18524
rect 26564 18522 26588 18524
rect 26644 18522 26650 18524
rect 26404 18470 26406 18522
rect 26586 18470 26588 18522
rect 26342 18468 26348 18470
rect 26404 18468 26428 18470
rect 26484 18468 26508 18470
rect 26564 18468 26588 18470
rect 26644 18468 26650 18470
rect 26342 18459 26650 18468
rect 23296 18352 23348 18358
rect 23296 18294 23348 18300
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 23388 18216 23440 18222
rect 25136 18216 25188 18222
rect 23440 18164 23612 18170
rect 23388 18158 23612 18164
rect 25136 18158 25188 18164
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 22756 17734 22876 17762
rect 22848 17610 22876 17734
rect 22940 17678 22968 18158
rect 23400 18142 23612 18158
rect 23168 17980 23476 17989
rect 23168 17978 23174 17980
rect 23230 17978 23254 17980
rect 23310 17978 23334 17980
rect 23390 17978 23414 17980
rect 23470 17978 23476 17980
rect 23230 17926 23232 17978
rect 23412 17926 23414 17978
rect 23168 17924 23174 17926
rect 23230 17924 23254 17926
rect 23310 17924 23334 17926
rect 23390 17924 23414 17926
rect 23470 17924 23476 17926
rect 23168 17915 23476 17924
rect 23584 17814 23612 18142
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 23572 17808 23624 17814
rect 23308 17756 23572 17762
rect 23308 17750 23624 17756
rect 23308 17734 23612 17750
rect 24136 17746 24164 18022
rect 25148 17954 25176 18158
rect 25056 17926 25176 17954
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24124 17740 24176 17746
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22836 17604 22888 17610
rect 22836 17546 22888 17552
rect 22848 17338 22876 17546
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22650 17232 22706 17241
rect 22650 17167 22652 17176
rect 22704 17167 22706 17176
rect 22652 17138 22704 17144
rect 22744 17128 22796 17134
rect 22744 17070 22796 17076
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22664 16658 22692 17002
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 22388 16250 22416 16458
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22388 15162 22416 15438
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22664 15094 22692 16594
rect 22756 16522 22784 17070
rect 22848 16658 22876 17274
rect 22940 17134 22968 17614
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22940 16726 22968 16934
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 22928 16516 22980 16522
rect 22928 16458 22980 16464
rect 22940 15978 22968 16458
rect 23032 16436 23060 17478
rect 23308 17202 23336 17734
rect 24124 17682 24176 17688
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 23572 17128 23624 17134
rect 23676 17105 23704 17478
rect 23572 17070 23624 17076
rect 23662 17096 23718 17105
rect 23168 16892 23476 16901
rect 23168 16890 23174 16892
rect 23230 16890 23254 16892
rect 23310 16890 23334 16892
rect 23390 16890 23414 16892
rect 23470 16890 23476 16892
rect 23230 16838 23232 16890
rect 23412 16838 23414 16890
rect 23168 16836 23174 16838
rect 23230 16836 23254 16838
rect 23310 16836 23334 16838
rect 23390 16836 23414 16838
rect 23470 16836 23476 16838
rect 23168 16827 23476 16836
rect 23584 16794 23612 17070
rect 23662 17031 23718 17040
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 23572 16516 23624 16522
rect 23676 16504 23704 17031
rect 23624 16476 23704 16504
rect 23572 16458 23624 16464
rect 23112 16448 23164 16454
rect 23032 16408 23112 16436
rect 23032 16250 23060 16408
rect 23112 16390 23164 16396
rect 23400 16250 23428 16458
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23492 16182 23520 16458
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 22928 15972 22980 15978
rect 22928 15914 22980 15920
rect 23168 15804 23476 15813
rect 23168 15802 23174 15804
rect 23230 15802 23254 15804
rect 23310 15802 23334 15804
rect 23390 15802 23414 15804
rect 23470 15802 23476 15804
rect 23230 15750 23232 15802
rect 23412 15750 23414 15802
rect 23168 15748 23174 15750
rect 23230 15748 23254 15750
rect 23310 15748 23334 15750
rect 23390 15748 23414 15750
rect 23470 15748 23476 15750
rect 23168 15739 23476 15748
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22652 15088 22704 15094
rect 22652 15030 22704 15036
rect 22848 14618 22876 15098
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22204 13938 22232 14486
rect 23032 14482 23060 14894
rect 23124 14822 23152 15506
rect 23676 15162 23704 16476
rect 23768 16640 23796 17478
rect 23940 16652 23992 16658
rect 23768 16612 23940 16640
rect 23768 16182 23796 16612
rect 23940 16594 23992 16600
rect 24044 16522 24072 17478
rect 24136 17354 24164 17682
rect 24136 17338 24256 17354
rect 24136 17332 24268 17338
rect 24136 17326 24216 17332
rect 24216 17274 24268 17280
rect 24872 17202 24900 17818
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24032 16516 24084 16522
rect 24032 16458 24084 16464
rect 24044 16250 24072 16458
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23756 16176 23808 16182
rect 23756 16118 23808 16124
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23768 15076 23796 16118
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23848 15088 23900 15094
rect 23768 15048 23848 15076
rect 23664 14884 23716 14890
rect 23664 14826 23716 14832
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23168 14716 23476 14725
rect 23168 14714 23174 14716
rect 23230 14714 23254 14716
rect 23310 14714 23334 14716
rect 23390 14714 23414 14716
rect 23470 14714 23476 14716
rect 23230 14662 23232 14714
rect 23412 14662 23414 14714
rect 23168 14660 23174 14662
rect 23230 14660 23254 14662
rect 23310 14660 23334 14662
rect 23390 14660 23414 14662
rect 23470 14660 23476 14662
rect 23168 14651 23476 14660
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22664 13870 22692 14214
rect 23032 14006 23060 14418
rect 23584 14414 23612 14758
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23676 14006 23704 14826
rect 23768 14618 23796 15048
rect 23848 15030 23900 15036
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23860 14618 23888 14758
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23848 14612 23900 14618
rect 23848 14554 23900 14560
rect 23952 14074 23980 15438
rect 24044 14618 24072 16186
rect 24228 15434 24256 16934
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24596 15910 24624 16050
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24596 15570 24624 15846
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24136 14822 24164 14962
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24228 14414 24256 15370
rect 24492 15360 24544 15366
rect 24492 15302 24544 15308
rect 24504 15094 24532 15302
rect 24872 15094 24900 17138
rect 24964 16794 24992 17546
rect 25056 17542 25084 17926
rect 25044 17536 25096 17542
rect 26148 17536 26200 17542
rect 25096 17484 25176 17490
rect 25044 17478 25176 17484
rect 26148 17478 26200 17484
rect 25056 17462 25176 17478
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 25056 16658 25084 17274
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 25056 16266 25084 16594
rect 24964 16250 25084 16266
rect 24952 16244 25084 16250
rect 25004 16238 25084 16244
rect 24952 16186 25004 16192
rect 25056 16114 25084 16238
rect 25148 16182 25176 17462
rect 26160 17202 26188 17478
rect 26342 17436 26650 17445
rect 26342 17434 26348 17436
rect 26404 17434 26428 17436
rect 26484 17434 26508 17436
rect 26564 17434 26588 17436
rect 26644 17434 26650 17436
rect 26404 17382 26406 17434
rect 26586 17382 26588 17434
rect 26342 17380 26348 17382
rect 26404 17380 26428 17382
rect 26484 17380 26508 17382
rect 26564 17380 26588 17382
rect 26644 17380 26650 17382
rect 26342 17371 26650 17380
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25332 16096 25360 17138
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25504 16720 25556 16726
rect 25504 16662 25556 16668
rect 25516 16522 25544 16662
rect 25976 16658 26004 16934
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25424 16250 25452 16458
rect 25516 16250 25544 16458
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25596 16176 25648 16182
rect 25596 16118 25648 16124
rect 25412 16108 25464 16114
rect 25332 16068 25412 16096
rect 25332 15910 25360 16068
rect 25412 16050 25464 16056
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24964 15162 24992 15438
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24492 15088 24544 15094
rect 24492 15030 24544 15036
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 23664 14000 23716 14006
rect 23664 13942 23716 13948
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21744 12850 21772 13738
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20456 11626 20484 12038
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 19994 10908 20302 10917
rect 19994 10906 20000 10908
rect 20056 10906 20080 10908
rect 20136 10906 20160 10908
rect 20216 10906 20240 10908
rect 20296 10906 20302 10908
rect 20056 10854 20058 10906
rect 20238 10854 20240 10906
rect 19994 10852 20000 10854
rect 20056 10852 20080 10854
rect 20136 10852 20160 10854
rect 20216 10852 20240 10854
rect 20296 10852 20302 10854
rect 19994 10843 20302 10852
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19616 10056 19668 10062
rect 19444 10016 19616 10044
rect 19616 9998 19668 10004
rect 19628 9518 19656 9998
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7478 18736 7754
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 18708 6798 18736 7414
rect 18892 7206 18920 7822
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17420 5710 17448 6190
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 16500 5386 16528 5578
rect 16316 5358 16528 5386
rect 16960 5370 16988 5578
rect 16580 5364 16632 5370
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15672 4826 15792 4842
rect 15856 4826 15884 5170
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16132 4826 16160 4966
rect 15384 4820 15436 4826
rect 15672 4820 15804 4826
rect 15672 4814 15752 4820
rect 15384 4762 15436 4768
rect 15752 4762 15804 4768
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15198 4176 15254 4185
rect 15198 4111 15254 4120
rect 15304 4010 15332 4558
rect 15488 4554 15516 4694
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15672 4282 15700 4422
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 3194 15700 3878
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15016 3120 15068 3126
rect 15014 3088 15016 3097
rect 15108 3120 15160 3126
rect 15068 3088 15070 3097
rect 15108 3062 15160 3068
rect 15856 3058 15884 4422
rect 16040 4078 16068 4558
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16132 4078 16160 4490
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16120 4072 16172 4078
rect 16172 4020 16252 4026
rect 16120 4014 16252 4020
rect 15948 3738 15976 4014
rect 16132 3998 16252 4014
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16132 3058 16160 3878
rect 16224 3738 16252 3998
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16316 3466 16344 5358
rect 16580 5306 16632 5312
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16396 5296 16448 5302
rect 16448 5244 16528 5250
rect 16396 5238 16528 5244
rect 16408 5222 16528 5238
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16408 4622 16436 5102
rect 16500 4622 16528 5222
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16592 4282 16620 5306
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 16820 4924 17128 4933
rect 16820 4922 16826 4924
rect 16882 4922 16906 4924
rect 16962 4922 16986 4924
rect 17042 4922 17066 4924
rect 17122 4922 17128 4924
rect 16882 4870 16884 4922
rect 17064 4870 17066 4922
rect 16820 4868 16826 4870
rect 16882 4868 16906 4870
rect 16962 4868 16986 4870
rect 17042 4868 17066 4870
rect 17122 4868 17128 4870
rect 16820 4859 17128 4868
rect 17236 4826 17264 5170
rect 17328 5166 17356 5646
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16684 4146 16712 4490
rect 16776 4146 16804 4762
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3194 16436 3334
rect 16684 3194 16712 4082
rect 17144 4078 17172 4558
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17236 4010 17264 4490
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 16820 3836 17128 3845
rect 16820 3834 16826 3836
rect 16882 3834 16906 3836
rect 16962 3834 16986 3836
rect 17042 3834 17066 3836
rect 17122 3834 17128 3836
rect 16882 3782 16884 3834
rect 17064 3782 17066 3834
rect 16820 3780 16826 3782
rect 16882 3780 16906 3782
rect 16962 3780 16986 3782
rect 17042 3780 17066 3782
rect 17122 3780 17128 3782
rect 16820 3771 17128 3780
rect 17328 3602 17356 5102
rect 17420 4622 17448 5646
rect 17512 4622 17540 5646
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17604 4826 17632 5238
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17696 4706 17724 4966
rect 17604 4678 17724 4706
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17604 4486 17632 4678
rect 17880 4486 17908 5510
rect 18708 5234 18736 6734
rect 18892 6458 18920 7142
rect 19352 6798 19380 7686
rect 19536 7546 19564 7958
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19720 6866 19748 8366
rect 19812 7886 19840 10134
rect 19994 9820 20302 9829
rect 19994 9818 20000 9820
rect 20056 9818 20080 9820
rect 20136 9818 20160 9820
rect 20216 9818 20240 9820
rect 20296 9818 20302 9820
rect 20056 9766 20058 9818
rect 20238 9766 20240 9818
rect 19994 9764 20000 9766
rect 20056 9764 20080 9766
rect 20136 9764 20160 9766
rect 20216 9764 20240 9766
rect 20296 9764 20302 9766
rect 19994 9755 20302 9764
rect 19994 8732 20302 8741
rect 19994 8730 20000 8732
rect 20056 8730 20080 8732
rect 20136 8730 20160 8732
rect 20216 8730 20240 8732
rect 20296 8730 20302 8732
rect 20056 8678 20058 8730
rect 20238 8678 20240 8730
rect 19994 8676 20000 8678
rect 20056 8676 20080 8678
rect 20136 8676 20160 8678
rect 20216 8676 20240 8678
rect 20296 8676 20302 8678
rect 19994 8667 20302 8676
rect 20364 8634 20392 10610
rect 20916 10130 20944 12242
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21192 11762 21220 12038
rect 21560 11914 21588 12106
rect 21744 12102 21772 12786
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21928 12434 21956 12582
rect 21836 12406 21956 12434
rect 21836 12238 21864 12406
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21836 11914 21864 12174
rect 21560 11886 21864 11914
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21284 11218 21312 11494
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20456 8838 20484 9862
rect 21192 9722 21220 9930
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20548 9042 20576 9386
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20640 8634 20668 8910
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19904 7954 19932 8298
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19904 7546 19932 7890
rect 19994 7644 20302 7653
rect 19994 7642 20000 7644
rect 20056 7642 20080 7644
rect 20136 7642 20160 7644
rect 20216 7642 20240 7644
rect 20296 7642 20302 7644
rect 20056 7590 20058 7642
rect 20238 7590 20240 7642
rect 19994 7588 20000 7590
rect 20056 7588 20080 7590
rect 20136 7588 20160 7590
rect 20216 7588 20240 7590
rect 20296 7588 20302 7590
rect 19994 7579 20302 7588
rect 20364 7546 20392 8434
rect 20640 7954 20668 8570
rect 20732 8566 20760 8910
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 21284 8430 21312 9522
rect 21560 8906 21588 11886
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21652 10742 21680 11086
rect 22112 11082 22140 12786
rect 22664 12714 22692 13670
rect 23168 13628 23476 13637
rect 23168 13626 23174 13628
rect 23230 13626 23254 13628
rect 23310 13626 23334 13628
rect 23390 13626 23414 13628
rect 23470 13626 23476 13628
rect 23230 13574 23232 13626
rect 23412 13574 23414 13626
rect 23168 13572 23174 13574
rect 23230 13572 23254 13574
rect 23310 13572 23334 13574
rect 23390 13572 23414 13574
rect 23470 13572 23476 13574
rect 23168 13563 23476 13572
rect 23676 13530 23704 13942
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23860 13394 23888 13670
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 22652 12708 22704 12714
rect 22652 12650 22704 12656
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22756 11898 22784 12242
rect 23032 12170 23060 13126
rect 23860 12986 23888 13330
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 23572 12844 23624 12850
rect 23624 12804 23796 12832
rect 23572 12786 23624 12792
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23168 12540 23476 12549
rect 23168 12538 23174 12540
rect 23230 12538 23254 12540
rect 23310 12538 23334 12540
rect 23390 12538 23414 12540
rect 23470 12538 23476 12540
rect 23230 12486 23232 12538
rect 23412 12486 23414 12538
rect 23168 12484 23174 12486
rect 23230 12484 23254 12486
rect 23310 12484 23334 12486
rect 23390 12484 23414 12486
rect 23470 12484 23476 12486
rect 23168 12475 23476 12484
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22756 11354 22784 11834
rect 23492 11830 23520 12038
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23492 11642 23520 11766
rect 23676 11694 23704 12582
rect 23768 12170 23796 12804
rect 23860 12442 23888 12922
rect 23952 12918 23980 13874
rect 24044 13734 24072 14282
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24228 13258 24256 13466
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 24044 12782 24072 13194
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 24136 12170 24164 13126
rect 24320 12306 24348 14894
rect 24964 14346 24992 15098
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 24952 14340 25004 14346
rect 24952 14282 25004 14288
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24412 13326 24440 14214
rect 24780 14074 24808 14214
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 24872 13802 24900 13874
rect 24860 13796 24912 13802
rect 24860 13738 24912 13744
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24504 12782 24532 13466
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24596 12918 24624 13262
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 24688 12986 24716 13194
rect 24780 12986 24808 13194
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24872 12730 24900 13738
rect 24964 13326 24992 13874
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25056 13326 25084 13670
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25056 12850 25084 13262
rect 25148 13240 25176 14758
rect 25240 13870 25268 14894
rect 25424 14414 25452 15846
rect 25608 15026 25636 16118
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25700 14822 25728 16458
rect 25884 15978 25912 16526
rect 26342 16348 26650 16357
rect 26342 16346 26348 16348
rect 26404 16346 26428 16348
rect 26484 16346 26508 16348
rect 26564 16346 26588 16348
rect 26644 16346 26650 16348
rect 26404 16294 26406 16346
rect 26586 16294 26588 16346
rect 26342 16292 26348 16294
rect 26404 16292 26428 16294
rect 26484 16292 26508 16294
rect 26564 16292 26588 16294
rect 26644 16292 26650 16294
rect 26342 16283 26650 16292
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 25792 15570 25820 15846
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26068 15162 26096 15438
rect 26342 15260 26650 15269
rect 26342 15258 26348 15260
rect 26404 15258 26428 15260
rect 26484 15258 26508 15260
rect 26564 15258 26588 15260
rect 26644 15258 26650 15260
rect 26404 15206 26406 15258
rect 26586 15206 26588 15258
rect 26342 15204 26348 15206
rect 26404 15204 26428 15206
rect 26484 15204 26508 15206
rect 26564 15204 26588 15206
rect 26644 15204 26650 15206
rect 26342 15195 26650 15204
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 25516 14006 25544 14214
rect 26342 14172 26650 14181
rect 26342 14170 26348 14172
rect 26404 14170 26428 14172
rect 26484 14170 26508 14172
rect 26564 14170 26588 14172
rect 26644 14170 26650 14172
rect 26404 14118 26406 14170
rect 26586 14118 26588 14170
rect 26342 14116 26348 14118
rect 26404 14116 26428 14118
rect 26484 14116 26508 14118
rect 26564 14116 26588 14118
rect 26644 14116 26650 14118
rect 26342 14107 26650 14116
rect 25504 14000 25556 14006
rect 25504 13942 25556 13948
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25516 13258 25544 13942
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 25228 13252 25280 13258
rect 25148 13212 25228 13240
rect 25228 13194 25280 13200
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25148 12730 25176 12786
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 24124 12164 24176 12170
rect 24124 12106 24176 12112
rect 23664 11688 23716 11694
rect 23492 11614 23612 11642
rect 23664 11630 23716 11636
rect 23168 11452 23476 11461
rect 23168 11450 23174 11452
rect 23230 11450 23254 11452
rect 23310 11450 23334 11452
rect 23390 11450 23414 11452
rect 23470 11450 23476 11452
rect 23230 11398 23232 11450
rect 23412 11398 23414 11450
rect 23168 11396 23174 11398
rect 23230 11396 23254 11398
rect 23310 11396 23334 11398
rect 23390 11396 23414 11398
rect 23470 11396 23476 11398
rect 23168 11387 23476 11396
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 21640 10736 21692 10742
rect 21640 10678 21692 10684
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 22020 9178 22048 9522
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7546 20576 7686
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19352 6458 19380 6734
rect 19800 6724 19852 6730
rect 19800 6666 19852 6672
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19444 6186 19472 6598
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19628 5778 19656 6394
rect 19812 6390 19840 6666
rect 19994 6556 20302 6565
rect 19994 6554 20000 6556
rect 20056 6554 20080 6556
rect 20136 6554 20160 6556
rect 20216 6554 20240 6556
rect 20296 6554 20302 6556
rect 20056 6502 20058 6554
rect 20238 6502 20240 6554
rect 19994 6500 20000 6502
rect 20056 6500 20080 6502
rect 20136 6500 20160 6502
rect 20216 6500 20240 6502
rect 20296 6500 20302 6502
rect 19994 6491 20302 6500
rect 20640 6458 20668 7890
rect 20824 7818 20852 8298
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20732 7528 20760 7686
rect 20812 7540 20864 7546
rect 20732 7500 20812 7528
rect 20812 7482 20864 7488
rect 20824 7274 20852 7482
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 19904 5370 19932 5578
rect 19994 5468 20302 5477
rect 19994 5466 20000 5468
rect 20056 5466 20080 5468
rect 20136 5466 20160 5468
rect 20216 5466 20240 5468
rect 20296 5466 20302 5468
rect 20056 5414 20058 5466
rect 20238 5414 20240 5466
rect 19994 5412 20000 5414
rect 20056 5412 20080 5414
rect 20136 5412 20160 5414
rect 20216 5412 20240 5414
rect 20296 5412 20302 5414
rect 19994 5403 20302 5412
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18156 4622 18184 5102
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17604 4146 17632 4422
rect 17880 4146 17908 4422
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17038 3360 17094 3369
rect 17038 3295 17094 3304
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 17052 3058 17080 3295
rect 17144 3058 17172 3470
rect 17420 3398 17448 4082
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17788 3738 17816 3878
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17592 3460 17644 3466
rect 17592 3402 17644 3408
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 15014 3023 15070 3032
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17420 2990 17448 3334
rect 17604 3194 17632 3402
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17788 2922 17816 3674
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 16040 2514 16068 2790
rect 17972 2774 18000 3878
rect 16820 2748 17128 2757
rect 16820 2746 16826 2748
rect 16882 2746 16906 2748
rect 16962 2746 16986 2748
rect 17042 2746 17066 2748
rect 17122 2746 17128 2748
rect 17972 2746 18092 2774
rect 16882 2694 16884 2746
rect 17064 2694 17066 2746
rect 16820 2692 16826 2694
rect 16882 2692 16906 2694
rect 16962 2692 16986 2694
rect 17042 2692 17066 2694
rect 17122 2692 17128 2694
rect 16820 2683 17128 2692
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 14924 2508 14976 2514
rect 14924 2450 14976 2456
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 18064 2446 18092 2746
rect 18156 2446 18184 4082
rect 18248 2446 18276 4966
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18432 4010 18460 4558
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 18524 3942 18552 4490
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18616 4010 18644 4218
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18708 3534 18736 5170
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19260 4706 19288 4966
rect 19260 4678 19472 4706
rect 20640 4690 20668 6394
rect 21192 6322 21220 7754
rect 21284 7546 21312 8366
rect 22204 7750 22232 9930
rect 22572 9518 22600 10542
rect 23168 10364 23476 10373
rect 23168 10362 23174 10364
rect 23230 10362 23254 10364
rect 23310 10362 23334 10364
rect 23390 10362 23414 10364
rect 23470 10362 23476 10364
rect 23230 10310 23232 10362
rect 23412 10310 23414 10362
rect 23168 10308 23174 10310
rect 23230 10308 23254 10310
rect 23310 10308 23334 10310
rect 23390 10308 23414 10310
rect 23470 10308 23476 10310
rect 23168 10299 23476 10308
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22756 9722 22784 10202
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23584 10010 23612 11614
rect 23768 10130 23796 12106
rect 24504 11898 24532 12718
rect 24872 12702 25176 12730
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 25976 11626 26004 13126
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 26068 12442 26096 12786
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 26160 12345 26188 13262
rect 26342 13084 26650 13093
rect 26342 13082 26348 13084
rect 26404 13082 26428 13084
rect 26484 13082 26508 13084
rect 26564 13082 26588 13084
rect 26644 13082 26650 13084
rect 26404 13030 26406 13082
rect 26586 13030 26588 13082
rect 26342 13028 26348 13030
rect 26404 13028 26428 13030
rect 26484 13028 26508 13030
rect 26564 13028 26588 13030
rect 26644 13028 26650 13030
rect 26342 13019 26650 13028
rect 26146 12336 26202 12345
rect 26146 12271 26202 12280
rect 26342 11996 26650 12005
rect 26342 11994 26348 11996
rect 26404 11994 26428 11996
rect 26484 11994 26508 11996
rect 26564 11994 26588 11996
rect 26644 11994 26650 11996
rect 26404 11942 26406 11994
rect 26586 11942 26588 11994
rect 26342 11940 26348 11942
rect 26404 11940 26428 11942
rect 26484 11940 26508 11942
rect 26564 11940 26588 11942
rect 26644 11940 26650 11942
rect 26342 11931 26650 11940
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 26342 10908 26650 10917
rect 26342 10906 26348 10908
rect 26404 10906 26428 10908
rect 26484 10906 26508 10908
rect 26564 10906 26588 10908
rect 26644 10906 26650 10908
rect 26404 10854 26406 10906
rect 26586 10854 26588 10906
rect 26342 10852 26348 10854
rect 26404 10852 26428 10854
rect 26484 10852 26508 10854
rect 26564 10852 26588 10854
rect 26644 10852 26650 10854
rect 26342 10843 26650 10852
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 24584 10056 24636 10062
rect 22836 9988 22888 9994
rect 22836 9930 22888 9936
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22848 9518 22876 9930
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 23032 9722 23060 9862
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22836 9512 22888 9518
rect 23124 9466 23152 9998
rect 23584 9982 24072 10010
rect 24584 9998 24636 10004
rect 25504 10056 25556 10062
rect 25504 9998 25556 10004
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 22836 9454 22888 9460
rect 22572 8634 22600 9454
rect 22848 8974 22876 9454
rect 23032 9438 23152 9466
rect 23492 9466 23520 9862
rect 23584 9654 23612 9982
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23492 9438 23612 9466
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22388 7750 22416 8366
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21192 5642 21220 6258
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 21560 5370 21588 7142
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21744 6458 21772 6598
rect 21836 6458 21864 7346
rect 22388 7342 22416 7686
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 21732 6248 21784 6254
rect 21652 6196 21732 6202
rect 21652 6190 21784 6196
rect 21652 6174 21772 6190
rect 21652 5846 21680 6174
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21744 5914 21772 6054
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21640 5840 21692 5846
rect 21640 5782 21692 5788
rect 21916 5568 21968 5574
rect 21916 5510 21968 5516
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18984 4486 19012 4558
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18708 3126 18736 3470
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18340 2650 18368 2926
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 7298 2204 7606 2213
rect 7298 2202 7304 2204
rect 7360 2202 7384 2204
rect 7440 2202 7464 2204
rect 7520 2202 7544 2204
rect 7600 2202 7606 2204
rect 7360 2150 7362 2202
rect 7542 2150 7544 2202
rect 7298 2148 7304 2150
rect 7360 2148 7384 2150
rect 7440 2148 7464 2150
rect 7520 2148 7544 2150
rect 7600 2148 7606 2150
rect 7298 2139 7606 2148
rect 10428 1306 10456 2382
rect 18524 2378 18552 2790
rect 18800 2514 18828 3878
rect 18892 3602 18920 4422
rect 18984 4078 19012 4422
rect 19260 4282 19288 4678
rect 19444 4622 19472 4678
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19352 4078 19380 4558
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19628 4146 19656 4422
rect 19812 4282 19840 4558
rect 19994 4380 20302 4389
rect 19994 4378 20000 4380
rect 20056 4378 20080 4380
rect 20136 4378 20160 4380
rect 20216 4378 20240 4380
rect 20296 4378 20302 4380
rect 20056 4326 20058 4378
rect 20238 4326 20240 4378
rect 19994 4324 20000 4326
rect 20056 4324 20080 4326
rect 20136 4324 20160 4326
rect 20216 4324 20240 4326
rect 20296 4324 20302 4326
rect 19994 4315 20302 4324
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 19168 2446 19196 3470
rect 19352 3398 19380 4014
rect 19996 3738 20024 4082
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20088 3738 20116 3878
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19994 3292 20302 3301
rect 19994 3290 20000 3292
rect 20056 3290 20080 3292
rect 20136 3290 20160 3292
rect 20216 3290 20240 3292
rect 20296 3290 20302 3292
rect 20056 3238 20058 3290
rect 20238 3238 20240 3290
rect 19994 3236 20000 3238
rect 20056 3236 20080 3238
rect 20136 3236 20160 3238
rect 20216 3236 20240 3238
rect 20296 3236 20302 3238
rect 19994 3227 20302 3236
rect 20364 3194 20392 3878
rect 20640 3602 20668 4626
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20640 3058 20668 3538
rect 20916 3194 20944 4490
rect 21284 3602 21312 4966
rect 21928 4554 21956 5510
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 22020 4826 22048 5170
rect 22204 5166 22232 6258
rect 22296 5234 22324 7210
rect 22480 5302 22508 7686
rect 22572 6458 22600 7890
rect 22848 7868 22876 8910
rect 22940 8362 22968 9318
rect 23032 9178 23060 9438
rect 23168 9276 23476 9285
rect 23168 9274 23174 9276
rect 23230 9274 23254 9276
rect 23310 9274 23334 9276
rect 23390 9274 23414 9276
rect 23470 9274 23476 9276
rect 23230 9222 23232 9274
rect 23412 9222 23414 9274
rect 23168 9220 23174 9222
rect 23230 9220 23254 9222
rect 23310 9220 23334 9222
rect 23390 9220 23414 9222
rect 23470 9220 23476 9222
rect 23168 9211 23476 9220
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23216 8498 23244 8774
rect 23492 8566 23520 8978
rect 23584 8974 23612 9438
rect 23676 8974 23704 9862
rect 23940 9036 23992 9042
rect 23940 8978 23992 8984
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23480 8560 23532 8566
rect 23584 8537 23612 8774
rect 23480 8502 23532 8508
rect 23570 8528 23626 8537
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 23204 8492 23256 8498
rect 23570 8463 23626 8472
rect 23204 8434 23256 8440
rect 22928 8356 22980 8362
rect 22928 8298 22980 8304
rect 23032 8090 23060 8434
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 23168 8188 23476 8197
rect 23168 8186 23174 8188
rect 23230 8186 23254 8188
rect 23310 8186 23334 8188
rect 23390 8186 23414 8188
rect 23470 8186 23476 8188
rect 23230 8134 23232 8186
rect 23412 8134 23414 8186
rect 23168 8132 23174 8134
rect 23230 8132 23254 8134
rect 23310 8132 23334 8134
rect 23390 8132 23414 8134
rect 23470 8132 23476 8134
rect 23168 8123 23476 8132
rect 23584 8090 23612 8366
rect 23676 8294 23704 8910
rect 23768 8634 23796 8910
rect 23848 8900 23900 8906
rect 23848 8842 23900 8848
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23768 8430 23796 8570
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23020 7880 23072 7886
rect 22848 7840 23020 7868
rect 23020 7822 23072 7828
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23032 7410 23060 7822
rect 23400 7546 23428 7822
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 22652 7404 22704 7410
rect 23020 7404 23072 7410
rect 22652 7346 22704 7352
rect 22940 7364 23020 7392
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22468 5296 22520 5302
rect 22572 5284 22600 6054
rect 22664 5574 22692 7346
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22848 6458 22876 6598
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 22848 5914 22876 6258
rect 22940 6254 22968 7364
rect 23020 7346 23072 7352
rect 23168 7100 23476 7109
rect 23168 7098 23174 7100
rect 23230 7098 23254 7100
rect 23310 7098 23334 7100
rect 23390 7098 23414 7100
rect 23470 7098 23476 7100
rect 23230 7046 23232 7098
rect 23412 7046 23414 7098
rect 23168 7044 23174 7046
rect 23230 7044 23254 7046
rect 23310 7044 23334 7046
rect 23390 7044 23414 7046
rect 23470 7044 23476 7046
rect 23168 7035 23476 7044
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 22928 6248 22980 6254
rect 22928 6190 22980 6196
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 22940 5914 22968 6054
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 22756 5370 22784 5850
rect 23032 5710 23060 6122
rect 23492 6118 23520 6734
rect 23584 6322 23612 6938
rect 23768 6798 23796 8366
rect 23860 7750 23888 8842
rect 23952 7886 23980 8978
rect 24044 8906 24072 9982
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 24308 9376 24360 9382
rect 24308 9318 24360 9324
rect 24320 9042 24348 9318
rect 24308 9036 24360 9042
rect 24308 8978 24360 8984
rect 24032 8900 24084 8906
rect 24032 8842 24084 8848
rect 24308 8832 24360 8838
rect 24308 8774 24360 8780
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 7410 23888 7686
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23952 7002 23980 7822
rect 24044 7818 24072 8570
rect 24032 7812 24084 7818
rect 24032 7754 24084 7760
rect 24044 7002 24072 7754
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24228 7546 24256 7686
rect 24320 7546 24348 8774
rect 24412 8566 24440 9862
rect 24400 8560 24452 8566
rect 24400 8502 24452 8508
rect 24596 8430 24624 9998
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24872 9722 24900 9930
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25056 9722 25084 9862
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 24872 9178 24900 9522
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24676 8900 24728 8906
rect 24676 8842 24728 8848
rect 24688 8566 24716 8842
rect 24964 8838 24992 9318
rect 25332 9042 25360 9862
rect 25516 9722 25544 9998
rect 26342 9820 26650 9829
rect 26342 9818 26348 9820
rect 26404 9818 26428 9820
rect 26484 9818 26508 9820
rect 26564 9818 26588 9820
rect 26644 9818 26650 9820
rect 26404 9766 26406 9818
rect 26586 9766 26588 9818
rect 26342 9764 26348 9766
rect 26404 9764 26428 9766
rect 26484 9764 26508 9766
rect 26564 9764 26588 9766
rect 26644 9764 26650 9766
rect 26342 9755 26650 9764
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 25872 9512 25924 9518
rect 25872 9454 25924 9460
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24858 8528 24914 8537
rect 24858 8463 24914 8472
rect 24872 8430 24900 8463
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 23952 6882 23980 6938
rect 23860 6854 23980 6882
rect 23860 6798 23888 6854
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23848 6792 23900 6798
rect 23848 6734 23900 6740
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23480 6112 23532 6118
rect 23532 6072 23612 6100
rect 23480 6054 23532 6060
rect 23168 6012 23476 6021
rect 23168 6010 23174 6012
rect 23230 6010 23254 6012
rect 23310 6010 23334 6012
rect 23390 6010 23414 6012
rect 23470 6010 23476 6012
rect 23230 5958 23232 6010
rect 23412 5958 23414 6010
rect 23168 5956 23174 5958
rect 23230 5956 23254 5958
rect 23310 5956 23334 5958
rect 23390 5956 23414 5958
rect 23470 5956 23476 5958
rect 23168 5947 23476 5956
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 22836 5636 22888 5642
rect 22836 5578 22888 5584
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22652 5296 22704 5302
rect 22572 5256 22652 5284
rect 22468 5238 22520 5244
rect 22652 5238 22704 5244
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22744 5228 22796 5234
rect 22848 5216 22876 5578
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23216 5370 23244 5510
rect 23584 5370 23612 6072
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 22928 5228 22980 5234
rect 22848 5188 22928 5216
rect 22744 5170 22796 5176
rect 22928 5170 22980 5176
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 21916 4548 21968 4554
rect 21916 4490 21968 4496
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 21836 3194 21864 3878
rect 21928 3602 21956 4490
rect 22296 4486 22324 5170
rect 22756 4622 22784 5170
rect 22940 4622 22968 5170
rect 23168 4924 23476 4933
rect 23168 4922 23174 4924
rect 23230 4922 23254 4924
rect 23310 4922 23334 4924
rect 23390 4922 23414 4924
rect 23470 4922 23476 4924
rect 23230 4870 23232 4922
rect 23412 4870 23414 4922
rect 23168 4868 23174 4870
rect 23230 4868 23254 4870
rect 23310 4868 23334 4870
rect 23390 4868 23414 4870
rect 23470 4868 23476 4870
rect 23168 4859 23476 4868
rect 23584 4758 23612 5306
rect 23676 5234 23704 6598
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 23572 4752 23624 4758
rect 23572 4694 23624 4700
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22296 4282 22324 4422
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 22664 3194 22692 3878
rect 22756 3738 22784 4558
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 22940 4060 22968 4422
rect 23032 4214 23060 4422
rect 23308 4214 23336 4422
rect 23584 4214 23612 4694
rect 23676 4554 23704 5170
rect 23664 4548 23716 4554
rect 23664 4490 23716 4496
rect 23020 4208 23072 4214
rect 23020 4150 23072 4156
rect 23296 4208 23348 4214
rect 23572 4208 23624 4214
rect 23296 4150 23348 4156
rect 23400 4156 23572 4162
rect 23400 4150 23624 4156
rect 23400 4146 23612 4150
rect 23676 4146 23704 4490
rect 23768 4146 23796 6734
rect 23860 6458 23888 6734
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 24320 6390 24348 6734
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24412 6322 24440 7142
rect 24504 6322 24532 7346
rect 24596 6390 24624 7482
rect 24964 7206 24992 8774
rect 25884 8634 25912 9454
rect 26342 8732 26650 8741
rect 26342 8730 26348 8732
rect 26404 8730 26428 8732
rect 26484 8730 26508 8732
rect 26564 8730 26588 8732
rect 26644 8730 26650 8732
rect 26404 8678 26406 8730
rect 26586 8678 26588 8730
rect 26342 8676 26348 8678
rect 26404 8676 26428 8678
rect 26484 8676 26508 8678
rect 26564 8676 26588 8678
rect 26644 8676 26650 8678
rect 26342 8667 26650 8676
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 25780 8356 25832 8362
rect 25780 8298 25832 8304
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 24952 7200 25004 7206
rect 24952 7142 25004 7148
rect 24872 6882 24900 7142
rect 24780 6866 24900 6882
rect 24768 6860 24900 6866
rect 24820 6854 24900 6860
rect 24768 6802 24820 6808
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24688 6458 24716 6666
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24584 6384 24636 6390
rect 24584 6326 24636 6332
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24216 5296 24268 5302
rect 24216 5238 24268 5244
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 23940 5024 23992 5030
rect 23940 4966 23992 4972
rect 23860 4282 23888 4966
rect 23952 4622 23980 4966
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 24228 4554 24256 5238
rect 24504 4622 24532 6258
rect 24964 5778 24992 7142
rect 25056 7002 25084 7346
rect 25044 6996 25096 7002
rect 25044 6938 25096 6944
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 25056 5710 25084 6938
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 25148 5370 25176 6190
rect 25240 5914 25268 7346
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25240 5302 25268 5850
rect 25412 5364 25464 5370
rect 25412 5306 25464 5312
rect 25228 5296 25280 5302
rect 25228 5238 25280 5244
rect 25240 4690 25268 5238
rect 25228 4684 25280 4690
rect 25228 4626 25280 4632
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 24216 4548 24268 4554
rect 24216 4490 24268 4496
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 24860 4480 24912 4486
rect 24860 4422 24912 4428
rect 23848 4276 23900 4282
rect 23848 4218 23900 4224
rect 23388 4140 23612 4146
rect 23440 4134 23612 4140
rect 23664 4140 23716 4146
rect 23388 4082 23440 4088
rect 23664 4082 23716 4088
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23020 4072 23072 4078
rect 22940 4032 23020 4060
rect 23020 4014 23072 4020
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 23032 3534 23060 4014
rect 23168 3836 23476 3845
rect 23168 3834 23174 3836
rect 23230 3834 23254 3836
rect 23310 3834 23334 3836
rect 23390 3834 23414 3836
rect 23470 3834 23476 3836
rect 23230 3782 23232 3834
rect 23412 3782 23414 3834
rect 23168 3780 23174 3782
rect 23230 3780 23254 3782
rect 23310 3780 23334 3782
rect 23390 3780 23414 3782
rect 23470 3780 23476 3782
rect 23168 3771 23476 3780
rect 23584 3738 23612 4014
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23860 3534 23888 4218
rect 24308 4208 24360 4214
rect 24308 4150 24360 4156
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 24044 3738 24072 4014
rect 24320 3738 24348 4150
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23768 3194 23796 3334
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 24320 3126 24348 3674
rect 24596 3602 24624 4422
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 24872 3534 24900 4422
rect 25240 4298 25268 4626
rect 25240 4282 25360 4298
rect 25240 4276 25372 4282
rect 25240 4270 25320 4276
rect 25320 4218 25372 4224
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 24860 3528 24912 3534
rect 25240 3516 25268 3878
rect 25332 3738 25360 4218
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25424 3534 25452 5306
rect 25700 4214 25728 6666
rect 25688 4208 25740 4214
rect 25688 4150 25740 4156
rect 25320 3528 25372 3534
rect 25240 3488 25320 3516
rect 24860 3470 24912 3476
rect 25320 3470 25372 3476
rect 25412 3528 25464 3534
rect 25412 3470 25464 3476
rect 25700 3194 25728 4150
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 23168 2748 23476 2757
rect 23168 2746 23174 2748
rect 23230 2746 23254 2748
rect 23310 2746 23334 2748
rect 23390 2746 23414 2748
rect 23470 2746 23476 2748
rect 23230 2694 23232 2746
rect 23412 2694 23414 2746
rect 23168 2692 23174 2694
rect 23230 2692 23254 2694
rect 23310 2692 23334 2694
rect 23390 2692 23414 2694
rect 23470 2692 23476 2694
rect 23168 2683 23476 2692
rect 25792 2446 25820 8298
rect 26342 7644 26650 7653
rect 26342 7642 26348 7644
rect 26404 7642 26428 7644
rect 26484 7642 26508 7644
rect 26564 7642 26588 7644
rect 26644 7642 26650 7644
rect 26404 7590 26406 7642
rect 26586 7590 26588 7642
rect 26342 7588 26348 7590
rect 26404 7588 26428 7590
rect 26484 7588 26508 7590
rect 26564 7588 26588 7590
rect 26644 7588 26650 7590
rect 26342 7579 26650 7588
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 26068 6322 26096 6938
rect 26342 6556 26650 6565
rect 26342 6554 26348 6556
rect 26404 6554 26428 6556
rect 26484 6554 26508 6556
rect 26564 6554 26588 6556
rect 26644 6554 26650 6556
rect 26404 6502 26406 6554
rect 26586 6502 26588 6554
rect 26342 6500 26348 6502
rect 26404 6500 26428 6502
rect 26484 6500 26508 6502
rect 26564 6500 26588 6502
rect 26644 6500 26650 6502
rect 26342 6491 26650 6500
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 26342 5468 26650 5477
rect 26342 5466 26348 5468
rect 26404 5466 26428 5468
rect 26484 5466 26508 5468
rect 26564 5466 26588 5468
rect 26644 5466 26650 5468
rect 26404 5414 26406 5466
rect 26586 5414 26588 5466
rect 26342 5412 26348 5414
rect 26404 5412 26428 5414
rect 26484 5412 26508 5414
rect 26564 5412 26588 5414
rect 26644 5412 26650 5414
rect 26342 5403 26650 5412
rect 26516 5024 26568 5030
rect 26516 4966 26568 4972
rect 26528 4865 26556 4966
rect 26514 4856 26570 4865
rect 26514 4791 26570 4800
rect 26342 4380 26650 4389
rect 26342 4378 26348 4380
rect 26404 4378 26428 4380
rect 26484 4378 26508 4380
rect 26564 4378 26588 4380
rect 26644 4378 26650 4380
rect 26404 4326 26406 4378
rect 26586 4326 26588 4378
rect 26342 4324 26348 4326
rect 26404 4324 26428 4326
rect 26484 4324 26508 4326
rect 26564 4324 26588 4326
rect 26644 4324 26650 4326
rect 26342 4315 26650 4324
rect 26342 3292 26650 3301
rect 26342 3290 26348 3292
rect 26404 3290 26428 3292
rect 26484 3290 26508 3292
rect 26564 3290 26588 3292
rect 26644 3290 26650 3292
rect 26404 3238 26406 3290
rect 26586 3238 26588 3290
rect 26342 3236 26348 3238
rect 26404 3236 26428 3238
rect 26484 3236 26508 3238
rect 26564 3236 26588 3238
rect 26644 3236 26650 3238
rect 26342 3227 26650 3236
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 13646 2204 13954 2213
rect 13646 2202 13652 2204
rect 13708 2202 13732 2204
rect 13788 2202 13812 2204
rect 13868 2202 13892 2204
rect 13948 2202 13954 2204
rect 13708 2150 13710 2202
rect 13890 2150 13892 2202
rect 13646 2148 13652 2150
rect 13708 2148 13732 2150
rect 13788 2148 13812 2150
rect 13868 2148 13892 2150
rect 13948 2148 13954 2150
rect 13646 2139 13954 2148
rect 10336 1278 10456 1306
rect 10336 800 10364 1278
rect 18064 800 18092 2246
rect 19994 2204 20302 2213
rect 19994 2202 20000 2204
rect 20056 2202 20080 2204
rect 20136 2202 20160 2204
rect 20216 2202 20240 2204
rect 20296 2202 20302 2204
rect 20056 2150 20058 2202
rect 20238 2150 20240 2202
rect 19994 2148 20000 2150
rect 20056 2148 20080 2150
rect 20136 2148 20160 2150
rect 20216 2148 20240 2150
rect 20296 2148 20302 2150
rect 19994 2139 20302 2148
rect 18 0 74 800
rect 3238 0 3294 800
rect 7102 0 7158 800
rect 10322 0 10378 800
rect 14186 0 14242 800
rect 18050 0 18106 800
rect 21270 0 21326 800
rect 25134 0 25190 800
rect 26160 785 26188 2314
rect 26342 2204 26650 2213
rect 26342 2202 26348 2204
rect 26404 2202 26428 2204
rect 26484 2202 26508 2204
rect 26564 2202 26588 2204
rect 26644 2202 26650 2204
rect 26404 2150 26406 2202
rect 26586 2150 26588 2202
rect 26342 2148 26348 2150
rect 26404 2148 26428 2150
rect 26484 2148 26508 2150
rect 26564 2148 26588 2150
rect 26644 2148 26650 2150
rect 26342 2139 26650 2148
rect 26146 776 26202 785
rect 26146 711 26202 720
<< via2 >>
rect 7304 27226 7360 27228
rect 7384 27226 7440 27228
rect 7464 27226 7520 27228
rect 7544 27226 7600 27228
rect 7304 27174 7350 27226
rect 7350 27174 7360 27226
rect 7384 27174 7414 27226
rect 7414 27174 7426 27226
rect 7426 27174 7440 27226
rect 7464 27174 7478 27226
rect 7478 27174 7490 27226
rect 7490 27174 7520 27226
rect 7544 27174 7554 27226
rect 7554 27174 7600 27226
rect 7304 27172 7360 27174
rect 7384 27172 7440 27174
rect 7464 27172 7520 27174
rect 7544 27172 7600 27174
rect 13652 27226 13708 27228
rect 13732 27226 13788 27228
rect 13812 27226 13868 27228
rect 13892 27226 13948 27228
rect 13652 27174 13698 27226
rect 13698 27174 13708 27226
rect 13732 27174 13762 27226
rect 13762 27174 13774 27226
rect 13774 27174 13788 27226
rect 13812 27174 13826 27226
rect 13826 27174 13838 27226
rect 13838 27174 13868 27226
rect 13892 27174 13902 27226
rect 13902 27174 13948 27226
rect 13652 27172 13708 27174
rect 13732 27172 13788 27174
rect 13812 27172 13868 27174
rect 13892 27172 13948 27174
rect 20000 27226 20056 27228
rect 20080 27226 20136 27228
rect 20160 27226 20216 27228
rect 20240 27226 20296 27228
rect 20000 27174 20046 27226
rect 20046 27174 20056 27226
rect 20080 27174 20110 27226
rect 20110 27174 20122 27226
rect 20122 27174 20136 27226
rect 20160 27174 20174 27226
rect 20174 27174 20186 27226
rect 20186 27174 20216 27226
rect 20240 27174 20250 27226
rect 20250 27174 20296 27226
rect 20000 27172 20056 27174
rect 20080 27172 20136 27174
rect 20160 27172 20216 27174
rect 20240 27172 20296 27174
rect 26348 27226 26404 27228
rect 26428 27226 26484 27228
rect 26508 27226 26564 27228
rect 26588 27226 26644 27228
rect 26348 27174 26394 27226
rect 26394 27174 26404 27226
rect 26428 27174 26458 27226
rect 26458 27174 26470 27226
rect 26470 27174 26484 27226
rect 26508 27174 26522 27226
rect 26522 27174 26534 27226
rect 26534 27174 26564 27226
rect 26588 27174 26598 27226
rect 26598 27174 26644 27226
rect 26348 27172 26404 27174
rect 26428 27172 26484 27174
rect 26508 27172 26564 27174
rect 26588 27172 26644 27174
rect 4130 26682 4186 26684
rect 4210 26682 4266 26684
rect 4290 26682 4346 26684
rect 4370 26682 4426 26684
rect 4130 26630 4176 26682
rect 4176 26630 4186 26682
rect 4210 26630 4240 26682
rect 4240 26630 4252 26682
rect 4252 26630 4266 26682
rect 4290 26630 4304 26682
rect 4304 26630 4316 26682
rect 4316 26630 4346 26682
rect 4370 26630 4380 26682
rect 4380 26630 4426 26682
rect 4130 26628 4186 26630
rect 4210 26628 4266 26630
rect 4290 26628 4346 26630
rect 4370 26628 4426 26630
rect 10478 26682 10534 26684
rect 10558 26682 10614 26684
rect 10638 26682 10694 26684
rect 10718 26682 10774 26684
rect 10478 26630 10524 26682
rect 10524 26630 10534 26682
rect 10558 26630 10588 26682
rect 10588 26630 10600 26682
rect 10600 26630 10614 26682
rect 10638 26630 10652 26682
rect 10652 26630 10664 26682
rect 10664 26630 10694 26682
rect 10718 26630 10728 26682
rect 10728 26630 10774 26682
rect 10478 26628 10534 26630
rect 10558 26628 10614 26630
rect 10638 26628 10694 26630
rect 10718 26628 10774 26630
rect 938 26560 994 26616
rect 7304 26138 7360 26140
rect 7384 26138 7440 26140
rect 7464 26138 7520 26140
rect 7544 26138 7600 26140
rect 7304 26086 7350 26138
rect 7350 26086 7360 26138
rect 7384 26086 7414 26138
rect 7414 26086 7426 26138
rect 7426 26086 7440 26138
rect 7464 26086 7478 26138
rect 7478 26086 7490 26138
rect 7490 26086 7520 26138
rect 7544 26086 7554 26138
rect 7554 26086 7600 26138
rect 7304 26084 7360 26086
rect 7384 26084 7440 26086
rect 7464 26084 7520 26086
rect 7544 26084 7600 26086
rect 4130 25594 4186 25596
rect 4210 25594 4266 25596
rect 4290 25594 4346 25596
rect 4370 25594 4426 25596
rect 4130 25542 4176 25594
rect 4176 25542 4186 25594
rect 4210 25542 4240 25594
rect 4240 25542 4252 25594
rect 4252 25542 4266 25594
rect 4290 25542 4304 25594
rect 4304 25542 4316 25594
rect 4316 25542 4346 25594
rect 4370 25542 4380 25594
rect 4380 25542 4426 25594
rect 4130 25540 4186 25542
rect 4210 25540 4266 25542
rect 4290 25540 4346 25542
rect 4370 25540 4426 25542
rect 7304 25050 7360 25052
rect 7384 25050 7440 25052
rect 7464 25050 7520 25052
rect 7544 25050 7600 25052
rect 7304 24998 7350 25050
rect 7350 24998 7360 25050
rect 7384 24998 7414 25050
rect 7414 24998 7426 25050
rect 7426 24998 7440 25050
rect 7464 24998 7478 25050
rect 7478 24998 7490 25050
rect 7490 24998 7520 25050
rect 7544 24998 7554 25050
rect 7554 24998 7600 25050
rect 7304 24996 7360 24998
rect 7384 24996 7440 24998
rect 7464 24996 7520 24998
rect 7544 24996 7600 24998
rect 4130 24506 4186 24508
rect 4210 24506 4266 24508
rect 4290 24506 4346 24508
rect 4370 24506 4426 24508
rect 4130 24454 4176 24506
rect 4176 24454 4186 24506
rect 4210 24454 4240 24506
rect 4240 24454 4252 24506
rect 4252 24454 4266 24506
rect 4290 24454 4304 24506
rect 4304 24454 4316 24506
rect 4316 24454 4346 24506
rect 4370 24454 4380 24506
rect 4380 24454 4426 24506
rect 4130 24452 4186 24454
rect 4210 24452 4266 24454
rect 4290 24452 4346 24454
rect 4370 24452 4426 24454
rect 7304 23962 7360 23964
rect 7384 23962 7440 23964
rect 7464 23962 7520 23964
rect 7544 23962 7600 23964
rect 7304 23910 7350 23962
rect 7350 23910 7360 23962
rect 7384 23910 7414 23962
rect 7414 23910 7426 23962
rect 7426 23910 7440 23962
rect 7464 23910 7478 23962
rect 7478 23910 7490 23962
rect 7490 23910 7520 23962
rect 7544 23910 7554 23962
rect 7554 23910 7600 23962
rect 7304 23908 7360 23910
rect 7384 23908 7440 23910
rect 7464 23908 7520 23910
rect 7544 23908 7600 23910
rect 4130 23418 4186 23420
rect 4210 23418 4266 23420
rect 4290 23418 4346 23420
rect 4370 23418 4426 23420
rect 4130 23366 4176 23418
rect 4176 23366 4186 23418
rect 4210 23366 4240 23418
rect 4240 23366 4252 23418
rect 4252 23366 4266 23418
rect 4290 23366 4304 23418
rect 4304 23366 4316 23418
rect 4316 23366 4346 23418
rect 4370 23366 4380 23418
rect 4380 23366 4426 23418
rect 4130 23364 4186 23366
rect 4210 23364 4266 23366
rect 4290 23364 4346 23366
rect 4370 23364 4426 23366
rect 7304 22874 7360 22876
rect 7384 22874 7440 22876
rect 7464 22874 7520 22876
rect 7544 22874 7600 22876
rect 7304 22822 7350 22874
rect 7350 22822 7360 22874
rect 7384 22822 7414 22874
rect 7414 22822 7426 22874
rect 7426 22822 7440 22874
rect 7464 22822 7478 22874
rect 7478 22822 7490 22874
rect 7490 22822 7520 22874
rect 7544 22822 7554 22874
rect 7554 22822 7600 22874
rect 7304 22820 7360 22822
rect 7384 22820 7440 22822
rect 7464 22820 7520 22822
rect 7544 22820 7600 22822
rect 10478 25594 10534 25596
rect 10558 25594 10614 25596
rect 10638 25594 10694 25596
rect 10718 25594 10774 25596
rect 10478 25542 10524 25594
rect 10524 25542 10534 25594
rect 10558 25542 10588 25594
rect 10588 25542 10600 25594
rect 10600 25542 10614 25594
rect 10638 25542 10652 25594
rect 10652 25542 10664 25594
rect 10664 25542 10694 25594
rect 10718 25542 10728 25594
rect 10728 25542 10774 25594
rect 10478 25540 10534 25542
rect 10558 25540 10614 25542
rect 10638 25540 10694 25542
rect 10718 25540 10774 25542
rect 10478 24506 10534 24508
rect 10558 24506 10614 24508
rect 10638 24506 10694 24508
rect 10718 24506 10774 24508
rect 10478 24454 10524 24506
rect 10524 24454 10534 24506
rect 10558 24454 10588 24506
rect 10588 24454 10600 24506
rect 10600 24454 10614 24506
rect 10638 24454 10652 24506
rect 10652 24454 10664 24506
rect 10664 24454 10694 24506
rect 10718 24454 10728 24506
rect 10728 24454 10774 24506
rect 10478 24452 10534 24454
rect 10558 24452 10614 24454
rect 10638 24452 10694 24454
rect 10718 24452 10774 24454
rect 10478 23418 10534 23420
rect 10558 23418 10614 23420
rect 10638 23418 10694 23420
rect 10718 23418 10774 23420
rect 10478 23366 10524 23418
rect 10524 23366 10534 23418
rect 10558 23366 10588 23418
rect 10588 23366 10600 23418
rect 10600 23366 10614 23418
rect 10638 23366 10652 23418
rect 10652 23366 10664 23418
rect 10664 23366 10694 23418
rect 10718 23366 10728 23418
rect 10728 23366 10774 23418
rect 10478 23364 10534 23366
rect 10558 23364 10614 23366
rect 10638 23364 10694 23366
rect 10718 23364 10774 23366
rect 12438 25880 12494 25936
rect 12254 25780 12256 25800
rect 12256 25780 12308 25800
rect 12308 25780 12310 25800
rect 12254 25744 12310 25780
rect 13652 26138 13708 26140
rect 13732 26138 13788 26140
rect 13812 26138 13868 26140
rect 13892 26138 13948 26140
rect 13652 26086 13698 26138
rect 13698 26086 13708 26138
rect 13732 26086 13762 26138
rect 13762 26086 13774 26138
rect 13774 26086 13788 26138
rect 13812 26086 13826 26138
rect 13826 26086 13838 26138
rect 13838 26086 13868 26138
rect 13892 26086 13902 26138
rect 13902 26086 13948 26138
rect 13652 26084 13708 26086
rect 13732 26084 13788 26086
rect 13812 26084 13868 26086
rect 13892 26084 13948 26086
rect 13634 25880 13690 25936
rect 14462 25780 14464 25800
rect 14464 25780 14516 25800
rect 14516 25780 14518 25800
rect 14462 25744 14518 25780
rect 13652 25050 13708 25052
rect 13732 25050 13788 25052
rect 13812 25050 13868 25052
rect 13892 25050 13948 25052
rect 13652 24998 13698 25050
rect 13698 24998 13708 25050
rect 13732 24998 13762 25050
rect 13762 24998 13774 25050
rect 13774 24998 13788 25050
rect 13812 24998 13826 25050
rect 13826 24998 13838 25050
rect 13838 24998 13868 25050
rect 13892 24998 13902 25050
rect 13902 24998 13948 25050
rect 13652 24996 13708 24998
rect 13732 24996 13788 24998
rect 13812 24996 13868 24998
rect 13892 24996 13948 24998
rect 4130 22330 4186 22332
rect 4210 22330 4266 22332
rect 4290 22330 4346 22332
rect 4370 22330 4426 22332
rect 4130 22278 4176 22330
rect 4176 22278 4186 22330
rect 4210 22278 4240 22330
rect 4240 22278 4252 22330
rect 4252 22278 4266 22330
rect 4290 22278 4304 22330
rect 4304 22278 4316 22330
rect 4316 22278 4346 22330
rect 4370 22278 4380 22330
rect 4380 22278 4426 22330
rect 4130 22276 4186 22278
rect 4210 22276 4266 22278
rect 4290 22276 4346 22278
rect 4370 22276 4426 22278
rect 7304 21786 7360 21788
rect 7384 21786 7440 21788
rect 7464 21786 7520 21788
rect 7544 21786 7600 21788
rect 7304 21734 7350 21786
rect 7350 21734 7360 21786
rect 7384 21734 7414 21786
rect 7414 21734 7426 21786
rect 7426 21734 7440 21786
rect 7464 21734 7478 21786
rect 7478 21734 7490 21786
rect 7490 21734 7520 21786
rect 7544 21734 7554 21786
rect 7554 21734 7600 21786
rect 7304 21732 7360 21734
rect 7384 21732 7440 21734
rect 7464 21732 7520 21734
rect 7544 21732 7600 21734
rect 4130 21242 4186 21244
rect 4210 21242 4266 21244
rect 4290 21242 4346 21244
rect 4370 21242 4426 21244
rect 4130 21190 4176 21242
rect 4176 21190 4186 21242
rect 4210 21190 4240 21242
rect 4240 21190 4252 21242
rect 4252 21190 4266 21242
rect 4290 21190 4304 21242
rect 4304 21190 4316 21242
rect 4316 21190 4346 21242
rect 4370 21190 4380 21242
rect 4380 21190 4426 21242
rect 4130 21188 4186 21190
rect 4210 21188 4266 21190
rect 4290 21188 4346 21190
rect 4370 21188 4426 21190
rect 7304 20698 7360 20700
rect 7384 20698 7440 20700
rect 7464 20698 7520 20700
rect 7544 20698 7600 20700
rect 7304 20646 7350 20698
rect 7350 20646 7360 20698
rect 7384 20646 7414 20698
rect 7414 20646 7426 20698
rect 7426 20646 7440 20698
rect 7464 20646 7478 20698
rect 7478 20646 7490 20698
rect 7490 20646 7520 20698
rect 7544 20646 7554 20698
rect 7554 20646 7600 20698
rect 7304 20644 7360 20646
rect 7384 20644 7440 20646
rect 7464 20644 7520 20646
rect 7544 20644 7600 20646
rect 4130 20154 4186 20156
rect 4210 20154 4266 20156
rect 4290 20154 4346 20156
rect 4370 20154 4426 20156
rect 4130 20102 4176 20154
rect 4176 20102 4186 20154
rect 4210 20102 4240 20154
rect 4240 20102 4252 20154
rect 4252 20102 4266 20154
rect 4290 20102 4304 20154
rect 4304 20102 4316 20154
rect 4316 20102 4346 20154
rect 4370 20102 4380 20154
rect 4380 20102 4426 20154
rect 4130 20100 4186 20102
rect 4210 20100 4266 20102
rect 4290 20100 4346 20102
rect 4370 20100 4426 20102
rect 8574 20440 8630 20496
rect 938 19116 940 19136
rect 940 19116 992 19136
rect 992 19116 994 19136
rect 938 19080 994 19116
rect 4130 19066 4186 19068
rect 4210 19066 4266 19068
rect 4290 19066 4346 19068
rect 4370 19066 4426 19068
rect 4130 19014 4176 19066
rect 4176 19014 4186 19066
rect 4210 19014 4240 19066
rect 4240 19014 4252 19066
rect 4252 19014 4266 19066
rect 4290 19014 4304 19066
rect 4304 19014 4316 19066
rect 4316 19014 4346 19066
rect 4370 19014 4380 19066
rect 4380 19014 4426 19066
rect 4130 19012 4186 19014
rect 4210 19012 4266 19014
rect 4290 19012 4346 19014
rect 4370 19012 4426 19014
rect 4130 17978 4186 17980
rect 4210 17978 4266 17980
rect 4290 17978 4346 17980
rect 4370 17978 4426 17980
rect 4130 17926 4176 17978
rect 4176 17926 4186 17978
rect 4210 17926 4240 17978
rect 4240 17926 4252 17978
rect 4252 17926 4266 17978
rect 4290 17926 4304 17978
rect 4304 17926 4316 17978
rect 4316 17926 4346 17978
rect 4370 17926 4380 17978
rect 4380 17926 4426 17978
rect 4130 17924 4186 17926
rect 4210 17924 4266 17926
rect 4290 17924 4346 17926
rect 4370 17924 4426 17926
rect 4130 16890 4186 16892
rect 4210 16890 4266 16892
rect 4290 16890 4346 16892
rect 4370 16890 4426 16892
rect 4130 16838 4176 16890
rect 4176 16838 4186 16890
rect 4210 16838 4240 16890
rect 4240 16838 4252 16890
rect 4252 16838 4266 16890
rect 4290 16838 4304 16890
rect 4304 16838 4316 16890
rect 4316 16838 4346 16890
rect 4370 16838 4380 16890
rect 4380 16838 4426 16890
rect 4130 16836 4186 16838
rect 4210 16836 4266 16838
rect 4290 16836 4346 16838
rect 4370 16836 4426 16838
rect 1398 15136 1454 15192
rect 4130 15802 4186 15804
rect 4210 15802 4266 15804
rect 4290 15802 4346 15804
rect 4370 15802 4426 15804
rect 4130 15750 4176 15802
rect 4176 15750 4186 15802
rect 4210 15750 4240 15802
rect 4240 15750 4252 15802
rect 4252 15750 4266 15802
rect 4290 15750 4304 15802
rect 4304 15750 4316 15802
rect 4316 15750 4346 15802
rect 4370 15750 4380 15802
rect 4380 15750 4426 15802
rect 4130 15748 4186 15750
rect 4210 15748 4266 15750
rect 4290 15748 4346 15750
rect 4370 15748 4426 15750
rect 4130 14714 4186 14716
rect 4210 14714 4266 14716
rect 4290 14714 4346 14716
rect 4370 14714 4426 14716
rect 4130 14662 4176 14714
rect 4176 14662 4186 14714
rect 4210 14662 4240 14714
rect 4240 14662 4252 14714
rect 4252 14662 4266 14714
rect 4290 14662 4304 14714
rect 4304 14662 4316 14714
rect 4316 14662 4346 14714
rect 4370 14662 4380 14714
rect 4380 14662 4426 14714
rect 4130 14660 4186 14662
rect 4210 14660 4266 14662
rect 4290 14660 4346 14662
rect 4370 14660 4426 14662
rect 4130 13626 4186 13628
rect 4210 13626 4266 13628
rect 4290 13626 4346 13628
rect 4370 13626 4426 13628
rect 4130 13574 4176 13626
rect 4176 13574 4186 13626
rect 4210 13574 4240 13626
rect 4240 13574 4252 13626
rect 4252 13574 4266 13626
rect 4290 13574 4304 13626
rect 4304 13574 4316 13626
rect 4316 13574 4346 13626
rect 4370 13574 4380 13626
rect 4380 13574 4426 13626
rect 4130 13572 4186 13574
rect 4210 13572 4266 13574
rect 4290 13572 4346 13574
rect 4370 13572 4426 13574
rect 4130 12538 4186 12540
rect 4210 12538 4266 12540
rect 4290 12538 4346 12540
rect 4370 12538 4426 12540
rect 4130 12486 4176 12538
rect 4176 12486 4186 12538
rect 4210 12486 4240 12538
rect 4240 12486 4252 12538
rect 4252 12486 4266 12538
rect 4290 12486 4304 12538
rect 4304 12486 4316 12538
rect 4316 12486 4346 12538
rect 4370 12486 4380 12538
rect 4380 12486 4426 12538
rect 4130 12484 4186 12486
rect 4210 12484 4266 12486
rect 4290 12484 4346 12486
rect 4370 12484 4426 12486
rect 7304 19610 7360 19612
rect 7384 19610 7440 19612
rect 7464 19610 7520 19612
rect 7544 19610 7600 19612
rect 7304 19558 7350 19610
rect 7350 19558 7360 19610
rect 7384 19558 7414 19610
rect 7414 19558 7426 19610
rect 7426 19558 7440 19610
rect 7464 19558 7478 19610
rect 7478 19558 7490 19610
rect 7490 19558 7520 19610
rect 7544 19558 7554 19610
rect 7554 19558 7600 19610
rect 7304 19556 7360 19558
rect 7384 19556 7440 19558
rect 7464 19556 7520 19558
rect 7544 19556 7600 19558
rect 7304 18522 7360 18524
rect 7384 18522 7440 18524
rect 7464 18522 7520 18524
rect 7544 18522 7600 18524
rect 7304 18470 7350 18522
rect 7350 18470 7360 18522
rect 7384 18470 7414 18522
rect 7414 18470 7426 18522
rect 7426 18470 7440 18522
rect 7464 18470 7478 18522
rect 7478 18470 7490 18522
rect 7490 18470 7520 18522
rect 7544 18470 7554 18522
rect 7554 18470 7600 18522
rect 7304 18468 7360 18470
rect 7384 18468 7440 18470
rect 7464 18468 7520 18470
rect 7544 18468 7600 18470
rect 10478 22330 10534 22332
rect 10558 22330 10614 22332
rect 10638 22330 10694 22332
rect 10718 22330 10774 22332
rect 10478 22278 10524 22330
rect 10524 22278 10534 22330
rect 10558 22278 10588 22330
rect 10588 22278 10600 22330
rect 10600 22278 10614 22330
rect 10638 22278 10652 22330
rect 10652 22278 10664 22330
rect 10664 22278 10694 22330
rect 10718 22278 10728 22330
rect 10728 22278 10774 22330
rect 10478 22276 10534 22278
rect 10558 22276 10614 22278
rect 10638 22276 10694 22278
rect 10718 22276 10774 22278
rect 10478 21242 10534 21244
rect 10558 21242 10614 21244
rect 10638 21242 10694 21244
rect 10718 21242 10774 21244
rect 10478 21190 10524 21242
rect 10524 21190 10534 21242
rect 10558 21190 10588 21242
rect 10588 21190 10600 21242
rect 10600 21190 10614 21242
rect 10638 21190 10652 21242
rect 10652 21190 10664 21242
rect 10664 21190 10694 21242
rect 10718 21190 10728 21242
rect 10728 21190 10774 21242
rect 10478 21188 10534 21190
rect 10558 21188 10614 21190
rect 10638 21188 10694 21190
rect 10718 21188 10774 21190
rect 13652 23962 13708 23964
rect 13732 23962 13788 23964
rect 13812 23962 13868 23964
rect 13892 23962 13948 23964
rect 13652 23910 13698 23962
rect 13698 23910 13708 23962
rect 13732 23910 13762 23962
rect 13762 23910 13774 23962
rect 13774 23910 13788 23962
rect 13812 23910 13826 23962
rect 13826 23910 13838 23962
rect 13838 23910 13868 23962
rect 13892 23910 13902 23962
rect 13902 23910 13948 23962
rect 13652 23908 13708 23910
rect 13732 23908 13788 23910
rect 13812 23908 13868 23910
rect 13892 23908 13948 23910
rect 13652 22874 13708 22876
rect 13732 22874 13788 22876
rect 13812 22874 13868 22876
rect 13892 22874 13948 22876
rect 13652 22822 13698 22874
rect 13698 22822 13708 22874
rect 13732 22822 13762 22874
rect 13762 22822 13774 22874
rect 13774 22822 13788 22874
rect 13812 22822 13826 22874
rect 13826 22822 13838 22874
rect 13838 22822 13868 22874
rect 13892 22822 13902 22874
rect 13902 22822 13948 22874
rect 13652 22820 13708 22822
rect 13732 22820 13788 22822
rect 13812 22820 13868 22822
rect 13892 22820 13948 22822
rect 16826 26682 16882 26684
rect 16906 26682 16962 26684
rect 16986 26682 17042 26684
rect 17066 26682 17122 26684
rect 16826 26630 16872 26682
rect 16872 26630 16882 26682
rect 16906 26630 16936 26682
rect 16936 26630 16948 26682
rect 16948 26630 16962 26682
rect 16986 26630 17000 26682
rect 17000 26630 17012 26682
rect 17012 26630 17042 26682
rect 17066 26630 17076 26682
rect 17076 26630 17122 26682
rect 16826 26628 16882 26630
rect 16906 26628 16962 26630
rect 16986 26628 17042 26630
rect 17066 26628 17122 26630
rect 16826 25594 16882 25596
rect 16906 25594 16962 25596
rect 16986 25594 17042 25596
rect 17066 25594 17122 25596
rect 16826 25542 16872 25594
rect 16872 25542 16882 25594
rect 16906 25542 16936 25594
rect 16936 25542 16948 25594
rect 16948 25542 16962 25594
rect 16986 25542 17000 25594
rect 17000 25542 17012 25594
rect 17012 25542 17042 25594
rect 17066 25542 17076 25594
rect 17076 25542 17122 25594
rect 16826 25540 16882 25542
rect 16906 25540 16962 25542
rect 16986 25540 17042 25542
rect 17066 25540 17122 25542
rect 16826 24506 16882 24508
rect 16906 24506 16962 24508
rect 16986 24506 17042 24508
rect 17066 24506 17122 24508
rect 16826 24454 16872 24506
rect 16872 24454 16882 24506
rect 16906 24454 16936 24506
rect 16936 24454 16948 24506
rect 16948 24454 16962 24506
rect 16986 24454 17000 24506
rect 17000 24454 17012 24506
rect 17012 24454 17042 24506
rect 17066 24454 17076 24506
rect 17076 24454 17122 24506
rect 16826 24452 16882 24454
rect 16906 24452 16962 24454
rect 16986 24452 17042 24454
rect 17066 24452 17122 24454
rect 13652 21786 13708 21788
rect 13732 21786 13788 21788
rect 13812 21786 13868 21788
rect 13892 21786 13948 21788
rect 13652 21734 13698 21786
rect 13698 21734 13708 21786
rect 13732 21734 13762 21786
rect 13762 21734 13774 21786
rect 13774 21734 13788 21786
rect 13812 21734 13826 21786
rect 13826 21734 13838 21786
rect 13838 21734 13868 21786
rect 13892 21734 13902 21786
rect 13902 21734 13948 21786
rect 13652 21732 13708 21734
rect 13732 21732 13788 21734
rect 13812 21732 13868 21734
rect 13892 21732 13948 21734
rect 11610 20476 11612 20496
rect 11612 20476 11664 20496
rect 11664 20476 11666 20496
rect 7304 17434 7360 17436
rect 7384 17434 7440 17436
rect 7464 17434 7520 17436
rect 7544 17434 7600 17436
rect 7304 17382 7350 17434
rect 7350 17382 7360 17434
rect 7384 17382 7414 17434
rect 7414 17382 7426 17434
rect 7426 17382 7440 17434
rect 7464 17382 7478 17434
rect 7478 17382 7490 17434
rect 7490 17382 7520 17434
rect 7544 17382 7554 17434
rect 7554 17382 7600 17434
rect 7304 17380 7360 17382
rect 7384 17380 7440 17382
rect 7464 17380 7520 17382
rect 7544 17380 7600 17382
rect 7304 16346 7360 16348
rect 7384 16346 7440 16348
rect 7464 16346 7520 16348
rect 7544 16346 7600 16348
rect 7304 16294 7350 16346
rect 7350 16294 7360 16346
rect 7384 16294 7414 16346
rect 7414 16294 7426 16346
rect 7426 16294 7440 16346
rect 7464 16294 7478 16346
rect 7478 16294 7490 16346
rect 7490 16294 7520 16346
rect 7544 16294 7554 16346
rect 7554 16294 7600 16346
rect 7304 16292 7360 16294
rect 7384 16292 7440 16294
rect 7464 16292 7520 16294
rect 7544 16292 7600 16294
rect 4130 11450 4186 11452
rect 4210 11450 4266 11452
rect 4290 11450 4346 11452
rect 4370 11450 4426 11452
rect 4130 11398 4176 11450
rect 4176 11398 4186 11450
rect 4210 11398 4240 11450
rect 4240 11398 4252 11450
rect 4252 11398 4266 11450
rect 4290 11398 4304 11450
rect 4304 11398 4316 11450
rect 4316 11398 4346 11450
rect 4370 11398 4380 11450
rect 4380 11398 4426 11450
rect 4130 11396 4186 11398
rect 4210 11396 4266 11398
rect 4290 11396 4346 11398
rect 4370 11396 4426 11398
rect 4130 10362 4186 10364
rect 4210 10362 4266 10364
rect 4290 10362 4346 10364
rect 4370 10362 4426 10364
rect 4130 10310 4176 10362
rect 4176 10310 4186 10362
rect 4210 10310 4240 10362
rect 4240 10310 4252 10362
rect 4252 10310 4266 10362
rect 4290 10310 4304 10362
rect 4304 10310 4316 10362
rect 4316 10310 4346 10362
rect 4370 10310 4380 10362
rect 4380 10310 4426 10362
rect 4130 10308 4186 10310
rect 4210 10308 4266 10310
rect 4290 10308 4346 10310
rect 4370 10308 4426 10310
rect 11610 20440 11666 20476
rect 10478 20154 10534 20156
rect 10558 20154 10614 20156
rect 10638 20154 10694 20156
rect 10718 20154 10774 20156
rect 10478 20102 10524 20154
rect 10524 20102 10534 20154
rect 10558 20102 10588 20154
rect 10588 20102 10600 20154
rect 10600 20102 10614 20154
rect 10638 20102 10652 20154
rect 10652 20102 10664 20154
rect 10664 20102 10694 20154
rect 10718 20102 10728 20154
rect 10728 20102 10774 20154
rect 10478 20100 10534 20102
rect 10558 20100 10614 20102
rect 10638 20100 10694 20102
rect 10718 20100 10774 20102
rect 10414 19236 10470 19272
rect 10414 19216 10416 19236
rect 10416 19216 10468 19236
rect 10468 19216 10470 19236
rect 10478 19066 10534 19068
rect 10558 19066 10614 19068
rect 10638 19066 10694 19068
rect 10718 19066 10774 19068
rect 10478 19014 10524 19066
rect 10524 19014 10534 19066
rect 10558 19014 10588 19066
rect 10588 19014 10600 19066
rect 10600 19014 10614 19066
rect 10638 19014 10652 19066
rect 10652 19014 10664 19066
rect 10664 19014 10694 19066
rect 10718 19014 10728 19066
rect 10728 19014 10774 19066
rect 10478 19012 10534 19014
rect 10558 19012 10614 19014
rect 10638 19012 10694 19014
rect 10718 19012 10774 19014
rect 10478 17978 10534 17980
rect 10558 17978 10614 17980
rect 10638 17978 10694 17980
rect 10718 17978 10774 17980
rect 10478 17926 10524 17978
rect 10524 17926 10534 17978
rect 10558 17926 10588 17978
rect 10588 17926 10600 17978
rect 10600 17926 10614 17978
rect 10638 17926 10652 17978
rect 10652 17926 10664 17978
rect 10664 17926 10694 17978
rect 10718 17926 10728 17978
rect 10728 17926 10774 17978
rect 10478 17924 10534 17926
rect 10558 17924 10614 17926
rect 10638 17924 10694 17926
rect 10718 17924 10774 17926
rect 13652 20698 13708 20700
rect 13732 20698 13788 20700
rect 13812 20698 13868 20700
rect 13892 20698 13948 20700
rect 13652 20646 13698 20698
rect 13698 20646 13708 20698
rect 13732 20646 13762 20698
rect 13762 20646 13774 20698
rect 13774 20646 13788 20698
rect 13812 20646 13826 20698
rect 13826 20646 13838 20698
rect 13838 20646 13868 20698
rect 13892 20646 13902 20698
rect 13902 20646 13948 20698
rect 13652 20644 13708 20646
rect 13732 20644 13788 20646
rect 13812 20644 13868 20646
rect 13892 20644 13948 20646
rect 10478 16890 10534 16892
rect 10558 16890 10614 16892
rect 10638 16890 10694 16892
rect 10718 16890 10774 16892
rect 10478 16838 10524 16890
rect 10524 16838 10534 16890
rect 10558 16838 10588 16890
rect 10588 16838 10600 16890
rect 10600 16838 10614 16890
rect 10638 16838 10652 16890
rect 10652 16838 10664 16890
rect 10664 16838 10694 16890
rect 10718 16838 10728 16890
rect 10728 16838 10774 16890
rect 10478 16836 10534 16838
rect 10558 16836 10614 16838
rect 10638 16836 10694 16838
rect 10718 16836 10774 16838
rect 12622 19216 12678 19272
rect 13652 19610 13708 19612
rect 13732 19610 13788 19612
rect 13812 19610 13868 19612
rect 13892 19610 13948 19612
rect 13652 19558 13698 19610
rect 13698 19558 13708 19610
rect 13732 19558 13762 19610
rect 13762 19558 13774 19610
rect 13774 19558 13788 19610
rect 13812 19558 13826 19610
rect 13826 19558 13838 19610
rect 13838 19558 13868 19610
rect 13892 19558 13902 19610
rect 13902 19558 13948 19610
rect 13652 19556 13708 19558
rect 13732 19556 13788 19558
rect 13812 19556 13868 19558
rect 13892 19556 13948 19558
rect 13652 18522 13708 18524
rect 13732 18522 13788 18524
rect 13812 18522 13868 18524
rect 13892 18522 13948 18524
rect 13652 18470 13698 18522
rect 13698 18470 13708 18522
rect 13732 18470 13762 18522
rect 13762 18470 13774 18522
rect 13774 18470 13788 18522
rect 13812 18470 13826 18522
rect 13826 18470 13838 18522
rect 13838 18470 13868 18522
rect 13892 18470 13902 18522
rect 13902 18470 13948 18522
rect 13652 18468 13708 18470
rect 13732 18468 13788 18470
rect 13812 18468 13868 18470
rect 13892 18468 13948 18470
rect 7304 15258 7360 15260
rect 7384 15258 7440 15260
rect 7464 15258 7520 15260
rect 7544 15258 7600 15260
rect 7304 15206 7350 15258
rect 7350 15206 7360 15258
rect 7384 15206 7414 15258
rect 7414 15206 7426 15258
rect 7426 15206 7440 15258
rect 7464 15206 7478 15258
rect 7478 15206 7490 15258
rect 7490 15206 7520 15258
rect 7544 15206 7554 15258
rect 7554 15206 7600 15258
rect 7304 15204 7360 15206
rect 7384 15204 7440 15206
rect 7464 15204 7520 15206
rect 7544 15204 7600 15206
rect 7304 14170 7360 14172
rect 7384 14170 7440 14172
rect 7464 14170 7520 14172
rect 7544 14170 7600 14172
rect 7304 14118 7350 14170
rect 7350 14118 7360 14170
rect 7384 14118 7414 14170
rect 7414 14118 7426 14170
rect 7426 14118 7440 14170
rect 7464 14118 7478 14170
rect 7478 14118 7490 14170
rect 7490 14118 7520 14170
rect 7544 14118 7554 14170
rect 7554 14118 7600 14170
rect 7304 14116 7360 14118
rect 7384 14116 7440 14118
rect 7464 14116 7520 14118
rect 7544 14116 7600 14118
rect 10478 15802 10534 15804
rect 10558 15802 10614 15804
rect 10638 15802 10694 15804
rect 10718 15802 10774 15804
rect 10478 15750 10524 15802
rect 10524 15750 10534 15802
rect 10558 15750 10588 15802
rect 10588 15750 10600 15802
rect 10600 15750 10614 15802
rect 10638 15750 10652 15802
rect 10652 15750 10664 15802
rect 10664 15750 10694 15802
rect 10718 15750 10728 15802
rect 10728 15750 10774 15802
rect 10478 15748 10534 15750
rect 10558 15748 10614 15750
rect 10638 15748 10694 15750
rect 10718 15748 10774 15750
rect 7304 13082 7360 13084
rect 7384 13082 7440 13084
rect 7464 13082 7520 13084
rect 7544 13082 7600 13084
rect 7304 13030 7350 13082
rect 7350 13030 7360 13082
rect 7384 13030 7414 13082
rect 7414 13030 7426 13082
rect 7426 13030 7440 13082
rect 7464 13030 7478 13082
rect 7478 13030 7490 13082
rect 7490 13030 7520 13082
rect 7544 13030 7554 13082
rect 7554 13030 7600 13082
rect 7304 13028 7360 13030
rect 7384 13028 7440 13030
rect 7464 13028 7520 13030
rect 7544 13028 7600 13030
rect 7304 11994 7360 11996
rect 7384 11994 7440 11996
rect 7464 11994 7520 11996
rect 7544 11994 7600 11996
rect 7304 11942 7350 11994
rect 7350 11942 7360 11994
rect 7384 11942 7414 11994
rect 7414 11942 7426 11994
rect 7426 11942 7440 11994
rect 7464 11942 7478 11994
rect 7478 11942 7490 11994
rect 7490 11942 7520 11994
rect 7544 11942 7554 11994
rect 7554 11942 7600 11994
rect 7304 11940 7360 11942
rect 7384 11940 7440 11942
rect 7464 11940 7520 11942
rect 7544 11940 7600 11942
rect 7304 10906 7360 10908
rect 7384 10906 7440 10908
rect 7464 10906 7520 10908
rect 7544 10906 7600 10908
rect 7304 10854 7350 10906
rect 7350 10854 7360 10906
rect 7384 10854 7414 10906
rect 7414 10854 7426 10906
rect 7426 10854 7440 10906
rect 7464 10854 7478 10906
rect 7478 10854 7490 10906
rect 7490 10854 7520 10906
rect 7544 10854 7554 10906
rect 7554 10854 7600 10906
rect 7304 10852 7360 10854
rect 7384 10852 7440 10854
rect 7464 10852 7520 10854
rect 7544 10852 7600 10854
rect 4130 9274 4186 9276
rect 4210 9274 4266 9276
rect 4290 9274 4346 9276
rect 4370 9274 4426 9276
rect 4130 9222 4176 9274
rect 4176 9222 4186 9274
rect 4210 9222 4240 9274
rect 4240 9222 4252 9274
rect 4252 9222 4266 9274
rect 4290 9222 4304 9274
rect 4304 9222 4316 9274
rect 4316 9222 4346 9274
rect 4370 9222 4380 9274
rect 4380 9222 4426 9274
rect 4130 9220 4186 9222
rect 4210 9220 4266 9222
rect 4290 9220 4346 9222
rect 4370 9220 4426 9222
rect 4130 8186 4186 8188
rect 4210 8186 4266 8188
rect 4290 8186 4346 8188
rect 4370 8186 4426 8188
rect 4130 8134 4176 8186
rect 4176 8134 4186 8186
rect 4210 8134 4240 8186
rect 4240 8134 4252 8186
rect 4252 8134 4266 8186
rect 4290 8134 4304 8186
rect 4304 8134 4316 8186
rect 4316 8134 4346 8186
rect 4370 8134 4380 8186
rect 4380 8134 4426 8186
rect 4130 8132 4186 8134
rect 4210 8132 4266 8134
rect 4290 8132 4346 8134
rect 4370 8132 4426 8134
rect 4066 7520 4122 7576
rect 4130 7098 4186 7100
rect 4210 7098 4266 7100
rect 4290 7098 4346 7100
rect 4370 7098 4426 7100
rect 4130 7046 4176 7098
rect 4176 7046 4186 7098
rect 4210 7046 4240 7098
rect 4240 7046 4252 7098
rect 4252 7046 4266 7098
rect 4290 7046 4304 7098
rect 4304 7046 4316 7098
rect 4316 7046 4346 7098
rect 4370 7046 4380 7098
rect 4380 7046 4426 7098
rect 4130 7044 4186 7046
rect 4210 7044 4266 7046
rect 4290 7044 4346 7046
rect 4370 7044 4426 7046
rect 7304 9818 7360 9820
rect 7384 9818 7440 9820
rect 7464 9818 7520 9820
rect 7544 9818 7600 9820
rect 7304 9766 7350 9818
rect 7350 9766 7360 9818
rect 7384 9766 7414 9818
rect 7414 9766 7426 9818
rect 7426 9766 7440 9818
rect 7464 9766 7478 9818
rect 7478 9766 7490 9818
rect 7490 9766 7520 9818
rect 7544 9766 7554 9818
rect 7554 9766 7600 9818
rect 7304 9764 7360 9766
rect 7384 9764 7440 9766
rect 7464 9764 7520 9766
rect 7544 9764 7600 9766
rect 4130 6010 4186 6012
rect 4210 6010 4266 6012
rect 4290 6010 4346 6012
rect 4370 6010 4426 6012
rect 4130 5958 4176 6010
rect 4176 5958 4186 6010
rect 4210 5958 4240 6010
rect 4240 5958 4252 6010
rect 4252 5958 4266 6010
rect 4290 5958 4304 6010
rect 4304 5958 4316 6010
rect 4316 5958 4346 6010
rect 4370 5958 4380 6010
rect 4380 5958 4426 6010
rect 4130 5956 4186 5958
rect 4210 5956 4266 5958
rect 4290 5956 4346 5958
rect 4370 5956 4426 5958
rect 4130 4922 4186 4924
rect 4210 4922 4266 4924
rect 4290 4922 4346 4924
rect 4370 4922 4426 4924
rect 4130 4870 4176 4922
rect 4176 4870 4186 4922
rect 4210 4870 4240 4922
rect 4240 4870 4252 4922
rect 4252 4870 4266 4922
rect 4290 4870 4304 4922
rect 4304 4870 4316 4922
rect 4316 4870 4346 4922
rect 4370 4870 4380 4922
rect 4380 4870 4426 4922
rect 4130 4868 4186 4870
rect 4210 4868 4266 4870
rect 4290 4868 4346 4870
rect 4370 4868 4426 4870
rect 4130 3834 4186 3836
rect 4210 3834 4266 3836
rect 4290 3834 4346 3836
rect 4370 3834 4426 3836
rect 4130 3782 4176 3834
rect 4176 3782 4186 3834
rect 4210 3782 4240 3834
rect 4240 3782 4252 3834
rect 4252 3782 4266 3834
rect 4290 3782 4304 3834
rect 4304 3782 4316 3834
rect 4316 3782 4346 3834
rect 4370 3782 4380 3834
rect 4380 3782 4426 3834
rect 4130 3780 4186 3782
rect 4210 3780 4266 3782
rect 4290 3780 4346 3782
rect 4370 3780 4426 3782
rect 7304 8730 7360 8732
rect 7384 8730 7440 8732
rect 7464 8730 7520 8732
rect 7544 8730 7600 8732
rect 7304 8678 7350 8730
rect 7350 8678 7360 8730
rect 7384 8678 7414 8730
rect 7414 8678 7426 8730
rect 7426 8678 7440 8730
rect 7464 8678 7478 8730
rect 7478 8678 7490 8730
rect 7490 8678 7520 8730
rect 7544 8678 7554 8730
rect 7554 8678 7600 8730
rect 7304 8676 7360 8678
rect 7384 8676 7440 8678
rect 7464 8676 7520 8678
rect 7544 8676 7600 8678
rect 10478 14714 10534 14716
rect 10558 14714 10614 14716
rect 10638 14714 10694 14716
rect 10718 14714 10774 14716
rect 10478 14662 10524 14714
rect 10524 14662 10534 14714
rect 10558 14662 10588 14714
rect 10588 14662 10600 14714
rect 10600 14662 10614 14714
rect 10638 14662 10652 14714
rect 10652 14662 10664 14714
rect 10664 14662 10694 14714
rect 10718 14662 10728 14714
rect 10728 14662 10774 14714
rect 10478 14660 10534 14662
rect 10558 14660 10614 14662
rect 10638 14660 10694 14662
rect 10718 14660 10774 14662
rect 10478 13626 10534 13628
rect 10558 13626 10614 13628
rect 10638 13626 10694 13628
rect 10718 13626 10774 13628
rect 10478 13574 10524 13626
rect 10524 13574 10534 13626
rect 10558 13574 10588 13626
rect 10588 13574 10600 13626
rect 10600 13574 10614 13626
rect 10638 13574 10652 13626
rect 10652 13574 10664 13626
rect 10664 13574 10694 13626
rect 10718 13574 10728 13626
rect 10728 13574 10774 13626
rect 10478 13572 10534 13574
rect 10558 13572 10614 13574
rect 10638 13572 10694 13574
rect 10718 13572 10774 13574
rect 12622 16088 12678 16144
rect 7304 7642 7360 7644
rect 7384 7642 7440 7644
rect 7464 7642 7520 7644
rect 7544 7642 7600 7644
rect 7304 7590 7350 7642
rect 7350 7590 7360 7642
rect 7384 7590 7414 7642
rect 7414 7590 7426 7642
rect 7426 7590 7440 7642
rect 7464 7590 7478 7642
rect 7478 7590 7490 7642
rect 7490 7590 7520 7642
rect 7544 7590 7554 7642
rect 7554 7590 7600 7642
rect 7304 7588 7360 7590
rect 7384 7588 7440 7590
rect 7464 7588 7520 7590
rect 7544 7588 7600 7590
rect 7304 6554 7360 6556
rect 7384 6554 7440 6556
rect 7464 6554 7520 6556
rect 7544 6554 7600 6556
rect 7304 6502 7350 6554
rect 7350 6502 7360 6554
rect 7384 6502 7414 6554
rect 7414 6502 7426 6554
rect 7426 6502 7440 6554
rect 7464 6502 7478 6554
rect 7478 6502 7490 6554
rect 7490 6502 7520 6554
rect 7544 6502 7554 6554
rect 7554 6502 7600 6554
rect 7304 6500 7360 6502
rect 7384 6500 7440 6502
rect 7464 6500 7520 6502
rect 7544 6500 7600 6502
rect 10478 12538 10534 12540
rect 10558 12538 10614 12540
rect 10638 12538 10694 12540
rect 10718 12538 10774 12540
rect 10478 12486 10524 12538
rect 10524 12486 10534 12538
rect 10558 12486 10588 12538
rect 10588 12486 10600 12538
rect 10600 12486 10614 12538
rect 10638 12486 10652 12538
rect 10652 12486 10664 12538
rect 10664 12486 10694 12538
rect 10718 12486 10728 12538
rect 10728 12486 10774 12538
rect 10478 12484 10534 12486
rect 10558 12484 10614 12486
rect 10638 12484 10694 12486
rect 10718 12484 10774 12486
rect 10478 11450 10534 11452
rect 10558 11450 10614 11452
rect 10638 11450 10694 11452
rect 10718 11450 10774 11452
rect 10478 11398 10524 11450
rect 10524 11398 10534 11450
rect 10558 11398 10588 11450
rect 10588 11398 10600 11450
rect 10600 11398 10614 11450
rect 10638 11398 10652 11450
rect 10652 11398 10664 11450
rect 10664 11398 10694 11450
rect 10718 11398 10728 11450
rect 10728 11398 10774 11450
rect 10478 11396 10534 11398
rect 10558 11396 10614 11398
rect 10638 11396 10694 11398
rect 10718 11396 10774 11398
rect 10478 10362 10534 10364
rect 10558 10362 10614 10364
rect 10638 10362 10694 10364
rect 10718 10362 10774 10364
rect 10478 10310 10524 10362
rect 10524 10310 10534 10362
rect 10558 10310 10588 10362
rect 10588 10310 10600 10362
rect 10600 10310 10614 10362
rect 10638 10310 10652 10362
rect 10652 10310 10664 10362
rect 10664 10310 10694 10362
rect 10718 10310 10728 10362
rect 10728 10310 10774 10362
rect 10478 10308 10534 10310
rect 10558 10308 10614 10310
rect 10638 10308 10694 10310
rect 10718 10308 10774 10310
rect 10478 9274 10534 9276
rect 10558 9274 10614 9276
rect 10638 9274 10694 9276
rect 10718 9274 10774 9276
rect 10478 9222 10524 9274
rect 10524 9222 10534 9274
rect 10558 9222 10588 9274
rect 10588 9222 10600 9274
rect 10600 9222 10614 9274
rect 10638 9222 10652 9274
rect 10652 9222 10664 9274
rect 10664 9222 10694 9274
rect 10718 9222 10728 9274
rect 10728 9222 10774 9274
rect 10478 9220 10534 9222
rect 10558 9220 10614 9222
rect 10638 9220 10694 9222
rect 10718 9220 10774 9222
rect 13652 17434 13708 17436
rect 13732 17434 13788 17436
rect 13812 17434 13868 17436
rect 13892 17434 13948 17436
rect 13652 17382 13698 17434
rect 13698 17382 13708 17434
rect 13732 17382 13762 17434
rect 13762 17382 13774 17434
rect 13774 17382 13788 17434
rect 13812 17382 13826 17434
rect 13826 17382 13838 17434
rect 13838 17382 13868 17434
rect 13892 17382 13902 17434
rect 13902 17382 13948 17434
rect 13652 17380 13708 17382
rect 13732 17380 13788 17382
rect 13812 17380 13868 17382
rect 13892 17380 13948 17382
rect 13652 16346 13708 16348
rect 13732 16346 13788 16348
rect 13812 16346 13868 16348
rect 13892 16346 13948 16348
rect 13652 16294 13698 16346
rect 13698 16294 13708 16346
rect 13732 16294 13762 16346
rect 13762 16294 13774 16346
rect 13774 16294 13788 16346
rect 13812 16294 13826 16346
rect 13826 16294 13838 16346
rect 13838 16294 13868 16346
rect 13892 16294 13902 16346
rect 13902 16294 13948 16346
rect 13652 16292 13708 16294
rect 13732 16292 13788 16294
rect 13812 16292 13868 16294
rect 13892 16292 13948 16294
rect 16826 23418 16882 23420
rect 16906 23418 16962 23420
rect 16986 23418 17042 23420
rect 17066 23418 17122 23420
rect 16826 23366 16872 23418
rect 16872 23366 16882 23418
rect 16906 23366 16936 23418
rect 16936 23366 16948 23418
rect 16948 23366 16962 23418
rect 16986 23366 17000 23418
rect 17000 23366 17012 23418
rect 17012 23366 17042 23418
rect 17066 23366 17076 23418
rect 17076 23366 17122 23418
rect 16826 23364 16882 23366
rect 16906 23364 16962 23366
rect 16986 23364 17042 23366
rect 17066 23364 17122 23366
rect 16826 22330 16882 22332
rect 16906 22330 16962 22332
rect 16986 22330 17042 22332
rect 17066 22330 17122 22332
rect 16826 22278 16872 22330
rect 16872 22278 16882 22330
rect 16906 22278 16936 22330
rect 16936 22278 16948 22330
rect 16948 22278 16962 22330
rect 16986 22278 17000 22330
rect 17000 22278 17012 22330
rect 17012 22278 17042 22330
rect 17066 22278 17076 22330
rect 17076 22278 17122 22330
rect 16826 22276 16882 22278
rect 16906 22276 16962 22278
rect 16986 22276 17042 22278
rect 17066 22276 17122 22278
rect 14646 16088 14702 16144
rect 13652 15258 13708 15260
rect 13732 15258 13788 15260
rect 13812 15258 13868 15260
rect 13892 15258 13948 15260
rect 13652 15206 13698 15258
rect 13698 15206 13708 15258
rect 13732 15206 13762 15258
rect 13762 15206 13774 15258
rect 13774 15206 13788 15258
rect 13812 15206 13826 15258
rect 13826 15206 13838 15258
rect 13838 15206 13868 15258
rect 13892 15206 13902 15258
rect 13902 15206 13948 15258
rect 13652 15204 13708 15206
rect 13732 15204 13788 15206
rect 13812 15204 13868 15206
rect 13892 15204 13948 15206
rect 13652 14170 13708 14172
rect 13732 14170 13788 14172
rect 13812 14170 13868 14172
rect 13892 14170 13948 14172
rect 13652 14118 13698 14170
rect 13698 14118 13708 14170
rect 13732 14118 13762 14170
rect 13762 14118 13774 14170
rect 13774 14118 13788 14170
rect 13812 14118 13826 14170
rect 13826 14118 13838 14170
rect 13838 14118 13868 14170
rect 13892 14118 13902 14170
rect 13902 14118 13948 14170
rect 13652 14116 13708 14118
rect 13732 14116 13788 14118
rect 13812 14116 13868 14118
rect 13892 14116 13948 14118
rect 13652 13082 13708 13084
rect 13732 13082 13788 13084
rect 13812 13082 13868 13084
rect 13892 13082 13948 13084
rect 13652 13030 13698 13082
rect 13698 13030 13708 13082
rect 13732 13030 13762 13082
rect 13762 13030 13774 13082
rect 13774 13030 13788 13082
rect 13812 13030 13826 13082
rect 13826 13030 13838 13082
rect 13838 13030 13868 13082
rect 13892 13030 13902 13082
rect 13902 13030 13948 13082
rect 13652 13028 13708 13030
rect 13732 13028 13788 13030
rect 13812 13028 13868 13030
rect 13892 13028 13948 13030
rect 13652 11994 13708 11996
rect 13732 11994 13788 11996
rect 13812 11994 13868 11996
rect 13892 11994 13948 11996
rect 13652 11942 13698 11994
rect 13698 11942 13708 11994
rect 13732 11942 13762 11994
rect 13762 11942 13774 11994
rect 13774 11942 13788 11994
rect 13812 11942 13826 11994
rect 13826 11942 13838 11994
rect 13838 11942 13868 11994
rect 13892 11942 13902 11994
rect 13902 11942 13948 11994
rect 13652 11940 13708 11942
rect 13732 11940 13788 11942
rect 13812 11940 13868 11942
rect 13892 11940 13948 11942
rect 13652 10906 13708 10908
rect 13732 10906 13788 10908
rect 13812 10906 13868 10908
rect 13892 10906 13948 10908
rect 13652 10854 13698 10906
rect 13698 10854 13708 10906
rect 13732 10854 13762 10906
rect 13762 10854 13774 10906
rect 13774 10854 13788 10906
rect 13812 10854 13826 10906
rect 13826 10854 13838 10906
rect 13838 10854 13868 10906
rect 13892 10854 13902 10906
rect 13902 10854 13948 10906
rect 13652 10852 13708 10854
rect 13732 10852 13788 10854
rect 13812 10852 13868 10854
rect 13892 10852 13948 10854
rect 11150 8744 11206 8800
rect 10478 8186 10534 8188
rect 10558 8186 10614 8188
rect 10638 8186 10694 8188
rect 10718 8186 10774 8188
rect 10478 8134 10524 8186
rect 10524 8134 10534 8186
rect 10558 8134 10588 8186
rect 10588 8134 10600 8186
rect 10600 8134 10614 8186
rect 10638 8134 10652 8186
rect 10652 8134 10664 8186
rect 10664 8134 10694 8186
rect 10718 8134 10728 8186
rect 10728 8134 10774 8186
rect 10478 8132 10534 8134
rect 10558 8132 10614 8134
rect 10638 8132 10694 8134
rect 10718 8132 10774 8134
rect 10478 7098 10534 7100
rect 10558 7098 10614 7100
rect 10638 7098 10694 7100
rect 10718 7098 10774 7100
rect 10478 7046 10524 7098
rect 10524 7046 10534 7098
rect 10558 7046 10588 7098
rect 10588 7046 10600 7098
rect 10600 7046 10614 7098
rect 10638 7046 10652 7098
rect 10652 7046 10664 7098
rect 10664 7046 10694 7098
rect 10718 7046 10728 7098
rect 10728 7046 10774 7098
rect 10478 7044 10534 7046
rect 10558 7044 10614 7046
rect 10638 7044 10694 7046
rect 10718 7044 10774 7046
rect 7304 5466 7360 5468
rect 7384 5466 7440 5468
rect 7464 5466 7520 5468
rect 7544 5466 7600 5468
rect 7304 5414 7350 5466
rect 7350 5414 7360 5466
rect 7384 5414 7414 5466
rect 7414 5414 7426 5466
rect 7426 5414 7440 5466
rect 7464 5414 7478 5466
rect 7478 5414 7490 5466
rect 7490 5414 7520 5466
rect 7544 5414 7554 5466
rect 7554 5414 7600 5466
rect 7304 5412 7360 5414
rect 7384 5412 7440 5414
rect 7464 5412 7520 5414
rect 7544 5412 7600 5414
rect 7304 4378 7360 4380
rect 7384 4378 7440 4380
rect 7464 4378 7520 4380
rect 7544 4378 7600 4380
rect 7304 4326 7350 4378
rect 7350 4326 7360 4378
rect 7384 4326 7414 4378
rect 7414 4326 7426 4378
rect 7426 4326 7440 4378
rect 7464 4326 7478 4378
rect 7478 4326 7490 4378
rect 7490 4326 7520 4378
rect 7544 4326 7554 4378
rect 7554 4326 7600 4378
rect 7304 4324 7360 4326
rect 7384 4324 7440 4326
rect 7464 4324 7520 4326
rect 7544 4324 7600 4326
rect 7304 3290 7360 3292
rect 7384 3290 7440 3292
rect 7464 3290 7520 3292
rect 7544 3290 7600 3292
rect 7304 3238 7350 3290
rect 7350 3238 7360 3290
rect 7384 3238 7414 3290
rect 7414 3238 7426 3290
rect 7426 3238 7440 3290
rect 7464 3238 7478 3290
rect 7478 3238 7490 3290
rect 7490 3238 7520 3290
rect 7544 3238 7554 3290
rect 7554 3238 7600 3290
rect 7304 3236 7360 3238
rect 7384 3236 7440 3238
rect 7464 3236 7520 3238
rect 7544 3236 7600 3238
rect 12438 9016 12494 9072
rect 12898 8780 12900 8800
rect 12900 8780 12952 8800
rect 12952 8780 12954 8800
rect 12898 8744 12954 8780
rect 10478 6010 10534 6012
rect 10558 6010 10614 6012
rect 10638 6010 10694 6012
rect 10718 6010 10774 6012
rect 10478 5958 10524 6010
rect 10524 5958 10534 6010
rect 10558 5958 10588 6010
rect 10588 5958 10600 6010
rect 10600 5958 10614 6010
rect 10638 5958 10652 6010
rect 10652 5958 10664 6010
rect 10664 5958 10694 6010
rect 10718 5958 10728 6010
rect 10728 5958 10774 6010
rect 10478 5956 10534 5958
rect 10558 5956 10614 5958
rect 10638 5956 10694 5958
rect 10718 5956 10774 5958
rect 13652 9818 13708 9820
rect 13732 9818 13788 9820
rect 13812 9818 13868 9820
rect 13892 9818 13948 9820
rect 13652 9766 13698 9818
rect 13698 9766 13708 9818
rect 13732 9766 13762 9818
rect 13762 9766 13774 9818
rect 13774 9766 13788 9818
rect 13812 9766 13826 9818
rect 13826 9766 13838 9818
rect 13838 9766 13868 9818
rect 13892 9766 13902 9818
rect 13902 9766 13948 9818
rect 13652 9764 13708 9766
rect 13732 9764 13788 9766
rect 13812 9764 13868 9766
rect 13892 9764 13948 9766
rect 13358 9016 13414 9072
rect 13652 8730 13708 8732
rect 13732 8730 13788 8732
rect 13812 8730 13868 8732
rect 13892 8730 13948 8732
rect 13652 8678 13698 8730
rect 13698 8678 13708 8730
rect 13732 8678 13762 8730
rect 13762 8678 13774 8730
rect 13774 8678 13788 8730
rect 13812 8678 13826 8730
rect 13826 8678 13838 8730
rect 13838 8678 13868 8730
rect 13892 8678 13902 8730
rect 13902 8678 13948 8730
rect 13652 8676 13708 8678
rect 13732 8676 13788 8678
rect 13812 8676 13868 8678
rect 13892 8676 13948 8678
rect 16762 21548 16818 21584
rect 16762 21528 16764 21548
rect 16764 21528 16816 21548
rect 16816 21528 16818 21548
rect 17682 21528 17738 21584
rect 17222 21412 17278 21448
rect 17222 21392 17224 21412
rect 17224 21392 17276 21412
rect 17276 21392 17278 21412
rect 16826 21242 16882 21244
rect 16906 21242 16962 21244
rect 16986 21242 17042 21244
rect 17066 21242 17122 21244
rect 16826 21190 16872 21242
rect 16872 21190 16882 21242
rect 16906 21190 16936 21242
rect 16936 21190 16948 21242
rect 16948 21190 16962 21242
rect 16986 21190 17000 21242
rect 17000 21190 17012 21242
rect 17012 21190 17042 21242
rect 17066 21190 17076 21242
rect 17076 21190 17122 21242
rect 16826 21188 16882 21190
rect 16906 21188 16962 21190
rect 16986 21188 17042 21190
rect 17066 21188 17122 21190
rect 16946 20576 17002 20632
rect 16826 20154 16882 20156
rect 16906 20154 16962 20156
rect 16986 20154 17042 20156
rect 17066 20154 17122 20156
rect 16826 20102 16872 20154
rect 16872 20102 16882 20154
rect 16906 20102 16936 20154
rect 16936 20102 16948 20154
rect 16948 20102 16962 20154
rect 16986 20102 17000 20154
rect 17000 20102 17012 20154
rect 17012 20102 17042 20154
rect 17066 20102 17076 20154
rect 17076 20102 17122 20154
rect 16826 20100 16882 20102
rect 16906 20100 16962 20102
rect 16986 20100 17042 20102
rect 17066 20100 17122 20102
rect 16826 19066 16882 19068
rect 16906 19066 16962 19068
rect 16986 19066 17042 19068
rect 17066 19066 17122 19068
rect 16826 19014 16872 19066
rect 16872 19014 16882 19066
rect 16906 19014 16936 19066
rect 16936 19014 16948 19066
rect 16948 19014 16962 19066
rect 16986 19014 17000 19066
rect 17000 19014 17012 19066
rect 17012 19014 17042 19066
rect 17066 19014 17076 19066
rect 17076 19014 17122 19066
rect 16826 19012 16882 19014
rect 16906 19012 16962 19014
rect 16986 19012 17042 19014
rect 17066 19012 17122 19014
rect 20000 26138 20056 26140
rect 20080 26138 20136 26140
rect 20160 26138 20216 26140
rect 20240 26138 20296 26140
rect 20000 26086 20046 26138
rect 20046 26086 20056 26138
rect 20080 26086 20110 26138
rect 20110 26086 20122 26138
rect 20122 26086 20136 26138
rect 20160 26086 20174 26138
rect 20174 26086 20186 26138
rect 20186 26086 20216 26138
rect 20240 26086 20250 26138
rect 20250 26086 20296 26138
rect 20000 26084 20056 26086
rect 20080 26084 20136 26086
rect 20160 26084 20216 26086
rect 20240 26084 20296 26086
rect 20000 25050 20056 25052
rect 20080 25050 20136 25052
rect 20160 25050 20216 25052
rect 20240 25050 20296 25052
rect 20000 24998 20046 25050
rect 20046 24998 20056 25050
rect 20080 24998 20110 25050
rect 20110 24998 20122 25050
rect 20122 24998 20136 25050
rect 20160 24998 20174 25050
rect 20174 24998 20186 25050
rect 20186 24998 20216 25050
rect 20240 24998 20250 25050
rect 20250 24998 20296 25050
rect 20000 24996 20056 24998
rect 20080 24996 20136 24998
rect 20160 24996 20216 24998
rect 20240 24996 20296 24998
rect 20000 23962 20056 23964
rect 20080 23962 20136 23964
rect 20160 23962 20216 23964
rect 20240 23962 20296 23964
rect 20000 23910 20046 23962
rect 20046 23910 20056 23962
rect 20080 23910 20110 23962
rect 20110 23910 20122 23962
rect 20122 23910 20136 23962
rect 20160 23910 20174 23962
rect 20174 23910 20186 23962
rect 20186 23910 20216 23962
rect 20240 23910 20250 23962
rect 20250 23910 20296 23962
rect 20000 23908 20056 23910
rect 20080 23908 20136 23910
rect 20160 23908 20216 23910
rect 20240 23908 20296 23910
rect 23174 26682 23230 26684
rect 23254 26682 23310 26684
rect 23334 26682 23390 26684
rect 23414 26682 23470 26684
rect 23174 26630 23220 26682
rect 23220 26630 23230 26682
rect 23254 26630 23284 26682
rect 23284 26630 23296 26682
rect 23296 26630 23310 26682
rect 23334 26630 23348 26682
rect 23348 26630 23360 26682
rect 23360 26630 23390 26682
rect 23414 26630 23424 26682
rect 23424 26630 23470 26682
rect 23174 26628 23230 26630
rect 23254 26628 23310 26630
rect 23334 26628 23390 26630
rect 23414 26628 23470 26630
rect 26348 26138 26404 26140
rect 26428 26138 26484 26140
rect 26508 26138 26564 26140
rect 26588 26138 26644 26140
rect 26348 26086 26394 26138
rect 26394 26086 26404 26138
rect 26428 26086 26458 26138
rect 26458 26086 26470 26138
rect 26470 26086 26484 26138
rect 26508 26086 26522 26138
rect 26522 26086 26534 26138
rect 26534 26086 26564 26138
rect 26588 26086 26598 26138
rect 26598 26086 26644 26138
rect 26348 26084 26404 26086
rect 26428 26084 26484 26086
rect 26508 26084 26564 26086
rect 26588 26084 26644 26086
rect 23174 25594 23230 25596
rect 23254 25594 23310 25596
rect 23334 25594 23390 25596
rect 23414 25594 23470 25596
rect 23174 25542 23220 25594
rect 23220 25542 23230 25594
rect 23254 25542 23284 25594
rect 23284 25542 23296 25594
rect 23296 25542 23310 25594
rect 23334 25542 23348 25594
rect 23348 25542 23360 25594
rect 23360 25542 23390 25594
rect 23414 25542 23424 25594
rect 23424 25542 23470 25594
rect 23174 25540 23230 25542
rect 23254 25540 23310 25542
rect 23334 25540 23390 25542
rect 23414 25540 23470 25542
rect 20000 22874 20056 22876
rect 20080 22874 20136 22876
rect 20160 22874 20216 22876
rect 20240 22874 20296 22876
rect 20000 22822 20046 22874
rect 20046 22822 20056 22874
rect 20080 22822 20110 22874
rect 20110 22822 20122 22874
rect 20122 22822 20136 22874
rect 20160 22822 20174 22874
rect 20174 22822 20186 22874
rect 20186 22822 20216 22874
rect 20240 22822 20250 22874
rect 20250 22822 20296 22874
rect 20000 22820 20056 22822
rect 20080 22820 20136 22822
rect 20160 22820 20216 22822
rect 20240 22820 20296 22822
rect 20000 21786 20056 21788
rect 20080 21786 20136 21788
rect 20160 21786 20216 21788
rect 20240 21786 20296 21788
rect 20000 21734 20046 21786
rect 20046 21734 20056 21786
rect 20080 21734 20110 21786
rect 20110 21734 20122 21786
rect 20122 21734 20136 21786
rect 20160 21734 20174 21786
rect 20174 21734 20186 21786
rect 20186 21734 20216 21786
rect 20240 21734 20250 21786
rect 20250 21734 20296 21786
rect 20000 21732 20056 21734
rect 20080 21732 20136 21734
rect 20160 21732 20216 21734
rect 20240 21732 20296 21734
rect 18326 21548 18382 21584
rect 18326 21528 18328 21548
rect 18328 21528 18380 21548
rect 18380 21528 18382 21548
rect 18602 21412 18658 21448
rect 18602 21392 18604 21412
rect 18604 21392 18656 21412
rect 18656 21392 18658 21412
rect 18510 20596 18566 20632
rect 18510 20576 18512 20596
rect 18512 20576 18564 20596
rect 18564 20576 18566 20596
rect 20000 20698 20056 20700
rect 20080 20698 20136 20700
rect 20160 20698 20216 20700
rect 20240 20698 20296 20700
rect 20000 20646 20046 20698
rect 20046 20646 20056 20698
rect 20080 20646 20110 20698
rect 20110 20646 20122 20698
rect 20122 20646 20136 20698
rect 20160 20646 20174 20698
rect 20174 20646 20186 20698
rect 20186 20646 20216 20698
rect 20240 20646 20250 20698
rect 20250 20646 20296 20698
rect 20000 20644 20056 20646
rect 20080 20644 20136 20646
rect 20160 20644 20216 20646
rect 20240 20644 20296 20646
rect 16826 17978 16882 17980
rect 16906 17978 16962 17980
rect 16986 17978 17042 17980
rect 17066 17978 17122 17980
rect 16826 17926 16872 17978
rect 16872 17926 16882 17978
rect 16906 17926 16936 17978
rect 16936 17926 16948 17978
rect 16948 17926 16962 17978
rect 16986 17926 17000 17978
rect 17000 17926 17012 17978
rect 17012 17926 17042 17978
rect 17066 17926 17076 17978
rect 17076 17926 17122 17978
rect 16826 17924 16882 17926
rect 16906 17924 16962 17926
rect 16986 17924 17042 17926
rect 17066 17924 17122 17926
rect 15750 17040 15806 17096
rect 15106 11736 15162 11792
rect 14186 11192 14242 11248
rect 14554 11056 14610 11112
rect 13652 7642 13708 7644
rect 13732 7642 13788 7644
rect 13812 7642 13868 7644
rect 13892 7642 13948 7644
rect 13652 7590 13698 7642
rect 13698 7590 13708 7642
rect 13732 7590 13762 7642
rect 13762 7590 13774 7642
rect 13774 7590 13788 7642
rect 13812 7590 13826 7642
rect 13826 7590 13838 7642
rect 13838 7590 13868 7642
rect 13892 7590 13902 7642
rect 13902 7590 13948 7642
rect 13652 7588 13708 7590
rect 13732 7588 13788 7590
rect 13812 7588 13868 7590
rect 13892 7588 13948 7590
rect 10478 4922 10534 4924
rect 10558 4922 10614 4924
rect 10638 4922 10694 4924
rect 10718 4922 10774 4924
rect 10478 4870 10524 4922
rect 10524 4870 10534 4922
rect 10558 4870 10588 4922
rect 10588 4870 10600 4922
rect 10600 4870 10614 4922
rect 10638 4870 10652 4922
rect 10652 4870 10664 4922
rect 10664 4870 10694 4922
rect 10718 4870 10728 4922
rect 10728 4870 10774 4922
rect 10478 4868 10534 4870
rect 10558 4868 10614 4870
rect 10638 4868 10694 4870
rect 10718 4868 10774 4870
rect 10478 3834 10534 3836
rect 10558 3834 10614 3836
rect 10638 3834 10694 3836
rect 10718 3834 10774 3836
rect 10478 3782 10524 3834
rect 10524 3782 10534 3834
rect 10558 3782 10588 3834
rect 10588 3782 10600 3834
rect 10600 3782 10614 3834
rect 10638 3782 10652 3834
rect 10652 3782 10664 3834
rect 10664 3782 10694 3834
rect 10718 3782 10728 3834
rect 10728 3782 10774 3834
rect 10478 3780 10534 3782
rect 10558 3780 10614 3782
rect 10638 3780 10694 3782
rect 10718 3780 10774 3782
rect 4130 2746 4186 2748
rect 4210 2746 4266 2748
rect 4290 2746 4346 2748
rect 4370 2746 4426 2748
rect 4130 2694 4176 2746
rect 4176 2694 4186 2746
rect 4210 2694 4240 2746
rect 4240 2694 4252 2746
rect 4252 2694 4266 2746
rect 4290 2694 4304 2746
rect 4304 2694 4316 2746
rect 4316 2694 4346 2746
rect 4370 2694 4380 2746
rect 4380 2694 4426 2746
rect 4130 2692 4186 2694
rect 4210 2692 4266 2694
rect 4290 2692 4346 2694
rect 4370 2692 4426 2694
rect 13652 6554 13708 6556
rect 13732 6554 13788 6556
rect 13812 6554 13868 6556
rect 13892 6554 13948 6556
rect 13652 6502 13698 6554
rect 13698 6502 13708 6554
rect 13732 6502 13762 6554
rect 13762 6502 13774 6554
rect 13774 6502 13788 6554
rect 13812 6502 13826 6554
rect 13826 6502 13838 6554
rect 13838 6502 13868 6554
rect 13892 6502 13902 6554
rect 13902 6502 13948 6554
rect 13652 6500 13708 6502
rect 13732 6500 13788 6502
rect 13812 6500 13868 6502
rect 13892 6500 13948 6502
rect 13652 5466 13708 5468
rect 13732 5466 13788 5468
rect 13812 5466 13868 5468
rect 13892 5466 13948 5468
rect 13652 5414 13698 5466
rect 13698 5414 13708 5466
rect 13732 5414 13762 5466
rect 13762 5414 13774 5466
rect 13774 5414 13788 5466
rect 13812 5414 13826 5466
rect 13826 5414 13838 5466
rect 13838 5414 13868 5466
rect 13892 5414 13902 5466
rect 13902 5414 13948 5466
rect 13652 5412 13708 5414
rect 13732 5412 13788 5414
rect 13812 5412 13868 5414
rect 13892 5412 13948 5414
rect 13652 4378 13708 4380
rect 13732 4378 13788 4380
rect 13812 4378 13868 4380
rect 13892 4378 13948 4380
rect 13652 4326 13698 4378
rect 13698 4326 13708 4378
rect 13732 4326 13762 4378
rect 13762 4326 13774 4378
rect 13774 4326 13788 4378
rect 13812 4326 13826 4378
rect 13826 4326 13838 4378
rect 13838 4326 13868 4378
rect 13892 4326 13902 4378
rect 13902 4326 13948 4378
rect 13652 4324 13708 4326
rect 13732 4324 13788 4326
rect 13812 4324 13868 4326
rect 13892 4324 13948 4326
rect 13910 4156 13912 4176
rect 13912 4156 13964 4176
rect 13964 4156 13966 4176
rect 13910 4120 13966 4156
rect 13358 3068 13360 3088
rect 13360 3068 13412 3088
rect 13412 3068 13414 3088
rect 13358 3032 13414 3068
rect 13652 3290 13708 3292
rect 13732 3290 13788 3292
rect 13812 3290 13868 3292
rect 13892 3290 13948 3292
rect 13652 3238 13698 3290
rect 13698 3238 13708 3290
rect 13732 3238 13762 3290
rect 13762 3238 13774 3290
rect 13774 3238 13788 3290
rect 13812 3238 13826 3290
rect 13826 3238 13838 3290
rect 13838 3238 13868 3290
rect 13892 3238 13902 3290
rect 13902 3238 13948 3290
rect 13652 3236 13708 3238
rect 13732 3236 13788 3238
rect 13812 3236 13868 3238
rect 13892 3236 13948 3238
rect 10478 2746 10534 2748
rect 10558 2746 10614 2748
rect 10638 2746 10694 2748
rect 10718 2746 10774 2748
rect 10478 2694 10524 2746
rect 10524 2694 10534 2746
rect 10558 2694 10588 2746
rect 10588 2694 10600 2746
rect 10600 2694 10614 2746
rect 10638 2694 10652 2746
rect 10652 2694 10664 2746
rect 10664 2694 10694 2746
rect 10718 2694 10728 2746
rect 10728 2694 10774 2746
rect 10478 2692 10534 2694
rect 10558 2692 10614 2694
rect 10638 2692 10694 2694
rect 10718 2692 10774 2694
rect 14462 3340 14464 3360
rect 14464 3340 14516 3360
rect 14516 3340 14518 3360
rect 14462 3304 14518 3340
rect 16826 16890 16882 16892
rect 16906 16890 16962 16892
rect 16986 16890 17042 16892
rect 17066 16890 17122 16892
rect 16826 16838 16872 16890
rect 16872 16838 16882 16890
rect 16906 16838 16936 16890
rect 16936 16838 16948 16890
rect 16948 16838 16962 16890
rect 16986 16838 17000 16890
rect 17000 16838 17012 16890
rect 17012 16838 17042 16890
rect 17066 16838 17076 16890
rect 17076 16838 17122 16890
rect 16826 16836 16882 16838
rect 16906 16836 16962 16838
rect 16986 16836 17042 16838
rect 17066 16836 17122 16838
rect 16210 16088 16266 16144
rect 20000 19610 20056 19612
rect 20080 19610 20136 19612
rect 20160 19610 20216 19612
rect 20240 19610 20296 19612
rect 20000 19558 20046 19610
rect 20046 19558 20056 19610
rect 20080 19558 20110 19610
rect 20110 19558 20122 19610
rect 20122 19558 20136 19610
rect 20160 19558 20174 19610
rect 20174 19558 20186 19610
rect 20186 19558 20216 19610
rect 20240 19558 20250 19610
rect 20250 19558 20296 19610
rect 20000 19556 20056 19558
rect 20080 19556 20136 19558
rect 20160 19556 20216 19558
rect 20240 19556 20296 19558
rect 16826 15802 16882 15804
rect 16906 15802 16962 15804
rect 16986 15802 17042 15804
rect 17066 15802 17122 15804
rect 16826 15750 16872 15802
rect 16872 15750 16882 15802
rect 16906 15750 16936 15802
rect 16936 15750 16948 15802
rect 16948 15750 16962 15802
rect 16986 15750 17000 15802
rect 17000 15750 17012 15802
rect 17012 15750 17042 15802
rect 17066 15750 17076 15802
rect 17076 15750 17122 15802
rect 16826 15748 16882 15750
rect 16906 15748 16962 15750
rect 16986 15748 17042 15750
rect 17066 15748 17122 15750
rect 18694 17196 18750 17232
rect 18694 17176 18696 17196
rect 18696 17176 18748 17196
rect 18748 17176 18750 17196
rect 19062 17176 19118 17232
rect 19246 17076 19248 17096
rect 19248 17076 19300 17096
rect 19300 17076 19302 17096
rect 19246 17040 19302 17076
rect 20000 18522 20056 18524
rect 20080 18522 20136 18524
rect 20160 18522 20216 18524
rect 20240 18522 20296 18524
rect 20000 18470 20046 18522
rect 20046 18470 20056 18522
rect 20080 18470 20110 18522
rect 20110 18470 20122 18522
rect 20122 18470 20136 18522
rect 20160 18470 20174 18522
rect 20174 18470 20186 18522
rect 20186 18470 20216 18522
rect 20240 18470 20250 18522
rect 20250 18470 20296 18522
rect 20000 18468 20056 18470
rect 20080 18468 20136 18470
rect 20160 18468 20216 18470
rect 20240 18468 20296 18470
rect 20000 17434 20056 17436
rect 20080 17434 20136 17436
rect 20160 17434 20216 17436
rect 20240 17434 20296 17436
rect 20000 17382 20046 17434
rect 20046 17382 20056 17434
rect 20080 17382 20110 17434
rect 20110 17382 20122 17434
rect 20122 17382 20136 17434
rect 20160 17382 20174 17434
rect 20174 17382 20186 17434
rect 20186 17382 20216 17434
rect 20240 17382 20250 17434
rect 20250 17382 20296 17434
rect 20000 17380 20056 17382
rect 20080 17380 20136 17382
rect 20160 17380 20216 17382
rect 20240 17380 20296 17382
rect 22282 22636 22338 22672
rect 26348 25050 26404 25052
rect 26428 25050 26484 25052
rect 26508 25050 26564 25052
rect 26588 25050 26644 25052
rect 26348 24998 26394 25050
rect 26394 24998 26404 25050
rect 26428 24998 26458 25050
rect 26458 24998 26470 25050
rect 26470 24998 26484 25050
rect 26508 24998 26522 25050
rect 26522 24998 26534 25050
rect 26534 24998 26564 25050
rect 26588 24998 26598 25050
rect 26598 24998 26644 25050
rect 26348 24996 26404 24998
rect 26428 24996 26484 24998
rect 26508 24996 26564 24998
rect 26588 24996 26644 24998
rect 23174 24506 23230 24508
rect 23254 24506 23310 24508
rect 23334 24506 23390 24508
rect 23414 24506 23470 24508
rect 23174 24454 23220 24506
rect 23220 24454 23230 24506
rect 23254 24454 23284 24506
rect 23284 24454 23296 24506
rect 23296 24454 23310 24506
rect 23334 24454 23348 24506
rect 23348 24454 23360 24506
rect 23360 24454 23390 24506
rect 23414 24454 23424 24506
rect 23424 24454 23470 24506
rect 23174 24452 23230 24454
rect 23254 24452 23310 24454
rect 23334 24452 23390 24454
rect 23414 24452 23470 24454
rect 22282 22616 22284 22636
rect 22284 22616 22336 22636
rect 22336 22616 22338 22636
rect 23174 23418 23230 23420
rect 23254 23418 23310 23420
rect 23334 23418 23390 23420
rect 23414 23418 23470 23420
rect 23174 23366 23220 23418
rect 23220 23366 23230 23418
rect 23254 23366 23284 23418
rect 23284 23366 23296 23418
rect 23296 23366 23310 23418
rect 23334 23366 23348 23418
rect 23348 23366 23360 23418
rect 23360 23366 23390 23418
rect 23414 23366 23424 23418
rect 23424 23366 23470 23418
rect 23174 23364 23230 23366
rect 23254 23364 23310 23366
rect 23334 23364 23390 23366
rect 23414 23364 23470 23366
rect 23110 22616 23166 22672
rect 26348 23962 26404 23964
rect 26428 23962 26484 23964
rect 26508 23962 26564 23964
rect 26588 23962 26644 23964
rect 26348 23910 26394 23962
rect 26394 23910 26404 23962
rect 26428 23910 26458 23962
rect 26458 23910 26470 23962
rect 26470 23910 26484 23962
rect 26508 23910 26522 23962
rect 26522 23910 26534 23962
rect 26534 23910 26564 23962
rect 26588 23910 26598 23962
rect 26598 23910 26644 23962
rect 26348 23908 26404 23910
rect 26428 23908 26484 23910
rect 26508 23908 26564 23910
rect 26588 23908 26644 23910
rect 26146 23704 26202 23760
rect 23174 22330 23230 22332
rect 23254 22330 23310 22332
rect 23334 22330 23390 22332
rect 23414 22330 23470 22332
rect 23174 22278 23220 22330
rect 23220 22278 23230 22330
rect 23254 22278 23284 22330
rect 23284 22278 23296 22330
rect 23296 22278 23310 22330
rect 23334 22278 23348 22330
rect 23348 22278 23360 22330
rect 23360 22278 23390 22330
rect 23414 22278 23424 22330
rect 23424 22278 23470 22330
rect 23174 22276 23230 22278
rect 23254 22276 23310 22278
rect 23334 22276 23390 22278
rect 23414 22276 23470 22278
rect 23174 21242 23230 21244
rect 23254 21242 23310 21244
rect 23334 21242 23390 21244
rect 23414 21242 23470 21244
rect 23174 21190 23220 21242
rect 23220 21190 23230 21242
rect 23254 21190 23284 21242
rect 23284 21190 23296 21242
rect 23296 21190 23310 21242
rect 23334 21190 23348 21242
rect 23348 21190 23360 21242
rect 23360 21190 23390 21242
rect 23414 21190 23424 21242
rect 23424 21190 23470 21242
rect 23174 21188 23230 21190
rect 23254 21188 23310 21190
rect 23334 21188 23390 21190
rect 23414 21188 23470 21190
rect 23174 20154 23230 20156
rect 23254 20154 23310 20156
rect 23334 20154 23390 20156
rect 23414 20154 23470 20156
rect 23174 20102 23220 20154
rect 23220 20102 23230 20154
rect 23254 20102 23284 20154
rect 23284 20102 23296 20154
rect 23296 20102 23310 20154
rect 23334 20102 23348 20154
rect 23348 20102 23360 20154
rect 23360 20102 23390 20154
rect 23414 20102 23424 20154
rect 23424 20102 23470 20154
rect 23174 20100 23230 20102
rect 23254 20100 23310 20102
rect 23334 20100 23390 20102
rect 23414 20100 23470 20102
rect 26348 22874 26404 22876
rect 26428 22874 26484 22876
rect 26508 22874 26564 22876
rect 26588 22874 26644 22876
rect 26348 22822 26394 22874
rect 26394 22822 26404 22874
rect 26428 22822 26458 22874
rect 26458 22822 26470 22874
rect 26470 22822 26484 22874
rect 26508 22822 26522 22874
rect 26522 22822 26534 22874
rect 26534 22822 26564 22874
rect 26588 22822 26598 22874
rect 26598 22822 26644 22874
rect 26348 22820 26404 22822
rect 26428 22820 26484 22822
rect 26508 22820 26564 22822
rect 26588 22820 26644 22822
rect 26348 21786 26404 21788
rect 26428 21786 26484 21788
rect 26508 21786 26564 21788
rect 26588 21786 26644 21788
rect 26348 21734 26394 21786
rect 26394 21734 26404 21786
rect 26428 21734 26458 21786
rect 26458 21734 26470 21786
rect 26470 21734 26484 21786
rect 26508 21734 26522 21786
rect 26522 21734 26534 21786
rect 26534 21734 26564 21786
rect 26588 21734 26598 21786
rect 26598 21734 26644 21786
rect 26348 21732 26404 21734
rect 26428 21732 26484 21734
rect 26508 21732 26564 21734
rect 26588 21732 26644 21734
rect 26348 20698 26404 20700
rect 26428 20698 26484 20700
rect 26508 20698 26564 20700
rect 26588 20698 26644 20700
rect 26348 20646 26394 20698
rect 26394 20646 26404 20698
rect 26428 20646 26458 20698
rect 26458 20646 26470 20698
rect 26470 20646 26484 20698
rect 26508 20646 26522 20698
rect 26522 20646 26534 20698
rect 26534 20646 26564 20698
rect 26588 20646 26598 20698
rect 26598 20646 26644 20698
rect 26348 20644 26404 20646
rect 26428 20644 26484 20646
rect 26508 20644 26564 20646
rect 26588 20644 26644 20646
rect 26348 19610 26404 19612
rect 26428 19610 26484 19612
rect 26508 19610 26564 19612
rect 26588 19610 26644 19612
rect 26348 19558 26394 19610
rect 26394 19558 26404 19610
rect 26428 19558 26458 19610
rect 26458 19558 26470 19610
rect 26470 19558 26484 19610
rect 26508 19558 26522 19610
rect 26522 19558 26534 19610
rect 26534 19558 26564 19610
rect 26588 19558 26598 19610
rect 26598 19558 26644 19610
rect 26348 19556 26404 19558
rect 26428 19556 26484 19558
rect 26508 19556 26564 19558
rect 26588 19556 26644 19558
rect 23174 19066 23230 19068
rect 23254 19066 23310 19068
rect 23334 19066 23390 19068
rect 23414 19066 23470 19068
rect 23174 19014 23220 19066
rect 23220 19014 23230 19066
rect 23254 19014 23284 19066
rect 23284 19014 23296 19066
rect 23296 19014 23310 19066
rect 23334 19014 23348 19066
rect 23348 19014 23360 19066
rect 23360 19014 23390 19066
rect 23414 19014 23424 19066
rect 23424 19014 23470 19066
rect 23174 19012 23230 19014
rect 23254 19012 23310 19014
rect 23334 19012 23390 19014
rect 23414 19012 23470 19014
rect 20000 16346 20056 16348
rect 20080 16346 20136 16348
rect 20160 16346 20216 16348
rect 20240 16346 20296 16348
rect 20000 16294 20046 16346
rect 20046 16294 20056 16346
rect 20080 16294 20110 16346
rect 20110 16294 20122 16346
rect 20122 16294 20136 16346
rect 20160 16294 20174 16346
rect 20174 16294 20186 16346
rect 20186 16294 20216 16346
rect 20240 16294 20250 16346
rect 20250 16294 20296 16346
rect 20000 16292 20056 16294
rect 20080 16292 20136 16294
rect 20160 16292 20216 16294
rect 20240 16292 20296 16294
rect 16826 14714 16882 14716
rect 16906 14714 16962 14716
rect 16986 14714 17042 14716
rect 17066 14714 17122 14716
rect 16826 14662 16872 14714
rect 16872 14662 16882 14714
rect 16906 14662 16936 14714
rect 16936 14662 16948 14714
rect 16948 14662 16962 14714
rect 16986 14662 17000 14714
rect 17000 14662 17012 14714
rect 17012 14662 17042 14714
rect 17066 14662 17076 14714
rect 17076 14662 17122 14714
rect 16826 14660 16882 14662
rect 16906 14660 16962 14662
rect 16986 14660 17042 14662
rect 17066 14660 17122 14662
rect 16826 13626 16882 13628
rect 16906 13626 16962 13628
rect 16986 13626 17042 13628
rect 17066 13626 17122 13628
rect 16826 13574 16872 13626
rect 16872 13574 16882 13626
rect 16906 13574 16936 13626
rect 16936 13574 16948 13626
rect 16948 13574 16962 13626
rect 16986 13574 17000 13626
rect 17000 13574 17012 13626
rect 17012 13574 17042 13626
rect 17066 13574 17076 13626
rect 17076 13574 17122 13626
rect 16826 13572 16882 13574
rect 16906 13572 16962 13574
rect 16986 13572 17042 13574
rect 17066 13572 17122 13574
rect 16826 12538 16882 12540
rect 16906 12538 16962 12540
rect 16986 12538 17042 12540
rect 17066 12538 17122 12540
rect 16826 12486 16872 12538
rect 16872 12486 16882 12538
rect 16906 12486 16936 12538
rect 16936 12486 16948 12538
rect 16948 12486 16962 12538
rect 16986 12486 17000 12538
rect 17000 12486 17012 12538
rect 17012 12486 17042 12538
rect 17066 12486 17076 12538
rect 17076 12486 17122 12538
rect 16826 12484 16882 12486
rect 16906 12484 16962 12486
rect 16986 12484 17042 12486
rect 17066 12484 17122 12486
rect 15842 11192 15898 11248
rect 20000 15258 20056 15260
rect 20080 15258 20136 15260
rect 20160 15258 20216 15260
rect 20240 15258 20296 15260
rect 20000 15206 20046 15258
rect 20046 15206 20056 15258
rect 20080 15206 20110 15258
rect 20110 15206 20122 15258
rect 20122 15206 20136 15258
rect 20160 15206 20174 15258
rect 20174 15206 20186 15258
rect 20186 15206 20216 15258
rect 20240 15206 20250 15258
rect 20250 15206 20296 15258
rect 20000 15204 20056 15206
rect 20080 15204 20136 15206
rect 20160 15204 20216 15206
rect 20240 15204 20296 15206
rect 20000 14170 20056 14172
rect 20080 14170 20136 14172
rect 20160 14170 20216 14172
rect 20240 14170 20296 14172
rect 20000 14118 20046 14170
rect 20046 14118 20056 14170
rect 20080 14118 20110 14170
rect 20110 14118 20122 14170
rect 20122 14118 20136 14170
rect 20160 14118 20174 14170
rect 20174 14118 20186 14170
rect 20186 14118 20216 14170
rect 20240 14118 20250 14170
rect 20250 14118 20296 14170
rect 20000 14116 20056 14118
rect 20080 14116 20136 14118
rect 20160 14116 20216 14118
rect 20240 14116 20296 14118
rect 20000 13082 20056 13084
rect 20080 13082 20136 13084
rect 20160 13082 20216 13084
rect 20240 13082 20296 13084
rect 20000 13030 20046 13082
rect 20046 13030 20056 13082
rect 20080 13030 20110 13082
rect 20110 13030 20122 13082
rect 20122 13030 20136 13082
rect 20160 13030 20174 13082
rect 20174 13030 20186 13082
rect 20186 13030 20216 13082
rect 20240 13030 20250 13082
rect 20250 13030 20296 13082
rect 20000 13028 20056 13030
rect 20080 13028 20136 13030
rect 20160 13028 20216 13030
rect 20240 13028 20296 13030
rect 16826 11450 16882 11452
rect 16906 11450 16962 11452
rect 16986 11450 17042 11452
rect 17066 11450 17122 11452
rect 16826 11398 16872 11450
rect 16872 11398 16882 11450
rect 16906 11398 16936 11450
rect 16936 11398 16948 11450
rect 16948 11398 16962 11450
rect 16986 11398 17000 11450
rect 17000 11398 17012 11450
rect 17012 11398 17042 11450
rect 17066 11398 17076 11450
rect 17076 11398 17122 11450
rect 16826 11396 16882 11398
rect 16906 11396 16962 11398
rect 16986 11396 17042 11398
rect 17066 11396 17122 11398
rect 17958 11756 18014 11792
rect 17958 11736 17960 11756
rect 17960 11736 18012 11756
rect 18012 11736 18014 11756
rect 16826 10362 16882 10364
rect 16906 10362 16962 10364
rect 16986 10362 17042 10364
rect 17066 10362 17122 10364
rect 16826 10310 16872 10362
rect 16872 10310 16882 10362
rect 16906 10310 16936 10362
rect 16936 10310 16948 10362
rect 16948 10310 16962 10362
rect 16986 10310 17000 10362
rect 17000 10310 17012 10362
rect 17012 10310 17042 10362
rect 17066 10310 17076 10362
rect 17076 10310 17122 10362
rect 16826 10308 16882 10310
rect 16906 10308 16962 10310
rect 16986 10308 17042 10310
rect 17066 10308 17122 10310
rect 16826 9274 16882 9276
rect 16906 9274 16962 9276
rect 16986 9274 17042 9276
rect 17066 9274 17122 9276
rect 16826 9222 16872 9274
rect 16872 9222 16882 9274
rect 16906 9222 16936 9274
rect 16936 9222 16948 9274
rect 16948 9222 16962 9274
rect 16986 9222 17000 9274
rect 17000 9222 17012 9274
rect 17012 9222 17042 9274
rect 17066 9222 17076 9274
rect 17076 9222 17122 9274
rect 16826 9220 16882 9222
rect 16906 9220 16962 9222
rect 16986 9220 17042 9222
rect 17066 9220 17122 9222
rect 19338 11056 19394 11112
rect 16826 8186 16882 8188
rect 16906 8186 16962 8188
rect 16986 8186 17042 8188
rect 17066 8186 17122 8188
rect 16826 8134 16872 8186
rect 16872 8134 16882 8186
rect 16906 8134 16936 8186
rect 16936 8134 16948 8186
rect 16948 8134 16962 8186
rect 16986 8134 17000 8186
rect 17000 8134 17012 8186
rect 17012 8134 17042 8186
rect 17066 8134 17076 8186
rect 17076 8134 17122 8186
rect 16826 8132 16882 8134
rect 16906 8132 16962 8134
rect 16986 8132 17042 8134
rect 17066 8132 17122 8134
rect 16826 7098 16882 7100
rect 16906 7098 16962 7100
rect 16986 7098 17042 7100
rect 17066 7098 17122 7100
rect 16826 7046 16872 7098
rect 16872 7046 16882 7098
rect 16906 7046 16936 7098
rect 16936 7046 16948 7098
rect 16948 7046 16962 7098
rect 16986 7046 17000 7098
rect 17000 7046 17012 7098
rect 17012 7046 17042 7098
rect 17066 7046 17076 7098
rect 17076 7046 17122 7098
rect 16826 7044 16882 7046
rect 16906 7044 16962 7046
rect 16986 7044 17042 7046
rect 17066 7044 17122 7046
rect 16826 6010 16882 6012
rect 16906 6010 16962 6012
rect 16986 6010 17042 6012
rect 17066 6010 17122 6012
rect 16826 5958 16872 6010
rect 16872 5958 16882 6010
rect 16906 5958 16936 6010
rect 16936 5958 16948 6010
rect 16948 5958 16962 6010
rect 16986 5958 17000 6010
rect 17000 5958 17012 6010
rect 17012 5958 17042 6010
rect 17066 5958 17076 6010
rect 17076 5958 17122 6010
rect 16826 5956 16882 5958
rect 16906 5956 16962 5958
rect 16986 5956 17042 5958
rect 17066 5956 17122 5958
rect 20000 11994 20056 11996
rect 20080 11994 20136 11996
rect 20160 11994 20216 11996
rect 20240 11994 20296 11996
rect 20000 11942 20046 11994
rect 20046 11942 20056 11994
rect 20080 11942 20110 11994
rect 20110 11942 20122 11994
rect 20122 11942 20136 11994
rect 20160 11942 20174 11994
rect 20174 11942 20186 11994
rect 20186 11942 20216 11994
rect 20240 11942 20250 11994
rect 20250 11942 20296 11994
rect 20000 11940 20056 11942
rect 20080 11940 20136 11942
rect 20160 11940 20216 11942
rect 20240 11940 20296 11942
rect 21638 17176 21694 17232
rect 22466 17040 22522 17096
rect 26348 18522 26404 18524
rect 26428 18522 26484 18524
rect 26508 18522 26564 18524
rect 26588 18522 26644 18524
rect 26348 18470 26394 18522
rect 26394 18470 26404 18522
rect 26428 18470 26458 18522
rect 26458 18470 26470 18522
rect 26470 18470 26484 18522
rect 26508 18470 26522 18522
rect 26522 18470 26534 18522
rect 26534 18470 26564 18522
rect 26588 18470 26598 18522
rect 26598 18470 26644 18522
rect 26348 18468 26404 18470
rect 26428 18468 26484 18470
rect 26508 18468 26564 18470
rect 26588 18468 26644 18470
rect 23174 17978 23230 17980
rect 23254 17978 23310 17980
rect 23334 17978 23390 17980
rect 23414 17978 23470 17980
rect 23174 17926 23220 17978
rect 23220 17926 23230 17978
rect 23254 17926 23284 17978
rect 23284 17926 23296 17978
rect 23296 17926 23310 17978
rect 23334 17926 23348 17978
rect 23348 17926 23360 17978
rect 23360 17926 23390 17978
rect 23414 17926 23424 17978
rect 23424 17926 23470 17978
rect 23174 17924 23230 17926
rect 23254 17924 23310 17926
rect 23334 17924 23390 17926
rect 23414 17924 23470 17926
rect 22650 17196 22706 17232
rect 22650 17176 22652 17196
rect 22652 17176 22704 17196
rect 22704 17176 22706 17196
rect 23174 16890 23230 16892
rect 23254 16890 23310 16892
rect 23334 16890 23390 16892
rect 23414 16890 23470 16892
rect 23174 16838 23220 16890
rect 23220 16838 23230 16890
rect 23254 16838 23284 16890
rect 23284 16838 23296 16890
rect 23296 16838 23310 16890
rect 23334 16838 23348 16890
rect 23348 16838 23360 16890
rect 23360 16838 23390 16890
rect 23414 16838 23424 16890
rect 23424 16838 23470 16890
rect 23174 16836 23230 16838
rect 23254 16836 23310 16838
rect 23334 16836 23390 16838
rect 23414 16836 23470 16838
rect 23662 17040 23718 17096
rect 23174 15802 23230 15804
rect 23254 15802 23310 15804
rect 23334 15802 23390 15804
rect 23414 15802 23470 15804
rect 23174 15750 23220 15802
rect 23220 15750 23230 15802
rect 23254 15750 23284 15802
rect 23284 15750 23296 15802
rect 23296 15750 23310 15802
rect 23334 15750 23348 15802
rect 23348 15750 23360 15802
rect 23360 15750 23390 15802
rect 23414 15750 23424 15802
rect 23424 15750 23470 15802
rect 23174 15748 23230 15750
rect 23254 15748 23310 15750
rect 23334 15748 23390 15750
rect 23414 15748 23470 15750
rect 23174 14714 23230 14716
rect 23254 14714 23310 14716
rect 23334 14714 23390 14716
rect 23414 14714 23470 14716
rect 23174 14662 23220 14714
rect 23220 14662 23230 14714
rect 23254 14662 23284 14714
rect 23284 14662 23296 14714
rect 23296 14662 23310 14714
rect 23334 14662 23348 14714
rect 23348 14662 23360 14714
rect 23360 14662 23390 14714
rect 23414 14662 23424 14714
rect 23424 14662 23470 14714
rect 23174 14660 23230 14662
rect 23254 14660 23310 14662
rect 23334 14660 23390 14662
rect 23414 14660 23470 14662
rect 26348 17434 26404 17436
rect 26428 17434 26484 17436
rect 26508 17434 26564 17436
rect 26588 17434 26644 17436
rect 26348 17382 26394 17434
rect 26394 17382 26404 17434
rect 26428 17382 26458 17434
rect 26458 17382 26470 17434
rect 26470 17382 26484 17434
rect 26508 17382 26522 17434
rect 26522 17382 26534 17434
rect 26534 17382 26564 17434
rect 26588 17382 26598 17434
rect 26598 17382 26644 17434
rect 26348 17380 26404 17382
rect 26428 17380 26484 17382
rect 26508 17380 26564 17382
rect 26588 17380 26644 17382
rect 20000 10906 20056 10908
rect 20080 10906 20136 10908
rect 20160 10906 20216 10908
rect 20240 10906 20296 10908
rect 20000 10854 20046 10906
rect 20046 10854 20056 10906
rect 20080 10854 20110 10906
rect 20110 10854 20122 10906
rect 20122 10854 20136 10906
rect 20160 10854 20174 10906
rect 20174 10854 20186 10906
rect 20186 10854 20216 10906
rect 20240 10854 20250 10906
rect 20250 10854 20296 10906
rect 20000 10852 20056 10854
rect 20080 10852 20136 10854
rect 20160 10852 20216 10854
rect 20240 10852 20296 10854
rect 15198 4120 15254 4176
rect 15014 3068 15016 3088
rect 15016 3068 15068 3088
rect 15068 3068 15070 3088
rect 15014 3032 15070 3068
rect 16826 4922 16882 4924
rect 16906 4922 16962 4924
rect 16986 4922 17042 4924
rect 17066 4922 17122 4924
rect 16826 4870 16872 4922
rect 16872 4870 16882 4922
rect 16906 4870 16936 4922
rect 16936 4870 16948 4922
rect 16948 4870 16962 4922
rect 16986 4870 17000 4922
rect 17000 4870 17012 4922
rect 17012 4870 17042 4922
rect 17066 4870 17076 4922
rect 17076 4870 17122 4922
rect 16826 4868 16882 4870
rect 16906 4868 16962 4870
rect 16986 4868 17042 4870
rect 17066 4868 17122 4870
rect 16826 3834 16882 3836
rect 16906 3834 16962 3836
rect 16986 3834 17042 3836
rect 17066 3834 17122 3836
rect 16826 3782 16872 3834
rect 16872 3782 16882 3834
rect 16906 3782 16936 3834
rect 16936 3782 16948 3834
rect 16948 3782 16962 3834
rect 16986 3782 17000 3834
rect 17000 3782 17012 3834
rect 17012 3782 17042 3834
rect 17066 3782 17076 3834
rect 17076 3782 17122 3834
rect 16826 3780 16882 3782
rect 16906 3780 16962 3782
rect 16986 3780 17042 3782
rect 17066 3780 17122 3782
rect 20000 9818 20056 9820
rect 20080 9818 20136 9820
rect 20160 9818 20216 9820
rect 20240 9818 20296 9820
rect 20000 9766 20046 9818
rect 20046 9766 20056 9818
rect 20080 9766 20110 9818
rect 20110 9766 20122 9818
rect 20122 9766 20136 9818
rect 20160 9766 20174 9818
rect 20174 9766 20186 9818
rect 20186 9766 20216 9818
rect 20240 9766 20250 9818
rect 20250 9766 20296 9818
rect 20000 9764 20056 9766
rect 20080 9764 20136 9766
rect 20160 9764 20216 9766
rect 20240 9764 20296 9766
rect 20000 8730 20056 8732
rect 20080 8730 20136 8732
rect 20160 8730 20216 8732
rect 20240 8730 20296 8732
rect 20000 8678 20046 8730
rect 20046 8678 20056 8730
rect 20080 8678 20110 8730
rect 20110 8678 20122 8730
rect 20122 8678 20136 8730
rect 20160 8678 20174 8730
rect 20174 8678 20186 8730
rect 20186 8678 20216 8730
rect 20240 8678 20250 8730
rect 20250 8678 20296 8730
rect 20000 8676 20056 8678
rect 20080 8676 20136 8678
rect 20160 8676 20216 8678
rect 20240 8676 20296 8678
rect 20000 7642 20056 7644
rect 20080 7642 20136 7644
rect 20160 7642 20216 7644
rect 20240 7642 20296 7644
rect 20000 7590 20046 7642
rect 20046 7590 20056 7642
rect 20080 7590 20110 7642
rect 20110 7590 20122 7642
rect 20122 7590 20136 7642
rect 20160 7590 20174 7642
rect 20174 7590 20186 7642
rect 20186 7590 20216 7642
rect 20240 7590 20250 7642
rect 20250 7590 20296 7642
rect 20000 7588 20056 7590
rect 20080 7588 20136 7590
rect 20160 7588 20216 7590
rect 20240 7588 20296 7590
rect 23174 13626 23230 13628
rect 23254 13626 23310 13628
rect 23334 13626 23390 13628
rect 23414 13626 23470 13628
rect 23174 13574 23220 13626
rect 23220 13574 23230 13626
rect 23254 13574 23284 13626
rect 23284 13574 23296 13626
rect 23296 13574 23310 13626
rect 23334 13574 23348 13626
rect 23348 13574 23360 13626
rect 23360 13574 23390 13626
rect 23414 13574 23424 13626
rect 23424 13574 23470 13626
rect 23174 13572 23230 13574
rect 23254 13572 23310 13574
rect 23334 13572 23390 13574
rect 23414 13572 23470 13574
rect 23174 12538 23230 12540
rect 23254 12538 23310 12540
rect 23334 12538 23390 12540
rect 23414 12538 23470 12540
rect 23174 12486 23220 12538
rect 23220 12486 23230 12538
rect 23254 12486 23284 12538
rect 23284 12486 23296 12538
rect 23296 12486 23310 12538
rect 23334 12486 23348 12538
rect 23348 12486 23360 12538
rect 23360 12486 23390 12538
rect 23414 12486 23424 12538
rect 23424 12486 23470 12538
rect 23174 12484 23230 12486
rect 23254 12484 23310 12486
rect 23334 12484 23390 12486
rect 23414 12484 23470 12486
rect 26348 16346 26404 16348
rect 26428 16346 26484 16348
rect 26508 16346 26564 16348
rect 26588 16346 26644 16348
rect 26348 16294 26394 16346
rect 26394 16294 26404 16346
rect 26428 16294 26458 16346
rect 26458 16294 26470 16346
rect 26470 16294 26484 16346
rect 26508 16294 26522 16346
rect 26522 16294 26534 16346
rect 26534 16294 26564 16346
rect 26588 16294 26598 16346
rect 26598 16294 26644 16346
rect 26348 16292 26404 16294
rect 26428 16292 26484 16294
rect 26508 16292 26564 16294
rect 26588 16292 26644 16294
rect 26348 15258 26404 15260
rect 26428 15258 26484 15260
rect 26508 15258 26564 15260
rect 26588 15258 26644 15260
rect 26348 15206 26394 15258
rect 26394 15206 26404 15258
rect 26428 15206 26458 15258
rect 26458 15206 26470 15258
rect 26470 15206 26484 15258
rect 26508 15206 26522 15258
rect 26522 15206 26534 15258
rect 26534 15206 26564 15258
rect 26588 15206 26598 15258
rect 26598 15206 26644 15258
rect 26348 15204 26404 15206
rect 26428 15204 26484 15206
rect 26508 15204 26564 15206
rect 26588 15204 26644 15206
rect 26348 14170 26404 14172
rect 26428 14170 26484 14172
rect 26508 14170 26564 14172
rect 26588 14170 26644 14172
rect 26348 14118 26394 14170
rect 26394 14118 26404 14170
rect 26428 14118 26458 14170
rect 26458 14118 26470 14170
rect 26470 14118 26484 14170
rect 26508 14118 26522 14170
rect 26522 14118 26534 14170
rect 26534 14118 26564 14170
rect 26588 14118 26598 14170
rect 26598 14118 26644 14170
rect 26348 14116 26404 14118
rect 26428 14116 26484 14118
rect 26508 14116 26564 14118
rect 26588 14116 26644 14118
rect 23174 11450 23230 11452
rect 23254 11450 23310 11452
rect 23334 11450 23390 11452
rect 23414 11450 23470 11452
rect 23174 11398 23220 11450
rect 23220 11398 23230 11450
rect 23254 11398 23284 11450
rect 23284 11398 23296 11450
rect 23296 11398 23310 11450
rect 23334 11398 23348 11450
rect 23348 11398 23360 11450
rect 23360 11398 23390 11450
rect 23414 11398 23424 11450
rect 23424 11398 23470 11450
rect 23174 11396 23230 11398
rect 23254 11396 23310 11398
rect 23334 11396 23390 11398
rect 23414 11396 23470 11398
rect 20000 6554 20056 6556
rect 20080 6554 20136 6556
rect 20160 6554 20216 6556
rect 20240 6554 20296 6556
rect 20000 6502 20046 6554
rect 20046 6502 20056 6554
rect 20080 6502 20110 6554
rect 20110 6502 20122 6554
rect 20122 6502 20136 6554
rect 20160 6502 20174 6554
rect 20174 6502 20186 6554
rect 20186 6502 20216 6554
rect 20240 6502 20250 6554
rect 20250 6502 20296 6554
rect 20000 6500 20056 6502
rect 20080 6500 20136 6502
rect 20160 6500 20216 6502
rect 20240 6500 20296 6502
rect 20000 5466 20056 5468
rect 20080 5466 20136 5468
rect 20160 5466 20216 5468
rect 20240 5466 20296 5468
rect 20000 5414 20046 5466
rect 20046 5414 20056 5466
rect 20080 5414 20110 5466
rect 20110 5414 20122 5466
rect 20122 5414 20136 5466
rect 20160 5414 20174 5466
rect 20174 5414 20186 5466
rect 20186 5414 20216 5466
rect 20240 5414 20250 5466
rect 20250 5414 20296 5466
rect 20000 5412 20056 5414
rect 20080 5412 20136 5414
rect 20160 5412 20216 5414
rect 20240 5412 20296 5414
rect 17038 3304 17094 3360
rect 16826 2746 16882 2748
rect 16906 2746 16962 2748
rect 16986 2746 17042 2748
rect 17066 2746 17122 2748
rect 16826 2694 16872 2746
rect 16872 2694 16882 2746
rect 16906 2694 16936 2746
rect 16936 2694 16948 2746
rect 16948 2694 16962 2746
rect 16986 2694 17000 2746
rect 17000 2694 17012 2746
rect 17012 2694 17042 2746
rect 17066 2694 17076 2746
rect 17076 2694 17122 2746
rect 16826 2692 16882 2694
rect 16906 2692 16962 2694
rect 16986 2692 17042 2694
rect 17066 2692 17122 2694
rect 23174 10362 23230 10364
rect 23254 10362 23310 10364
rect 23334 10362 23390 10364
rect 23414 10362 23470 10364
rect 23174 10310 23220 10362
rect 23220 10310 23230 10362
rect 23254 10310 23284 10362
rect 23284 10310 23296 10362
rect 23296 10310 23310 10362
rect 23334 10310 23348 10362
rect 23348 10310 23360 10362
rect 23360 10310 23390 10362
rect 23414 10310 23424 10362
rect 23424 10310 23470 10362
rect 23174 10308 23230 10310
rect 23254 10308 23310 10310
rect 23334 10308 23390 10310
rect 23414 10308 23470 10310
rect 26348 13082 26404 13084
rect 26428 13082 26484 13084
rect 26508 13082 26564 13084
rect 26588 13082 26644 13084
rect 26348 13030 26394 13082
rect 26394 13030 26404 13082
rect 26428 13030 26458 13082
rect 26458 13030 26470 13082
rect 26470 13030 26484 13082
rect 26508 13030 26522 13082
rect 26522 13030 26534 13082
rect 26534 13030 26564 13082
rect 26588 13030 26598 13082
rect 26598 13030 26644 13082
rect 26348 13028 26404 13030
rect 26428 13028 26484 13030
rect 26508 13028 26564 13030
rect 26588 13028 26644 13030
rect 26146 12280 26202 12336
rect 26348 11994 26404 11996
rect 26428 11994 26484 11996
rect 26508 11994 26564 11996
rect 26588 11994 26644 11996
rect 26348 11942 26394 11994
rect 26394 11942 26404 11994
rect 26428 11942 26458 11994
rect 26458 11942 26470 11994
rect 26470 11942 26484 11994
rect 26508 11942 26522 11994
rect 26522 11942 26534 11994
rect 26534 11942 26564 11994
rect 26588 11942 26598 11994
rect 26598 11942 26644 11994
rect 26348 11940 26404 11942
rect 26428 11940 26484 11942
rect 26508 11940 26564 11942
rect 26588 11940 26644 11942
rect 26348 10906 26404 10908
rect 26428 10906 26484 10908
rect 26508 10906 26564 10908
rect 26588 10906 26644 10908
rect 26348 10854 26394 10906
rect 26394 10854 26404 10906
rect 26428 10854 26458 10906
rect 26458 10854 26470 10906
rect 26470 10854 26484 10906
rect 26508 10854 26522 10906
rect 26522 10854 26534 10906
rect 26534 10854 26564 10906
rect 26588 10854 26598 10906
rect 26598 10854 26644 10906
rect 26348 10852 26404 10854
rect 26428 10852 26484 10854
rect 26508 10852 26564 10854
rect 26588 10852 26644 10854
rect 7304 2202 7360 2204
rect 7384 2202 7440 2204
rect 7464 2202 7520 2204
rect 7544 2202 7600 2204
rect 7304 2150 7350 2202
rect 7350 2150 7360 2202
rect 7384 2150 7414 2202
rect 7414 2150 7426 2202
rect 7426 2150 7440 2202
rect 7464 2150 7478 2202
rect 7478 2150 7490 2202
rect 7490 2150 7520 2202
rect 7544 2150 7554 2202
rect 7554 2150 7600 2202
rect 7304 2148 7360 2150
rect 7384 2148 7440 2150
rect 7464 2148 7520 2150
rect 7544 2148 7600 2150
rect 20000 4378 20056 4380
rect 20080 4378 20136 4380
rect 20160 4378 20216 4380
rect 20240 4378 20296 4380
rect 20000 4326 20046 4378
rect 20046 4326 20056 4378
rect 20080 4326 20110 4378
rect 20110 4326 20122 4378
rect 20122 4326 20136 4378
rect 20160 4326 20174 4378
rect 20174 4326 20186 4378
rect 20186 4326 20216 4378
rect 20240 4326 20250 4378
rect 20250 4326 20296 4378
rect 20000 4324 20056 4326
rect 20080 4324 20136 4326
rect 20160 4324 20216 4326
rect 20240 4324 20296 4326
rect 20000 3290 20056 3292
rect 20080 3290 20136 3292
rect 20160 3290 20216 3292
rect 20240 3290 20296 3292
rect 20000 3238 20046 3290
rect 20046 3238 20056 3290
rect 20080 3238 20110 3290
rect 20110 3238 20122 3290
rect 20122 3238 20136 3290
rect 20160 3238 20174 3290
rect 20174 3238 20186 3290
rect 20186 3238 20216 3290
rect 20240 3238 20250 3290
rect 20250 3238 20296 3290
rect 20000 3236 20056 3238
rect 20080 3236 20136 3238
rect 20160 3236 20216 3238
rect 20240 3236 20296 3238
rect 23174 9274 23230 9276
rect 23254 9274 23310 9276
rect 23334 9274 23390 9276
rect 23414 9274 23470 9276
rect 23174 9222 23220 9274
rect 23220 9222 23230 9274
rect 23254 9222 23284 9274
rect 23284 9222 23296 9274
rect 23296 9222 23310 9274
rect 23334 9222 23348 9274
rect 23348 9222 23360 9274
rect 23360 9222 23390 9274
rect 23414 9222 23424 9274
rect 23424 9222 23470 9274
rect 23174 9220 23230 9222
rect 23254 9220 23310 9222
rect 23334 9220 23390 9222
rect 23414 9220 23470 9222
rect 23570 8472 23626 8528
rect 23174 8186 23230 8188
rect 23254 8186 23310 8188
rect 23334 8186 23390 8188
rect 23414 8186 23470 8188
rect 23174 8134 23220 8186
rect 23220 8134 23230 8186
rect 23254 8134 23284 8186
rect 23284 8134 23296 8186
rect 23296 8134 23310 8186
rect 23334 8134 23348 8186
rect 23348 8134 23360 8186
rect 23360 8134 23390 8186
rect 23414 8134 23424 8186
rect 23424 8134 23470 8186
rect 23174 8132 23230 8134
rect 23254 8132 23310 8134
rect 23334 8132 23390 8134
rect 23414 8132 23470 8134
rect 23174 7098 23230 7100
rect 23254 7098 23310 7100
rect 23334 7098 23390 7100
rect 23414 7098 23470 7100
rect 23174 7046 23220 7098
rect 23220 7046 23230 7098
rect 23254 7046 23284 7098
rect 23284 7046 23296 7098
rect 23296 7046 23310 7098
rect 23334 7046 23348 7098
rect 23348 7046 23360 7098
rect 23360 7046 23390 7098
rect 23414 7046 23424 7098
rect 23424 7046 23470 7098
rect 23174 7044 23230 7046
rect 23254 7044 23310 7046
rect 23334 7044 23390 7046
rect 23414 7044 23470 7046
rect 26348 9818 26404 9820
rect 26428 9818 26484 9820
rect 26508 9818 26564 9820
rect 26588 9818 26644 9820
rect 26348 9766 26394 9818
rect 26394 9766 26404 9818
rect 26428 9766 26458 9818
rect 26458 9766 26470 9818
rect 26470 9766 26484 9818
rect 26508 9766 26522 9818
rect 26522 9766 26534 9818
rect 26534 9766 26564 9818
rect 26588 9766 26598 9818
rect 26598 9766 26644 9818
rect 26348 9764 26404 9766
rect 26428 9764 26484 9766
rect 26508 9764 26564 9766
rect 26588 9764 26644 9766
rect 24858 8472 24914 8528
rect 23174 6010 23230 6012
rect 23254 6010 23310 6012
rect 23334 6010 23390 6012
rect 23414 6010 23470 6012
rect 23174 5958 23220 6010
rect 23220 5958 23230 6010
rect 23254 5958 23284 6010
rect 23284 5958 23296 6010
rect 23296 5958 23310 6010
rect 23334 5958 23348 6010
rect 23348 5958 23360 6010
rect 23360 5958 23390 6010
rect 23414 5958 23424 6010
rect 23424 5958 23470 6010
rect 23174 5956 23230 5958
rect 23254 5956 23310 5958
rect 23334 5956 23390 5958
rect 23414 5956 23470 5958
rect 23174 4922 23230 4924
rect 23254 4922 23310 4924
rect 23334 4922 23390 4924
rect 23414 4922 23470 4924
rect 23174 4870 23220 4922
rect 23220 4870 23230 4922
rect 23254 4870 23284 4922
rect 23284 4870 23296 4922
rect 23296 4870 23310 4922
rect 23334 4870 23348 4922
rect 23348 4870 23360 4922
rect 23360 4870 23390 4922
rect 23414 4870 23424 4922
rect 23424 4870 23470 4922
rect 23174 4868 23230 4870
rect 23254 4868 23310 4870
rect 23334 4868 23390 4870
rect 23414 4868 23470 4870
rect 26348 8730 26404 8732
rect 26428 8730 26484 8732
rect 26508 8730 26564 8732
rect 26588 8730 26644 8732
rect 26348 8678 26394 8730
rect 26394 8678 26404 8730
rect 26428 8678 26458 8730
rect 26458 8678 26470 8730
rect 26470 8678 26484 8730
rect 26508 8678 26522 8730
rect 26522 8678 26534 8730
rect 26534 8678 26564 8730
rect 26588 8678 26598 8730
rect 26598 8678 26644 8730
rect 26348 8676 26404 8678
rect 26428 8676 26484 8678
rect 26508 8676 26564 8678
rect 26588 8676 26644 8678
rect 23174 3834 23230 3836
rect 23254 3834 23310 3836
rect 23334 3834 23390 3836
rect 23414 3834 23470 3836
rect 23174 3782 23220 3834
rect 23220 3782 23230 3834
rect 23254 3782 23284 3834
rect 23284 3782 23296 3834
rect 23296 3782 23310 3834
rect 23334 3782 23348 3834
rect 23348 3782 23360 3834
rect 23360 3782 23390 3834
rect 23414 3782 23424 3834
rect 23424 3782 23470 3834
rect 23174 3780 23230 3782
rect 23254 3780 23310 3782
rect 23334 3780 23390 3782
rect 23414 3780 23470 3782
rect 23174 2746 23230 2748
rect 23254 2746 23310 2748
rect 23334 2746 23390 2748
rect 23414 2746 23470 2748
rect 23174 2694 23220 2746
rect 23220 2694 23230 2746
rect 23254 2694 23284 2746
rect 23284 2694 23296 2746
rect 23296 2694 23310 2746
rect 23334 2694 23348 2746
rect 23348 2694 23360 2746
rect 23360 2694 23390 2746
rect 23414 2694 23424 2746
rect 23424 2694 23470 2746
rect 23174 2692 23230 2694
rect 23254 2692 23310 2694
rect 23334 2692 23390 2694
rect 23414 2692 23470 2694
rect 26348 7642 26404 7644
rect 26428 7642 26484 7644
rect 26508 7642 26564 7644
rect 26588 7642 26644 7644
rect 26348 7590 26394 7642
rect 26394 7590 26404 7642
rect 26428 7590 26458 7642
rect 26458 7590 26470 7642
rect 26470 7590 26484 7642
rect 26508 7590 26522 7642
rect 26522 7590 26534 7642
rect 26534 7590 26564 7642
rect 26588 7590 26598 7642
rect 26598 7590 26644 7642
rect 26348 7588 26404 7590
rect 26428 7588 26484 7590
rect 26508 7588 26564 7590
rect 26588 7588 26644 7590
rect 26348 6554 26404 6556
rect 26428 6554 26484 6556
rect 26508 6554 26564 6556
rect 26588 6554 26644 6556
rect 26348 6502 26394 6554
rect 26394 6502 26404 6554
rect 26428 6502 26458 6554
rect 26458 6502 26470 6554
rect 26470 6502 26484 6554
rect 26508 6502 26522 6554
rect 26522 6502 26534 6554
rect 26534 6502 26564 6554
rect 26588 6502 26598 6554
rect 26598 6502 26644 6554
rect 26348 6500 26404 6502
rect 26428 6500 26484 6502
rect 26508 6500 26564 6502
rect 26588 6500 26644 6502
rect 26348 5466 26404 5468
rect 26428 5466 26484 5468
rect 26508 5466 26564 5468
rect 26588 5466 26644 5468
rect 26348 5414 26394 5466
rect 26394 5414 26404 5466
rect 26428 5414 26458 5466
rect 26458 5414 26470 5466
rect 26470 5414 26484 5466
rect 26508 5414 26522 5466
rect 26522 5414 26534 5466
rect 26534 5414 26564 5466
rect 26588 5414 26598 5466
rect 26598 5414 26644 5466
rect 26348 5412 26404 5414
rect 26428 5412 26484 5414
rect 26508 5412 26564 5414
rect 26588 5412 26644 5414
rect 26514 4800 26570 4856
rect 26348 4378 26404 4380
rect 26428 4378 26484 4380
rect 26508 4378 26564 4380
rect 26588 4378 26644 4380
rect 26348 4326 26394 4378
rect 26394 4326 26404 4378
rect 26428 4326 26458 4378
rect 26458 4326 26470 4378
rect 26470 4326 26484 4378
rect 26508 4326 26522 4378
rect 26522 4326 26534 4378
rect 26534 4326 26564 4378
rect 26588 4326 26598 4378
rect 26598 4326 26644 4378
rect 26348 4324 26404 4326
rect 26428 4324 26484 4326
rect 26508 4324 26564 4326
rect 26588 4324 26644 4326
rect 26348 3290 26404 3292
rect 26428 3290 26484 3292
rect 26508 3290 26564 3292
rect 26588 3290 26644 3292
rect 26348 3238 26394 3290
rect 26394 3238 26404 3290
rect 26428 3238 26458 3290
rect 26458 3238 26470 3290
rect 26470 3238 26484 3290
rect 26508 3238 26522 3290
rect 26522 3238 26534 3290
rect 26534 3238 26564 3290
rect 26588 3238 26598 3290
rect 26598 3238 26644 3290
rect 26348 3236 26404 3238
rect 26428 3236 26484 3238
rect 26508 3236 26564 3238
rect 26588 3236 26644 3238
rect 13652 2202 13708 2204
rect 13732 2202 13788 2204
rect 13812 2202 13868 2204
rect 13892 2202 13948 2204
rect 13652 2150 13698 2202
rect 13698 2150 13708 2202
rect 13732 2150 13762 2202
rect 13762 2150 13774 2202
rect 13774 2150 13788 2202
rect 13812 2150 13826 2202
rect 13826 2150 13838 2202
rect 13838 2150 13868 2202
rect 13892 2150 13902 2202
rect 13902 2150 13948 2202
rect 13652 2148 13708 2150
rect 13732 2148 13788 2150
rect 13812 2148 13868 2150
rect 13892 2148 13948 2150
rect 20000 2202 20056 2204
rect 20080 2202 20136 2204
rect 20160 2202 20216 2204
rect 20240 2202 20296 2204
rect 20000 2150 20046 2202
rect 20046 2150 20056 2202
rect 20080 2150 20110 2202
rect 20110 2150 20122 2202
rect 20122 2150 20136 2202
rect 20160 2150 20174 2202
rect 20174 2150 20186 2202
rect 20186 2150 20216 2202
rect 20240 2150 20250 2202
rect 20250 2150 20296 2202
rect 20000 2148 20056 2150
rect 20080 2148 20136 2150
rect 20160 2148 20216 2150
rect 20240 2148 20296 2150
rect 26348 2202 26404 2204
rect 26428 2202 26484 2204
rect 26508 2202 26564 2204
rect 26588 2202 26644 2204
rect 26348 2150 26394 2202
rect 26394 2150 26404 2202
rect 26428 2150 26458 2202
rect 26458 2150 26470 2202
rect 26470 2150 26484 2202
rect 26508 2150 26522 2202
rect 26522 2150 26534 2202
rect 26534 2150 26564 2202
rect 26588 2150 26598 2202
rect 26598 2150 26644 2202
rect 26348 2148 26404 2150
rect 26428 2148 26484 2150
rect 26508 2148 26564 2150
rect 26588 2148 26644 2150
rect 26146 720 26202 776
<< metal3 >>
rect 26841 27888 27641 28008
rect 7294 27232 7610 27233
rect 7294 27168 7300 27232
rect 7364 27168 7380 27232
rect 7444 27168 7460 27232
rect 7524 27168 7540 27232
rect 7604 27168 7610 27232
rect 7294 27167 7610 27168
rect 13642 27232 13958 27233
rect 13642 27168 13648 27232
rect 13712 27168 13728 27232
rect 13792 27168 13808 27232
rect 13872 27168 13888 27232
rect 13952 27168 13958 27232
rect 13642 27167 13958 27168
rect 19990 27232 20306 27233
rect 19990 27168 19996 27232
rect 20060 27168 20076 27232
rect 20140 27168 20156 27232
rect 20220 27168 20236 27232
rect 20300 27168 20306 27232
rect 19990 27167 20306 27168
rect 26338 27232 26654 27233
rect 26338 27168 26344 27232
rect 26408 27168 26424 27232
rect 26488 27168 26504 27232
rect 26568 27168 26584 27232
rect 26648 27168 26654 27232
rect 26338 27167 26654 27168
rect 4120 26688 4436 26689
rect 0 26618 800 26648
rect 4120 26624 4126 26688
rect 4190 26624 4206 26688
rect 4270 26624 4286 26688
rect 4350 26624 4366 26688
rect 4430 26624 4436 26688
rect 4120 26623 4436 26624
rect 10468 26688 10784 26689
rect 10468 26624 10474 26688
rect 10538 26624 10554 26688
rect 10618 26624 10634 26688
rect 10698 26624 10714 26688
rect 10778 26624 10784 26688
rect 10468 26623 10784 26624
rect 16816 26688 17132 26689
rect 16816 26624 16822 26688
rect 16886 26624 16902 26688
rect 16966 26624 16982 26688
rect 17046 26624 17062 26688
rect 17126 26624 17132 26688
rect 16816 26623 17132 26624
rect 23164 26688 23480 26689
rect 23164 26624 23170 26688
rect 23234 26624 23250 26688
rect 23314 26624 23330 26688
rect 23394 26624 23410 26688
rect 23474 26624 23480 26688
rect 23164 26623 23480 26624
rect 933 26618 999 26621
rect 0 26616 999 26618
rect 0 26560 938 26616
rect 994 26560 999 26616
rect 0 26558 999 26560
rect 0 26528 800 26558
rect 933 26555 999 26558
rect 7294 26144 7610 26145
rect 7294 26080 7300 26144
rect 7364 26080 7380 26144
rect 7444 26080 7460 26144
rect 7524 26080 7540 26144
rect 7604 26080 7610 26144
rect 7294 26079 7610 26080
rect 13642 26144 13958 26145
rect 13642 26080 13648 26144
rect 13712 26080 13728 26144
rect 13792 26080 13808 26144
rect 13872 26080 13888 26144
rect 13952 26080 13958 26144
rect 13642 26079 13958 26080
rect 19990 26144 20306 26145
rect 19990 26080 19996 26144
rect 20060 26080 20076 26144
rect 20140 26080 20156 26144
rect 20220 26080 20236 26144
rect 20300 26080 20306 26144
rect 19990 26079 20306 26080
rect 26338 26144 26654 26145
rect 26338 26080 26344 26144
rect 26408 26080 26424 26144
rect 26488 26080 26504 26144
rect 26568 26080 26584 26144
rect 26648 26080 26654 26144
rect 26338 26079 26654 26080
rect 12433 25938 12499 25941
rect 13629 25938 13695 25941
rect 12433 25936 13695 25938
rect 12433 25880 12438 25936
rect 12494 25880 13634 25936
rect 13690 25880 13695 25936
rect 12433 25878 13695 25880
rect 12433 25875 12499 25878
rect 13629 25875 13695 25878
rect 12249 25802 12315 25805
rect 14457 25802 14523 25805
rect 12249 25800 14523 25802
rect 12249 25744 12254 25800
rect 12310 25744 14462 25800
rect 14518 25744 14523 25800
rect 12249 25742 14523 25744
rect 12249 25739 12315 25742
rect 14457 25739 14523 25742
rect 4120 25600 4436 25601
rect 4120 25536 4126 25600
rect 4190 25536 4206 25600
rect 4270 25536 4286 25600
rect 4350 25536 4366 25600
rect 4430 25536 4436 25600
rect 4120 25535 4436 25536
rect 10468 25600 10784 25601
rect 10468 25536 10474 25600
rect 10538 25536 10554 25600
rect 10618 25536 10634 25600
rect 10698 25536 10714 25600
rect 10778 25536 10784 25600
rect 10468 25535 10784 25536
rect 16816 25600 17132 25601
rect 16816 25536 16822 25600
rect 16886 25536 16902 25600
rect 16966 25536 16982 25600
rect 17046 25536 17062 25600
rect 17126 25536 17132 25600
rect 16816 25535 17132 25536
rect 23164 25600 23480 25601
rect 23164 25536 23170 25600
rect 23234 25536 23250 25600
rect 23314 25536 23330 25600
rect 23394 25536 23410 25600
rect 23474 25536 23480 25600
rect 23164 25535 23480 25536
rect 7294 25056 7610 25057
rect 7294 24992 7300 25056
rect 7364 24992 7380 25056
rect 7444 24992 7460 25056
rect 7524 24992 7540 25056
rect 7604 24992 7610 25056
rect 7294 24991 7610 24992
rect 13642 25056 13958 25057
rect 13642 24992 13648 25056
rect 13712 24992 13728 25056
rect 13792 24992 13808 25056
rect 13872 24992 13888 25056
rect 13952 24992 13958 25056
rect 13642 24991 13958 24992
rect 19990 25056 20306 25057
rect 19990 24992 19996 25056
rect 20060 24992 20076 25056
rect 20140 24992 20156 25056
rect 20220 24992 20236 25056
rect 20300 24992 20306 25056
rect 19990 24991 20306 24992
rect 26338 25056 26654 25057
rect 26338 24992 26344 25056
rect 26408 24992 26424 25056
rect 26488 24992 26504 25056
rect 26568 24992 26584 25056
rect 26648 24992 26654 25056
rect 26338 24991 26654 24992
rect 4120 24512 4436 24513
rect 4120 24448 4126 24512
rect 4190 24448 4206 24512
rect 4270 24448 4286 24512
rect 4350 24448 4366 24512
rect 4430 24448 4436 24512
rect 4120 24447 4436 24448
rect 10468 24512 10784 24513
rect 10468 24448 10474 24512
rect 10538 24448 10554 24512
rect 10618 24448 10634 24512
rect 10698 24448 10714 24512
rect 10778 24448 10784 24512
rect 10468 24447 10784 24448
rect 16816 24512 17132 24513
rect 16816 24448 16822 24512
rect 16886 24448 16902 24512
rect 16966 24448 16982 24512
rect 17046 24448 17062 24512
rect 17126 24448 17132 24512
rect 16816 24447 17132 24448
rect 23164 24512 23480 24513
rect 23164 24448 23170 24512
rect 23234 24448 23250 24512
rect 23314 24448 23330 24512
rect 23394 24448 23410 24512
rect 23474 24448 23480 24512
rect 23164 24447 23480 24448
rect 7294 23968 7610 23969
rect 7294 23904 7300 23968
rect 7364 23904 7380 23968
rect 7444 23904 7460 23968
rect 7524 23904 7540 23968
rect 7604 23904 7610 23968
rect 7294 23903 7610 23904
rect 13642 23968 13958 23969
rect 13642 23904 13648 23968
rect 13712 23904 13728 23968
rect 13792 23904 13808 23968
rect 13872 23904 13888 23968
rect 13952 23904 13958 23968
rect 13642 23903 13958 23904
rect 19990 23968 20306 23969
rect 19990 23904 19996 23968
rect 20060 23904 20076 23968
rect 20140 23904 20156 23968
rect 20220 23904 20236 23968
rect 20300 23904 20306 23968
rect 19990 23903 20306 23904
rect 26338 23968 26654 23969
rect 26338 23904 26344 23968
rect 26408 23904 26424 23968
rect 26488 23904 26504 23968
rect 26568 23904 26584 23968
rect 26648 23904 26654 23968
rect 26338 23903 26654 23904
rect 26841 23864 27641 23928
rect 26742 23808 27641 23864
rect 26742 23804 26986 23808
rect 26141 23762 26207 23765
rect 26742 23762 26802 23804
rect 26141 23760 26802 23762
rect 26141 23704 26146 23760
rect 26202 23704 26802 23760
rect 26141 23702 26802 23704
rect 26141 23699 26207 23702
rect 4120 23424 4436 23425
rect 4120 23360 4126 23424
rect 4190 23360 4206 23424
rect 4270 23360 4286 23424
rect 4350 23360 4366 23424
rect 4430 23360 4436 23424
rect 4120 23359 4436 23360
rect 10468 23424 10784 23425
rect 10468 23360 10474 23424
rect 10538 23360 10554 23424
rect 10618 23360 10634 23424
rect 10698 23360 10714 23424
rect 10778 23360 10784 23424
rect 10468 23359 10784 23360
rect 16816 23424 17132 23425
rect 16816 23360 16822 23424
rect 16886 23360 16902 23424
rect 16966 23360 16982 23424
rect 17046 23360 17062 23424
rect 17126 23360 17132 23424
rect 16816 23359 17132 23360
rect 23164 23424 23480 23425
rect 23164 23360 23170 23424
rect 23234 23360 23250 23424
rect 23314 23360 23330 23424
rect 23394 23360 23410 23424
rect 23474 23360 23480 23424
rect 23164 23359 23480 23360
rect 7294 22880 7610 22881
rect 7294 22816 7300 22880
rect 7364 22816 7380 22880
rect 7444 22816 7460 22880
rect 7524 22816 7540 22880
rect 7604 22816 7610 22880
rect 7294 22815 7610 22816
rect 13642 22880 13958 22881
rect 13642 22816 13648 22880
rect 13712 22816 13728 22880
rect 13792 22816 13808 22880
rect 13872 22816 13888 22880
rect 13952 22816 13958 22880
rect 13642 22815 13958 22816
rect 19990 22880 20306 22881
rect 19990 22816 19996 22880
rect 20060 22816 20076 22880
rect 20140 22816 20156 22880
rect 20220 22816 20236 22880
rect 20300 22816 20306 22880
rect 19990 22815 20306 22816
rect 26338 22880 26654 22881
rect 26338 22816 26344 22880
rect 26408 22816 26424 22880
rect 26488 22816 26504 22880
rect 26568 22816 26584 22880
rect 26648 22816 26654 22880
rect 26338 22815 26654 22816
rect 22277 22674 22343 22677
rect 23105 22674 23171 22677
rect 22277 22672 23171 22674
rect 22277 22616 22282 22672
rect 22338 22616 23110 22672
rect 23166 22616 23171 22672
rect 22277 22614 23171 22616
rect 22277 22611 22343 22614
rect 23105 22611 23171 22614
rect 0 22448 800 22568
rect 4120 22336 4436 22337
rect 4120 22272 4126 22336
rect 4190 22272 4206 22336
rect 4270 22272 4286 22336
rect 4350 22272 4366 22336
rect 4430 22272 4436 22336
rect 4120 22271 4436 22272
rect 10468 22336 10784 22337
rect 10468 22272 10474 22336
rect 10538 22272 10554 22336
rect 10618 22272 10634 22336
rect 10698 22272 10714 22336
rect 10778 22272 10784 22336
rect 10468 22271 10784 22272
rect 16816 22336 17132 22337
rect 16816 22272 16822 22336
rect 16886 22272 16902 22336
rect 16966 22272 16982 22336
rect 17046 22272 17062 22336
rect 17126 22272 17132 22336
rect 16816 22271 17132 22272
rect 23164 22336 23480 22337
rect 23164 22272 23170 22336
rect 23234 22272 23250 22336
rect 23314 22272 23330 22336
rect 23394 22272 23410 22336
rect 23474 22272 23480 22336
rect 23164 22271 23480 22272
rect 7294 21792 7610 21793
rect 7294 21728 7300 21792
rect 7364 21728 7380 21792
rect 7444 21728 7460 21792
rect 7524 21728 7540 21792
rect 7604 21728 7610 21792
rect 7294 21727 7610 21728
rect 13642 21792 13958 21793
rect 13642 21728 13648 21792
rect 13712 21728 13728 21792
rect 13792 21728 13808 21792
rect 13872 21728 13888 21792
rect 13952 21728 13958 21792
rect 13642 21727 13958 21728
rect 19990 21792 20306 21793
rect 19990 21728 19996 21792
rect 20060 21728 20076 21792
rect 20140 21728 20156 21792
rect 20220 21728 20236 21792
rect 20300 21728 20306 21792
rect 19990 21727 20306 21728
rect 26338 21792 26654 21793
rect 26338 21728 26344 21792
rect 26408 21728 26424 21792
rect 26488 21728 26504 21792
rect 26568 21728 26584 21792
rect 26648 21728 26654 21792
rect 26338 21727 26654 21728
rect 16757 21586 16823 21589
rect 17677 21586 17743 21589
rect 18321 21586 18387 21589
rect 16757 21584 18387 21586
rect 16757 21528 16762 21584
rect 16818 21528 17682 21584
rect 17738 21528 18326 21584
rect 18382 21528 18387 21584
rect 16757 21526 18387 21528
rect 16757 21523 16823 21526
rect 17677 21523 17743 21526
rect 18321 21523 18387 21526
rect 17217 21450 17283 21453
rect 18597 21450 18663 21453
rect 17217 21448 18663 21450
rect 17217 21392 17222 21448
rect 17278 21392 18602 21448
rect 18658 21392 18663 21448
rect 17217 21390 18663 21392
rect 17217 21387 17283 21390
rect 18597 21387 18663 21390
rect 4120 21248 4436 21249
rect 4120 21184 4126 21248
rect 4190 21184 4206 21248
rect 4270 21184 4286 21248
rect 4350 21184 4366 21248
rect 4430 21184 4436 21248
rect 4120 21183 4436 21184
rect 10468 21248 10784 21249
rect 10468 21184 10474 21248
rect 10538 21184 10554 21248
rect 10618 21184 10634 21248
rect 10698 21184 10714 21248
rect 10778 21184 10784 21248
rect 10468 21183 10784 21184
rect 16816 21248 17132 21249
rect 16816 21184 16822 21248
rect 16886 21184 16902 21248
rect 16966 21184 16982 21248
rect 17046 21184 17062 21248
rect 17126 21184 17132 21248
rect 16816 21183 17132 21184
rect 23164 21248 23480 21249
rect 23164 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23480 21248
rect 23164 21183 23480 21184
rect 7294 20704 7610 20705
rect 7294 20640 7300 20704
rect 7364 20640 7380 20704
rect 7444 20640 7460 20704
rect 7524 20640 7540 20704
rect 7604 20640 7610 20704
rect 7294 20639 7610 20640
rect 13642 20704 13958 20705
rect 13642 20640 13648 20704
rect 13712 20640 13728 20704
rect 13792 20640 13808 20704
rect 13872 20640 13888 20704
rect 13952 20640 13958 20704
rect 13642 20639 13958 20640
rect 19990 20704 20306 20705
rect 19990 20640 19996 20704
rect 20060 20640 20076 20704
rect 20140 20640 20156 20704
rect 20220 20640 20236 20704
rect 20300 20640 20306 20704
rect 19990 20639 20306 20640
rect 26338 20704 26654 20705
rect 26338 20640 26344 20704
rect 26408 20640 26424 20704
rect 26488 20640 26504 20704
rect 26568 20640 26584 20704
rect 26648 20640 26654 20704
rect 26338 20639 26654 20640
rect 16941 20634 17007 20637
rect 18505 20634 18571 20637
rect 16941 20632 18571 20634
rect 16941 20576 16946 20632
rect 17002 20576 18510 20632
rect 18566 20576 18571 20632
rect 16941 20574 18571 20576
rect 16941 20571 17007 20574
rect 18505 20571 18571 20574
rect 8569 20498 8635 20501
rect 11605 20498 11671 20501
rect 8569 20496 11671 20498
rect 8569 20440 8574 20496
rect 8630 20440 11610 20496
rect 11666 20440 11671 20496
rect 8569 20438 11671 20440
rect 8569 20435 8635 20438
rect 11605 20435 11671 20438
rect 4120 20160 4436 20161
rect 4120 20096 4126 20160
rect 4190 20096 4206 20160
rect 4270 20096 4286 20160
rect 4350 20096 4366 20160
rect 4430 20096 4436 20160
rect 4120 20095 4436 20096
rect 10468 20160 10784 20161
rect 10468 20096 10474 20160
rect 10538 20096 10554 20160
rect 10618 20096 10634 20160
rect 10698 20096 10714 20160
rect 10778 20096 10784 20160
rect 10468 20095 10784 20096
rect 16816 20160 17132 20161
rect 16816 20096 16822 20160
rect 16886 20096 16902 20160
rect 16966 20096 16982 20160
rect 17046 20096 17062 20160
rect 17126 20096 17132 20160
rect 16816 20095 17132 20096
rect 23164 20160 23480 20161
rect 23164 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23480 20160
rect 23164 20095 23480 20096
rect 26841 19728 27641 19848
rect 7294 19616 7610 19617
rect 7294 19552 7300 19616
rect 7364 19552 7380 19616
rect 7444 19552 7460 19616
rect 7524 19552 7540 19616
rect 7604 19552 7610 19616
rect 7294 19551 7610 19552
rect 13642 19616 13958 19617
rect 13642 19552 13648 19616
rect 13712 19552 13728 19616
rect 13792 19552 13808 19616
rect 13872 19552 13888 19616
rect 13952 19552 13958 19616
rect 13642 19551 13958 19552
rect 19990 19616 20306 19617
rect 19990 19552 19996 19616
rect 20060 19552 20076 19616
rect 20140 19552 20156 19616
rect 20220 19552 20236 19616
rect 20300 19552 20306 19616
rect 19990 19551 20306 19552
rect 26338 19616 26654 19617
rect 26338 19552 26344 19616
rect 26408 19552 26424 19616
rect 26488 19552 26504 19616
rect 26568 19552 26584 19616
rect 26648 19552 26654 19616
rect 26338 19551 26654 19552
rect 10409 19274 10475 19277
rect 12617 19274 12683 19277
rect 10409 19272 12683 19274
rect 10409 19216 10414 19272
rect 10470 19216 12622 19272
rect 12678 19216 12683 19272
rect 10409 19214 12683 19216
rect 10409 19211 10475 19214
rect 12617 19211 12683 19214
rect 0 19138 800 19168
rect 933 19138 999 19141
rect 0 19136 999 19138
rect 0 19080 938 19136
rect 994 19080 999 19136
rect 0 19078 999 19080
rect 0 19048 800 19078
rect 933 19075 999 19078
rect 4120 19072 4436 19073
rect 4120 19008 4126 19072
rect 4190 19008 4206 19072
rect 4270 19008 4286 19072
rect 4350 19008 4366 19072
rect 4430 19008 4436 19072
rect 4120 19007 4436 19008
rect 10468 19072 10784 19073
rect 10468 19008 10474 19072
rect 10538 19008 10554 19072
rect 10618 19008 10634 19072
rect 10698 19008 10714 19072
rect 10778 19008 10784 19072
rect 10468 19007 10784 19008
rect 16816 19072 17132 19073
rect 16816 19008 16822 19072
rect 16886 19008 16902 19072
rect 16966 19008 16982 19072
rect 17046 19008 17062 19072
rect 17126 19008 17132 19072
rect 16816 19007 17132 19008
rect 23164 19072 23480 19073
rect 23164 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23480 19072
rect 23164 19007 23480 19008
rect 7294 18528 7610 18529
rect 7294 18464 7300 18528
rect 7364 18464 7380 18528
rect 7444 18464 7460 18528
rect 7524 18464 7540 18528
rect 7604 18464 7610 18528
rect 7294 18463 7610 18464
rect 13642 18528 13958 18529
rect 13642 18464 13648 18528
rect 13712 18464 13728 18528
rect 13792 18464 13808 18528
rect 13872 18464 13888 18528
rect 13952 18464 13958 18528
rect 13642 18463 13958 18464
rect 19990 18528 20306 18529
rect 19990 18464 19996 18528
rect 20060 18464 20076 18528
rect 20140 18464 20156 18528
rect 20220 18464 20236 18528
rect 20300 18464 20306 18528
rect 19990 18463 20306 18464
rect 26338 18528 26654 18529
rect 26338 18464 26344 18528
rect 26408 18464 26424 18528
rect 26488 18464 26504 18528
rect 26568 18464 26584 18528
rect 26648 18464 26654 18528
rect 26338 18463 26654 18464
rect 4120 17984 4436 17985
rect 4120 17920 4126 17984
rect 4190 17920 4206 17984
rect 4270 17920 4286 17984
rect 4350 17920 4366 17984
rect 4430 17920 4436 17984
rect 4120 17919 4436 17920
rect 10468 17984 10784 17985
rect 10468 17920 10474 17984
rect 10538 17920 10554 17984
rect 10618 17920 10634 17984
rect 10698 17920 10714 17984
rect 10778 17920 10784 17984
rect 10468 17919 10784 17920
rect 16816 17984 17132 17985
rect 16816 17920 16822 17984
rect 16886 17920 16902 17984
rect 16966 17920 16982 17984
rect 17046 17920 17062 17984
rect 17126 17920 17132 17984
rect 16816 17919 17132 17920
rect 23164 17984 23480 17985
rect 23164 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23480 17984
rect 23164 17919 23480 17920
rect 7294 17440 7610 17441
rect 7294 17376 7300 17440
rect 7364 17376 7380 17440
rect 7444 17376 7460 17440
rect 7524 17376 7540 17440
rect 7604 17376 7610 17440
rect 7294 17375 7610 17376
rect 13642 17440 13958 17441
rect 13642 17376 13648 17440
rect 13712 17376 13728 17440
rect 13792 17376 13808 17440
rect 13872 17376 13888 17440
rect 13952 17376 13958 17440
rect 13642 17375 13958 17376
rect 19990 17440 20306 17441
rect 19990 17376 19996 17440
rect 20060 17376 20076 17440
rect 20140 17376 20156 17440
rect 20220 17376 20236 17440
rect 20300 17376 20306 17440
rect 19990 17375 20306 17376
rect 26338 17440 26654 17441
rect 26338 17376 26344 17440
rect 26408 17376 26424 17440
rect 26488 17376 26504 17440
rect 26568 17376 26584 17440
rect 26648 17376 26654 17440
rect 26338 17375 26654 17376
rect 18689 17234 18755 17237
rect 19057 17234 19123 17237
rect 18689 17232 19123 17234
rect 18689 17176 18694 17232
rect 18750 17176 19062 17232
rect 19118 17176 19123 17232
rect 18689 17174 19123 17176
rect 18689 17171 18755 17174
rect 19057 17171 19123 17174
rect 21633 17234 21699 17237
rect 22645 17234 22711 17237
rect 21633 17232 22711 17234
rect 21633 17176 21638 17232
rect 21694 17176 22650 17232
rect 22706 17176 22711 17232
rect 21633 17174 22711 17176
rect 21633 17171 21699 17174
rect 22645 17171 22711 17174
rect 15745 17098 15811 17101
rect 19241 17098 19307 17101
rect 15745 17096 19307 17098
rect 15745 17040 15750 17096
rect 15806 17040 19246 17096
rect 19302 17040 19307 17096
rect 15745 17038 19307 17040
rect 15745 17035 15811 17038
rect 19241 17035 19307 17038
rect 22461 17098 22527 17101
rect 23657 17098 23723 17101
rect 22461 17096 23723 17098
rect 22461 17040 22466 17096
rect 22522 17040 23662 17096
rect 23718 17040 23723 17096
rect 22461 17038 23723 17040
rect 22461 17035 22527 17038
rect 23657 17035 23723 17038
rect 4120 16896 4436 16897
rect 4120 16832 4126 16896
rect 4190 16832 4206 16896
rect 4270 16832 4286 16896
rect 4350 16832 4366 16896
rect 4430 16832 4436 16896
rect 4120 16831 4436 16832
rect 10468 16896 10784 16897
rect 10468 16832 10474 16896
rect 10538 16832 10554 16896
rect 10618 16832 10634 16896
rect 10698 16832 10714 16896
rect 10778 16832 10784 16896
rect 10468 16831 10784 16832
rect 16816 16896 17132 16897
rect 16816 16832 16822 16896
rect 16886 16832 16902 16896
rect 16966 16832 16982 16896
rect 17046 16832 17062 16896
rect 17126 16832 17132 16896
rect 16816 16831 17132 16832
rect 23164 16896 23480 16897
rect 23164 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23480 16896
rect 23164 16831 23480 16832
rect 7294 16352 7610 16353
rect 7294 16288 7300 16352
rect 7364 16288 7380 16352
rect 7444 16288 7460 16352
rect 7524 16288 7540 16352
rect 7604 16288 7610 16352
rect 7294 16287 7610 16288
rect 13642 16352 13958 16353
rect 13642 16288 13648 16352
rect 13712 16288 13728 16352
rect 13792 16288 13808 16352
rect 13872 16288 13888 16352
rect 13952 16288 13958 16352
rect 13642 16287 13958 16288
rect 19990 16352 20306 16353
rect 19990 16288 19996 16352
rect 20060 16288 20076 16352
rect 20140 16288 20156 16352
rect 20220 16288 20236 16352
rect 20300 16288 20306 16352
rect 19990 16287 20306 16288
rect 26338 16352 26654 16353
rect 26338 16288 26344 16352
rect 26408 16288 26424 16352
rect 26488 16288 26504 16352
rect 26568 16288 26584 16352
rect 26648 16288 26654 16352
rect 26841 16328 27641 16448
rect 26338 16287 26654 16288
rect 12617 16146 12683 16149
rect 14641 16146 14707 16149
rect 16205 16146 16271 16149
rect 12617 16144 16271 16146
rect 12617 16088 12622 16144
rect 12678 16088 14646 16144
rect 14702 16088 16210 16144
rect 16266 16088 16271 16144
rect 12617 16086 16271 16088
rect 12617 16083 12683 16086
rect 14641 16083 14707 16086
rect 16205 16083 16271 16086
rect 4120 15808 4436 15809
rect 4120 15744 4126 15808
rect 4190 15744 4206 15808
rect 4270 15744 4286 15808
rect 4350 15744 4366 15808
rect 4430 15744 4436 15808
rect 4120 15743 4436 15744
rect 10468 15808 10784 15809
rect 10468 15744 10474 15808
rect 10538 15744 10554 15808
rect 10618 15744 10634 15808
rect 10698 15744 10714 15808
rect 10778 15744 10784 15808
rect 10468 15743 10784 15744
rect 16816 15808 17132 15809
rect 16816 15744 16822 15808
rect 16886 15744 16902 15808
rect 16966 15744 16982 15808
rect 17046 15744 17062 15808
rect 17126 15744 17132 15808
rect 16816 15743 17132 15744
rect 23164 15808 23480 15809
rect 23164 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23480 15808
rect 23164 15743 23480 15744
rect 7294 15264 7610 15265
rect 7294 15200 7300 15264
rect 7364 15200 7380 15264
rect 7444 15200 7460 15264
rect 7524 15200 7540 15264
rect 7604 15200 7610 15264
rect 7294 15199 7610 15200
rect 13642 15264 13958 15265
rect 13642 15200 13648 15264
rect 13712 15200 13728 15264
rect 13792 15200 13808 15264
rect 13872 15200 13888 15264
rect 13952 15200 13958 15264
rect 13642 15199 13958 15200
rect 19990 15264 20306 15265
rect 19990 15200 19996 15264
rect 20060 15200 20076 15264
rect 20140 15200 20156 15264
rect 20220 15200 20236 15264
rect 20300 15200 20306 15264
rect 19990 15199 20306 15200
rect 26338 15264 26654 15265
rect 26338 15200 26344 15264
rect 26408 15200 26424 15264
rect 26488 15200 26504 15264
rect 26568 15200 26584 15264
rect 26648 15200 26654 15264
rect 26338 15199 26654 15200
rect 1393 15194 1459 15197
rect 798 15192 1459 15194
rect 798 15136 1398 15192
rect 1454 15136 1459 15192
rect 798 15134 1459 15136
rect 798 15088 858 15134
rect 1393 15131 1459 15134
rect 0 14998 858 15088
rect 0 14968 800 14998
rect 4120 14720 4436 14721
rect 4120 14656 4126 14720
rect 4190 14656 4206 14720
rect 4270 14656 4286 14720
rect 4350 14656 4366 14720
rect 4430 14656 4436 14720
rect 4120 14655 4436 14656
rect 10468 14720 10784 14721
rect 10468 14656 10474 14720
rect 10538 14656 10554 14720
rect 10618 14656 10634 14720
rect 10698 14656 10714 14720
rect 10778 14656 10784 14720
rect 10468 14655 10784 14656
rect 16816 14720 17132 14721
rect 16816 14656 16822 14720
rect 16886 14656 16902 14720
rect 16966 14656 16982 14720
rect 17046 14656 17062 14720
rect 17126 14656 17132 14720
rect 16816 14655 17132 14656
rect 23164 14720 23480 14721
rect 23164 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23480 14720
rect 23164 14655 23480 14656
rect 7294 14176 7610 14177
rect 7294 14112 7300 14176
rect 7364 14112 7380 14176
rect 7444 14112 7460 14176
rect 7524 14112 7540 14176
rect 7604 14112 7610 14176
rect 7294 14111 7610 14112
rect 13642 14176 13958 14177
rect 13642 14112 13648 14176
rect 13712 14112 13728 14176
rect 13792 14112 13808 14176
rect 13872 14112 13888 14176
rect 13952 14112 13958 14176
rect 13642 14111 13958 14112
rect 19990 14176 20306 14177
rect 19990 14112 19996 14176
rect 20060 14112 20076 14176
rect 20140 14112 20156 14176
rect 20220 14112 20236 14176
rect 20300 14112 20306 14176
rect 19990 14111 20306 14112
rect 26338 14176 26654 14177
rect 26338 14112 26344 14176
rect 26408 14112 26424 14176
rect 26488 14112 26504 14176
rect 26568 14112 26584 14176
rect 26648 14112 26654 14176
rect 26338 14111 26654 14112
rect 4120 13632 4436 13633
rect 4120 13568 4126 13632
rect 4190 13568 4206 13632
rect 4270 13568 4286 13632
rect 4350 13568 4366 13632
rect 4430 13568 4436 13632
rect 4120 13567 4436 13568
rect 10468 13632 10784 13633
rect 10468 13568 10474 13632
rect 10538 13568 10554 13632
rect 10618 13568 10634 13632
rect 10698 13568 10714 13632
rect 10778 13568 10784 13632
rect 10468 13567 10784 13568
rect 16816 13632 17132 13633
rect 16816 13568 16822 13632
rect 16886 13568 16902 13632
rect 16966 13568 16982 13632
rect 17046 13568 17062 13632
rect 17126 13568 17132 13632
rect 16816 13567 17132 13568
rect 23164 13632 23480 13633
rect 23164 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23480 13632
rect 23164 13567 23480 13568
rect 7294 13088 7610 13089
rect 7294 13024 7300 13088
rect 7364 13024 7380 13088
rect 7444 13024 7460 13088
rect 7524 13024 7540 13088
rect 7604 13024 7610 13088
rect 7294 13023 7610 13024
rect 13642 13088 13958 13089
rect 13642 13024 13648 13088
rect 13712 13024 13728 13088
rect 13792 13024 13808 13088
rect 13872 13024 13888 13088
rect 13952 13024 13958 13088
rect 13642 13023 13958 13024
rect 19990 13088 20306 13089
rect 19990 13024 19996 13088
rect 20060 13024 20076 13088
rect 20140 13024 20156 13088
rect 20220 13024 20236 13088
rect 20300 13024 20306 13088
rect 19990 13023 20306 13024
rect 26338 13088 26654 13089
rect 26338 13024 26344 13088
rect 26408 13024 26424 13088
rect 26488 13024 26504 13088
rect 26568 13024 26584 13088
rect 26648 13024 26654 13088
rect 26338 13023 26654 13024
rect 4120 12544 4436 12545
rect 4120 12480 4126 12544
rect 4190 12480 4206 12544
rect 4270 12480 4286 12544
rect 4350 12480 4366 12544
rect 4430 12480 4436 12544
rect 4120 12479 4436 12480
rect 10468 12544 10784 12545
rect 10468 12480 10474 12544
rect 10538 12480 10554 12544
rect 10618 12480 10634 12544
rect 10698 12480 10714 12544
rect 10778 12480 10784 12544
rect 10468 12479 10784 12480
rect 16816 12544 17132 12545
rect 16816 12480 16822 12544
rect 16886 12480 16902 12544
rect 16966 12480 16982 12544
rect 17046 12480 17062 12544
rect 17126 12480 17132 12544
rect 16816 12479 17132 12480
rect 23164 12544 23480 12545
rect 23164 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23480 12544
rect 23164 12479 23480 12480
rect 26141 12338 26207 12341
rect 26841 12338 27641 12368
rect 26141 12336 27641 12338
rect 26141 12280 26146 12336
rect 26202 12280 27641 12336
rect 26141 12278 27641 12280
rect 26141 12275 26207 12278
rect 26841 12248 27641 12278
rect 7294 12000 7610 12001
rect 7294 11936 7300 12000
rect 7364 11936 7380 12000
rect 7444 11936 7460 12000
rect 7524 11936 7540 12000
rect 7604 11936 7610 12000
rect 7294 11935 7610 11936
rect 13642 12000 13958 12001
rect 13642 11936 13648 12000
rect 13712 11936 13728 12000
rect 13792 11936 13808 12000
rect 13872 11936 13888 12000
rect 13952 11936 13958 12000
rect 13642 11935 13958 11936
rect 19990 12000 20306 12001
rect 19990 11936 19996 12000
rect 20060 11936 20076 12000
rect 20140 11936 20156 12000
rect 20220 11936 20236 12000
rect 20300 11936 20306 12000
rect 19990 11935 20306 11936
rect 26338 12000 26654 12001
rect 26338 11936 26344 12000
rect 26408 11936 26424 12000
rect 26488 11936 26504 12000
rect 26568 11936 26584 12000
rect 26648 11936 26654 12000
rect 26338 11935 26654 11936
rect 15101 11794 15167 11797
rect 17953 11794 18019 11797
rect 15101 11792 18019 11794
rect 15101 11736 15106 11792
rect 15162 11736 17958 11792
rect 18014 11736 18019 11792
rect 15101 11734 18019 11736
rect 15101 11731 15167 11734
rect 17953 11731 18019 11734
rect 4120 11456 4436 11457
rect 4120 11392 4126 11456
rect 4190 11392 4206 11456
rect 4270 11392 4286 11456
rect 4350 11392 4366 11456
rect 4430 11392 4436 11456
rect 4120 11391 4436 11392
rect 10468 11456 10784 11457
rect 10468 11392 10474 11456
rect 10538 11392 10554 11456
rect 10618 11392 10634 11456
rect 10698 11392 10714 11456
rect 10778 11392 10784 11456
rect 10468 11391 10784 11392
rect 16816 11456 17132 11457
rect 16816 11392 16822 11456
rect 16886 11392 16902 11456
rect 16966 11392 16982 11456
rect 17046 11392 17062 11456
rect 17126 11392 17132 11456
rect 16816 11391 17132 11392
rect 23164 11456 23480 11457
rect 23164 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23480 11456
rect 23164 11391 23480 11392
rect 14181 11250 14247 11253
rect 15837 11250 15903 11253
rect 14181 11248 15903 11250
rect 14181 11192 14186 11248
rect 14242 11192 15842 11248
rect 15898 11192 15903 11248
rect 14181 11190 15903 11192
rect 14181 11187 14247 11190
rect 15837 11187 15903 11190
rect 14549 11114 14615 11117
rect 19333 11114 19399 11117
rect 14549 11112 19399 11114
rect 14549 11056 14554 11112
rect 14610 11056 19338 11112
rect 19394 11056 19399 11112
rect 14549 11054 19399 11056
rect 14549 11051 14615 11054
rect 19333 11051 19399 11054
rect 0 10888 800 11008
rect 7294 10912 7610 10913
rect 7294 10848 7300 10912
rect 7364 10848 7380 10912
rect 7444 10848 7460 10912
rect 7524 10848 7540 10912
rect 7604 10848 7610 10912
rect 7294 10847 7610 10848
rect 13642 10912 13958 10913
rect 13642 10848 13648 10912
rect 13712 10848 13728 10912
rect 13792 10848 13808 10912
rect 13872 10848 13888 10912
rect 13952 10848 13958 10912
rect 13642 10847 13958 10848
rect 19990 10912 20306 10913
rect 19990 10848 19996 10912
rect 20060 10848 20076 10912
rect 20140 10848 20156 10912
rect 20220 10848 20236 10912
rect 20300 10848 20306 10912
rect 19990 10847 20306 10848
rect 26338 10912 26654 10913
rect 26338 10848 26344 10912
rect 26408 10848 26424 10912
rect 26488 10848 26504 10912
rect 26568 10848 26584 10912
rect 26648 10848 26654 10912
rect 26338 10847 26654 10848
rect 4120 10368 4436 10369
rect 4120 10304 4126 10368
rect 4190 10304 4206 10368
rect 4270 10304 4286 10368
rect 4350 10304 4366 10368
rect 4430 10304 4436 10368
rect 4120 10303 4436 10304
rect 10468 10368 10784 10369
rect 10468 10304 10474 10368
rect 10538 10304 10554 10368
rect 10618 10304 10634 10368
rect 10698 10304 10714 10368
rect 10778 10304 10784 10368
rect 10468 10303 10784 10304
rect 16816 10368 17132 10369
rect 16816 10304 16822 10368
rect 16886 10304 16902 10368
rect 16966 10304 16982 10368
rect 17046 10304 17062 10368
rect 17126 10304 17132 10368
rect 16816 10303 17132 10304
rect 23164 10368 23480 10369
rect 23164 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23480 10368
rect 23164 10303 23480 10304
rect 7294 9824 7610 9825
rect 7294 9760 7300 9824
rect 7364 9760 7380 9824
rect 7444 9760 7460 9824
rect 7524 9760 7540 9824
rect 7604 9760 7610 9824
rect 7294 9759 7610 9760
rect 13642 9824 13958 9825
rect 13642 9760 13648 9824
rect 13712 9760 13728 9824
rect 13792 9760 13808 9824
rect 13872 9760 13888 9824
rect 13952 9760 13958 9824
rect 13642 9759 13958 9760
rect 19990 9824 20306 9825
rect 19990 9760 19996 9824
rect 20060 9760 20076 9824
rect 20140 9760 20156 9824
rect 20220 9760 20236 9824
rect 20300 9760 20306 9824
rect 19990 9759 20306 9760
rect 26338 9824 26654 9825
rect 26338 9760 26344 9824
rect 26408 9760 26424 9824
rect 26488 9760 26504 9824
rect 26568 9760 26584 9824
rect 26648 9760 26654 9824
rect 26338 9759 26654 9760
rect 4120 9280 4436 9281
rect 4120 9216 4126 9280
rect 4190 9216 4206 9280
rect 4270 9216 4286 9280
rect 4350 9216 4366 9280
rect 4430 9216 4436 9280
rect 4120 9215 4436 9216
rect 10468 9280 10784 9281
rect 10468 9216 10474 9280
rect 10538 9216 10554 9280
rect 10618 9216 10634 9280
rect 10698 9216 10714 9280
rect 10778 9216 10784 9280
rect 10468 9215 10784 9216
rect 16816 9280 17132 9281
rect 16816 9216 16822 9280
rect 16886 9216 16902 9280
rect 16966 9216 16982 9280
rect 17046 9216 17062 9280
rect 17126 9216 17132 9280
rect 16816 9215 17132 9216
rect 23164 9280 23480 9281
rect 23164 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23480 9280
rect 23164 9215 23480 9216
rect 12433 9074 12499 9077
rect 13353 9074 13419 9077
rect 12433 9072 13419 9074
rect 12433 9016 12438 9072
rect 12494 9016 13358 9072
rect 13414 9016 13419 9072
rect 12433 9014 13419 9016
rect 12433 9011 12499 9014
rect 13353 9011 13419 9014
rect 26841 8848 27641 8968
rect 11145 8802 11211 8805
rect 12893 8802 12959 8805
rect 11145 8800 12959 8802
rect 11145 8744 11150 8800
rect 11206 8744 12898 8800
rect 12954 8744 12959 8800
rect 11145 8742 12959 8744
rect 11145 8739 11211 8742
rect 12893 8739 12959 8742
rect 7294 8736 7610 8737
rect 7294 8672 7300 8736
rect 7364 8672 7380 8736
rect 7444 8672 7460 8736
rect 7524 8672 7540 8736
rect 7604 8672 7610 8736
rect 7294 8671 7610 8672
rect 13642 8736 13958 8737
rect 13642 8672 13648 8736
rect 13712 8672 13728 8736
rect 13792 8672 13808 8736
rect 13872 8672 13888 8736
rect 13952 8672 13958 8736
rect 13642 8671 13958 8672
rect 19990 8736 20306 8737
rect 19990 8672 19996 8736
rect 20060 8672 20076 8736
rect 20140 8672 20156 8736
rect 20220 8672 20236 8736
rect 20300 8672 20306 8736
rect 19990 8671 20306 8672
rect 26338 8736 26654 8737
rect 26338 8672 26344 8736
rect 26408 8672 26424 8736
rect 26488 8672 26504 8736
rect 26568 8672 26584 8736
rect 26648 8672 26654 8736
rect 26338 8671 26654 8672
rect 23565 8530 23631 8533
rect 24853 8530 24919 8533
rect 23565 8528 24919 8530
rect 23565 8472 23570 8528
rect 23626 8472 24858 8528
rect 24914 8472 24919 8528
rect 23565 8470 24919 8472
rect 23565 8467 23631 8470
rect 24853 8467 24919 8470
rect 4120 8192 4436 8193
rect 4120 8128 4126 8192
rect 4190 8128 4206 8192
rect 4270 8128 4286 8192
rect 4350 8128 4366 8192
rect 4430 8128 4436 8192
rect 4120 8127 4436 8128
rect 10468 8192 10784 8193
rect 10468 8128 10474 8192
rect 10538 8128 10554 8192
rect 10618 8128 10634 8192
rect 10698 8128 10714 8192
rect 10778 8128 10784 8192
rect 10468 8127 10784 8128
rect 16816 8192 17132 8193
rect 16816 8128 16822 8192
rect 16886 8128 16902 8192
rect 16966 8128 16982 8192
rect 17046 8128 17062 8192
rect 17126 8128 17132 8192
rect 16816 8127 17132 8128
rect 23164 8192 23480 8193
rect 23164 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23480 8192
rect 23164 8127 23480 8128
rect 7294 7648 7610 7649
rect 0 7578 800 7608
rect 7294 7584 7300 7648
rect 7364 7584 7380 7648
rect 7444 7584 7460 7648
rect 7524 7584 7540 7648
rect 7604 7584 7610 7648
rect 7294 7583 7610 7584
rect 13642 7648 13958 7649
rect 13642 7584 13648 7648
rect 13712 7584 13728 7648
rect 13792 7584 13808 7648
rect 13872 7584 13888 7648
rect 13952 7584 13958 7648
rect 13642 7583 13958 7584
rect 19990 7648 20306 7649
rect 19990 7584 19996 7648
rect 20060 7584 20076 7648
rect 20140 7584 20156 7648
rect 20220 7584 20236 7648
rect 20300 7584 20306 7648
rect 19990 7583 20306 7584
rect 26338 7648 26654 7649
rect 26338 7584 26344 7648
rect 26408 7584 26424 7648
rect 26488 7584 26504 7648
rect 26568 7584 26584 7648
rect 26648 7584 26654 7648
rect 26338 7583 26654 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 800 7518
rect 4061 7515 4127 7518
rect 4120 7104 4436 7105
rect 4120 7040 4126 7104
rect 4190 7040 4206 7104
rect 4270 7040 4286 7104
rect 4350 7040 4366 7104
rect 4430 7040 4436 7104
rect 4120 7039 4436 7040
rect 10468 7104 10784 7105
rect 10468 7040 10474 7104
rect 10538 7040 10554 7104
rect 10618 7040 10634 7104
rect 10698 7040 10714 7104
rect 10778 7040 10784 7104
rect 10468 7039 10784 7040
rect 16816 7104 17132 7105
rect 16816 7040 16822 7104
rect 16886 7040 16902 7104
rect 16966 7040 16982 7104
rect 17046 7040 17062 7104
rect 17126 7040 17132 7104
rect 16816 7039 17132 7040
rect 23164 7104 23480 7105
rect 23164 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23480 7104
rect 23164 7039 23480 7040
rect 7294 6560 7610 6561
rect 7294 6496 7300 6560
rect 7364 6496 7380 6560
rect 7444 6496 7460 6560
rect 7524 6496 7540 6560
rect 7604 6496 7610 6560
rect 7294 6495 7610 6496
rect 13642 6560 13958 6561
rect 13642 6496 13648 6560
rect 13712 6496 13728 6560
rect 13792 6496 13808 6560
rect 13872 6496 13888 6560
rect 13952 6496 13958 6560
rect 13642 6495 13958 6496
rect 19990 6560 20306 6561
rect 19990 6496 19996 6560
rect 20060 6496 20076 6560
rect 20140 6496 20156 6560
rect 20220 6496 20236 6560
rect 20300 6496 20306 6560
rect 19990 6495 20306 6496
rect 26338 6560 26654 6561
rect 26338 6496 26344 6560
rect 26408 6496 26424 6560
rect 26488 6496 26504 6560
rect 26568 6496 26584 6560
rect 26648 6496 26654 6560
rect 26338 6495 26654 6496
rect 4120 6016 4436 6017
rect 4120 5952 4126 6016
rect 4190 5952 4206 6016
rect 4270 5952 4286 6016
rect 4350 5952 4366 6016
rect 4430 5952 4436 6016
rect 4120 5951 4436 5952
rect 10468 6016 10784 6017
rect 10468 5952 10474 6016
rect 10538 5952 10554 6016
rect 10618 5952 10634 6016
rect 10698 5952 10714 6016
rect 10778 5952 10784 6016
rect 10468 5951 10784 5952
rect 16816 6016 17132 6017
rect 16816 5952 16822 6016
rect 16886 5952 16902 6016
rect 16966 5952 16982 6016
rect 17046 5952 17062 6016
rect 17126 5952 17132 6016
rect 16816 5951 17132 5952
rect 23164 6016 23480 6017
rect 23164 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23480 6016
rect 23164 5951 23480 5952
rect 7294 5472 7610 5473
rect 7294 5408 7300 5472
rect 7364 5408 7380 5472
rect 7444 5408 7460 5472
rect 7524 5408 7540 5472
rect 7604 5408 7610 5472
rect 7294 5407 7610 5408
rect 13642 5472 13958 5473
rect 13642 5408 13648 5472
rect 13712 5408 13728 5472
rect 13792 5408 13808 5472
rect 13872 5408 13888 5472
rect 13952 5408 13958 5472
rect 13642 5407 13958 5408
rect 19990 5472 20306 5473
rect 19990 5408 19996 5472
rect 20060 5408 20076 5472
rect 20140 5408 20156 5472
rect 20220 5408 20236 5472
rect 20300 5408 20306 5472
rect 19990 5407 20306 5408
rect 26338 5472 26654 5473
rect 26338 5408 26344 5472
rect 26408 5408 26424 5472
rect 26488 5408 26504 5472
rect 26568 5408 26584 5472
rect 26648 5408 26654 5472
rect 26338 5407 26654 5408
rect 4120 4928 4436 4929
rect 4120 4864 4126 4928
rect 4190 4864 4206 4928
rect 4270 4864 4286 4928
rect 4350 4864 4366 4928
rect 4430 4864 4436 4928
rect 4120 4863 4436 4864
rect 10468 4928 10784 4929
rect 10468 4864 10474 4928
rect 10538 4864 10554 4928
rect 10618 4864 10634 4928
rect 10698 4864 10714 4928
rect 10778 4864 10784 4928
rect 10468 4863 10784 4864
rect 16816 4928 17132 4929
rect 16816 4864 16822 4928
rect 16886 4864 16902 4928
rect 16966 4864 16982 4928
rect 17046 4864 17062 4928
rect 17126 4864 17132 4928
rect 16816 4863 17132 4864
rect 23164 4928 23480 4929
rect 23164 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23480 4928
rect 23164 4863 23480 4864
rect 26509 4858 26575 4861
rect 26841 4858 27641 4888
rect 26509 4856 27641 4858
rect 26509 4800 26514 4856
rect 26570 4800 27641 4856
rect 26509 4798 27641 4800
rect 26509 4795 26575 4798
rect 26841 4768 27641 4798
rect 7294 4384 7610 4385
rect 7294 4320 7300 4384
rect 7364 4320 7380 4384
rect 7444 4320 7460 4384
rect 7524 4320 7540 4384
rect 7604 4320 7610 4384
rect 7294 4319 7610 4320
rect 13642 4384 13958 4385
rect 13642 4320 13648 4384
rect 13712 4320 13728 4384
rect 13792 4320 13808 4384
rect 13872 4320 13888 4384
rect 13952 4320 13958 4384
rect 13642 4319 13958 4320
rect 19990 4384 20306 4385
rect 19990 4320 19996 4384
rect 20060 4320 20076 4384
rect 20140 4320 20156 4384
rect 20220 4320 20236 4384
rect 20300 4320 20306 4384
rect 19990 4319 20306 4320
rect 26338 4384 26654 4385
rect 26338 4320 26344 4384
rect 26408 4320 26424 4384
rect 26488 4320 26504 4384
rect 26568 4320 26584 4384
rect 26648 4320 26654 4384
rect 26338 4319 26654 4320
rect 13905 4178 13971 4181
rect 15193 4178 15259 4181
rect 13905 4176 15259 4178
rect 13905 4120 13910 4176
rect 13966 4120 15198 4176
rect 15254 4120 15259 4176
rect 13905 4118 15259 4120
rect 13905 4115 13971 4118
rect 15193 4115 15259 4118
rect 4120 3840 4436 3841
rect 4120 3776 4126 3840
rect 4190 3776 4206 3840
rect 4270 3776 4286 3840
rect 4350 3776 4366 3840
rect 4430 3776 4436 3840
rect 4120 3775 4436 3776
rect 10468 3840 10784 3841
rect 10468 3776 10474 3840
rect 10538 3776 10554 3840
rect 10618 3776 10634 3840
rect 10698 3776 10714 3840
rect 10778 3776 10784 3840
rect 10468 3775 10784 3776
rect 16816 3840 17132 3841
rect 16816 3776 16822 3840
rect 16886 3776 16902 3840
rect 16966 3776 16982 3840
rect 17046 3776 17062 3840
rect 17126 3776 17132 3840
rect 16816 3775 17132 3776
rect 23164 3840 23480 3841
rect 23164 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23480 3840
rect 23164 3775 23480 3776
rect 0 3408 800 3528
rect 14457 3362 14523 3365
rect 17033 3362 17099 3365
rect 14457 3360 17099 3362
rect 14457 3304 14462 3360
rect 14518 3304 17038 3360
rect 17094 3304 17099 3360
rect 14457 3302 17099 3304
rect 14457 3299 14523 3302
rect 17033 3299 17099 3302
rect 7294 3296 7610 3297
rect 7294 3232 7300 3296
rect 7364 3232 7380 3296
rect 7444 3232 7460 3296
rect 7524 3232 7540 3296
rect 7604 3232 7610 3296
rect 7294 3231 7610 3232
rect 13642 3296 13958 3297
rect 13642 3232 13648 3296
rect 13712 3232 13728 3296
rect 13792 3232 13808 3296
rect 13872 3232 13888 3296
rect 13952 3232 13958 3296
rect 13642 3231 13958 3232
rect 19990 3296 20306 3297
rect 19990 3232 19996 3296
rect 20060 3232 20076 3296
rect 20140 3232 20156 3296
rect 20220 3232 20236 3296
rect 20300 3232 20306 3296
rect 19990 3231 20306 3232
rect 26338 3296 26654 3297
rect 26338 3232 26344 3296
rect 26408 3232 26424 3296
rect 26488 3232 26504 3296
rect 26568 3232 26584 3296
rect 26648 3232 26654 3296
rect 26338 3231 26654 3232
rect 13353 3090 13419 3093
rect 15009 3090 15075 3093
rect 13353 3088 15075 3090
rect 13353 3032 13358 3088
rect 13414 3032 15014 3088
rect 15070 3032 15075 3088
rect 13353 3030 15075 3032
rect 13353 3027 13419 3030
rect 15009 3027 15075 3030
rect 4120 2752 4436 2753
rect 4120 2688 4126 2752
rect 4190 2688 4206 2752
rect 4270 2688 4286 2752
rect 4350 2688 4366 2752
rect 4430 2688 4436 2752
rect 4120 2687 4436 2688
rect 10468 2752 10784 2753
rect 10468 2688 10474 2752
rect 10538 2688 10554 2752
rect 10618 2688 10634 2752
rect 10698 2688 10714 2752
rect 10778 2688 10784 2752
rect 10468 2687 10784 2688
rect 16816 2752 17132 2753
rect 16816 2688 16822 2752
rect 16886 2688 16902 2752
rect 16966 2688 16982 2752
rect 17046 2688 17062 2752
rect 17126 2688 17132 2752
rect 16816 2687 17132 2688
rect 23164 2752 23480 2753
rect 23164 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23480 2752
rect 23164 2687 23480 2688
rect 7294 2208 7610 2209
rect 7294 2144 7300 2208
rect 7364 2144 7380 2208
rect 7444 2144 7460 2208
rect 7524 2144 7540 2208
rect 7604 2144 7610 2208
rect 7294 2143 7610 2144
rect 13642 2208 13958 2209
rect 13642 2144 13648 2208
rect 13712 2144 13728 2208
rect 13792 2144 13808 2208
rect 13872 2144 13888 2208
rect 13952 2144 13958 2208
rect 13642 2143 13958 2144
rect 19990 2208 20306 2209
rect 19990 2144 19996 2208
rect 20060 2144 20076 2208
rect 20140 2144 20156 2208
rect 20220 2144 20236 2208
rect 20300 2144 20306 2208
rect 19990 2143 20306 2144
rect 26338 2208 26654 2209
rect 26338 2144 26344 2208
rect 26408 2144 26424 2208
rect 26488 2144 26504 2208
rect 26568 2144 26584 2208
rect 26648 2144 26654 2208
rect 26338 2143 26654 2144
rect 26141 778 26207 781
rect 26841 778 27641 808
rect 26141 776 27641 778
rect 26141 720 26146 776
rect 26202 720 27641 776
rect 26141 718 27641 720
rect 26141 715 26207 718
rect 26841 688 27641 718
<< via3 >>
rect 7300 27228 7364 27232
rect 7300 27172 7304 27228
rect 7304 27172 7360 27228
rect 7360 27172 7364 27228
rect 7300 27168 7364 27172
rect 7380 27228 7444 27232
rect 7380 27172 7384 27228
rect 7384 27172 7440 27228
rect 7440 27172 7444 27228
rect 7380 27168 7444 27172
rect 7460 27228 7524 27232
rect 7460 27172 7464 27228
rect 7464 27172 7520 27228
rect 7520 27172 7524 27228
rect 7460 27168 7524 27172
rect 7540 27228 7604 27232
rect 7540 27172 7544 27228
rect 7544 27172 7600 27228
rect 7600 27172 7604 27228
rect 7540 27168 7604 27172
rect 13648 27228 13712 27232
rect 13648 27172 13652 27228
rect 13652 27172 13708 27228
rect 13708 27172 13712 27228
rect 13648 27168 13712 27172
rect 13728 27228 13792 27232
rect 13728 27172 13732 27228
rect 13732 27172 13788 27228
rect 13788 27172 13792 27228
rect 13728 27168 13792 27172
rect 13808 27228 13872 27232
rect 13808 27172 13812 27228
rect 13812 27172 13868 27228
rect 13868 27172 13872 27228
rect 13808 27168 13872 27172
rect 13888 27228 13952 27232
rect 13888 27172 13892 27228
rect 13892 27172 13948 27228
rect 13948 27172 13952 27228
rect 13888 27168 13952 27172
rect 19996 27228 20060 27232
rect 19996 27172 20000 27228
rect 20000 27172 20056 27228
rect 20056 27172 20060 27228
rect 19996 27168 20060 27172
rect 20076 27228 20140 27232
rect 20076 27172 20080 27228
rect 20080 27172 20136 27228
rect 20136 27172 20140 27228
rect 20076 27168 20140 27172
rect 20156 27228 20220 27232
rect 20156 27172 20160 27228
rect 20160 27172 20216 27228
rect 20216 27172 20220 27228
rect 20156 27168 20220 27172
rect 20236 27228 20300 27232
rect 20236 27172 20240 27228
rect 20240 27172 20296 27228
rect 20296 27172 20300 27228
rect 20236 27168 20300 27172
rect 26344 27228 26408 27232
rect 26344 27172 26348 27228
rect 26348 27172 26404 27228
rect 26404 27172 26408 27228
rect 26344 27168 26408 27172
rect 26424 27228 26488 27232
rect 26424 27172 26428 27228
rect 26428 27172 26484 27228
rect 26484 27172 26488 27228
rect 26424 27168 26488 27172
rect 26504 27228 26568 27232
rect 26504 27172 26508 27228
rect 26508 27172 26564 27228
rect 26564 27172 26568 27228
rect 26504 27168 26568 27172
rect 26584 27228 26648 27232
rect 26584 27172 26588 27228
rect 26588 27172 26644 27228
rect 26644 27172 26648 27228
rect 26584 27168 26648 27172
rect 4126 26684 4190 26688
rect 4126 26628 4130 26684
rect 4130 26628 4186 26684
rect 4186 26628 4190 26684
rect 4126 26624 4190 26628
rect 4206 26684 4270 26688
rect 4206 26628 4210 26684
rect 4210 26628 4266 26684
rect 4266 26628 4270 26684
rect 4206 26624 4270 26628
rect 4286 26684 4350 26688
rect 4286 26628 4290 26684
rect 4290 26628 4346 26684
rect 4346 26628 4350 26684
rect 4286 26624 4350 26628
rect 4366 26684 4430 26688
rect 4366 26628 4370 26684
rect 4370 26628 4426 26684
rect 4426 26628 4430 26684
rect 4366 26624 4430 26628
rect 10474 26684 10538 26688
rect 10474 26628 10478 26684
rect 10478 26628 10534 26684
rect 10534 26628 10538 26684
rect 10474 26624 10538 26628
rect 10554 26684 10618 26688
rect 10554 26628 10558 26684
rect 10558 26628 10614 26684
rect 10614 26628 10618 26684
rect 10554 26624 10618 26628
rect 10634 26684 10698 26688
rect 10634 26628 10638 26684
rect 10638 26628 10694 26684
rect 10694 26628 10698 26684
rect 10634 26624 10698 26628
rect 10714 26684 10778 26688
rect 10714 26628 10718 26684
rect 10718 26628 10774 26684
rect 10774 26628 10778 26684
rect 10714 26624 10778 26628
rect 16822 26684 16886 26688
rect 16822 26628 16826 26684
rect 16826 26628 16882 26684
rect 16882 26628 16886 26684
rect 16822 26624 16886 26628
rect 16902 26684 16966 26688
rect 16902 26628 16906 26684
rect 16906 26628 16962 26684
rect 16962 26628 16966 26684
rect 16902 26624 16966 26628
rect 16982 26684 17046 26688
rect 16982 26628 16986 26684
rect 16986 26628 17042 26684
rect 17042 26628 17046 26684
rect 16982 26624 17046 26628
rect 17062 26684 17126 26688
rect 17062 26628 17066 26684
rect 17066 26628 17122 26684
rect 17122 26628 17126 26684
rect 17062 26624 17126 26628
rect 23170 26684 23234 26688
rect 23170 26628 23174 26684
rect 23174 26628 23230 26684
rect 23230 26628 23234 26684
rect 23170 26624 23234 26628
rect 23250 26684 23314 26688
rect 23250 26628 23254 26684
rect 23254 26628 23310 26684
rect 23310 26628 23314 26684
rect 23250 26624 23314 26628
rect 23330 26684 23394 26688
rect 23330 26628 23334 26684
rect 23334 26628 23390 26684
rect 23390 26628 23394 26684
rect 23330 26624 23394 26628
rect 23410 26684 23474 26688
rect 23410 26628 23414 26684
rect 23414 26628 23470 26684
rect 23470 26628 23474 26684
rect 23410 26624 23474 26628
rect 7300 26140 7364 26144
rect 7300 26084 7304 26140
rect 7304 26084 7360 26140
rect 7360 26084 7364 26140
rect 7300 26080 7364 26084
rect 7380 26140 7444 26144
rect 7380 26084 7384 26140
rect 7384 26084 7440 26140
rect 7440 26084 7444 26140
rect 7380 26080 7444 26084
rect 7460 26140 7524 26144
rect 7460 26084 7464 26140
rect 7464 26084 7520 26140
rect 7520 26084 7524 26140
rect 7460 26080 7524 26084
rect 7540 26140 7604 26144
rect 7540 26084 7544 26140
rect 7544 26084 7600 26140
rect 7600 26084 7604 26140
rect 7540 26080 7604 26084
rect 13648 26140 13712 26144
rect 13648 26084 13652 26140
rect 13652 26084 13708 26140
rect 13708 26084 13712 26140
rect 13648 26080 13712 26084
rect 13728 26140 13792 26144
rect 13728 26084 13732 26140
rect 13732 26084 13788 26140
rect 13788 26084 13792 26140
rect 13728 26080 13792 26084
rect 13808 26140 13872 26144
rect 13808 26084 13812 26140
rect 13812 26084 13868 26140
rect 13868 26084 13872 26140
rect 13808 26080 13872 26084
rect 13888 26140 13952 26144
rect 13888 26084 13892 26140
rect 13892 26084 13948 26140
rect 13948 26084 13952 26140
rect 13888 26080 13952 26084
rect 19996 26140 20060 26144
rect 19996 26084 20000 26140
rect 20000 26084 20056 26140
rect 20056 26084 20060 26140
rect 19996 26080 20060 26084
rect 20076 26140 20140 26144
rect 20076 26084 20080 26140
rect 20080 26084 20136 26140
rect 20136 26084 20140 26140
rect 20076 26080 20140 26084
rect 20156 26140 20220 26144
rect 20156 26084 20160 26140
rect 20160 26084 20216 26140
rect 20216 26084 20220 26140
rect 20156 26080 20220 26084
rect 20236 26140 20300 26144
rect 20236 26084 20240 26140
rect 20240 26084 20296 26140
rect 20296 26084 20300 26140
rect 20236 26080 20300 26084
rect 26344 26140 26408 26144
rect 26344 26084 26348 26140
rect 26348 26084 26404 26140
rect 26404 26084 26408 26140
rect 26344 26080 26408 26084
rect 26424 26140 26488 26144
rect 26424 26084 26428 26140
rect 26428 26084 26484 26140
rect 26484 26084 26488 26140
rect 26424 26080 26488 26084
rect 26504 26140 26568 26144
rect 26504 26084 26508 26140
rect 26508 26084 26564 26140
rect 26564 26084 26568 26140
rect 26504 26080 26568 26084
rect 26584 26140 26648 26144
rect 26584 26084 26588 26140
rect 26588 26084 26644 26140
rect 26644 26084 26648 26140
rect 26584 26080 26648 26084
rect 4126 25596 4190 25600
rect 4126 25540 4130 25596
rect 4130 25540 4186 25596
rect 4186 25540 4190 25596
rect 4126 25536 4190 25540
rect 4206 25596 4270 25600
rect 4206 25540 4210 25596
rect 4210 25540 4266 25596
rect 4266 25540 4270 25596
rect 4206 25536 4270 25540
rect 4286 25596 4350 25600
rect 4286 25540 4290 25596
rect 4290 25540 4346 25596
rect 4346 25540 4350 25596
rect 4286 25536 4350 25540
rect 4366 25596 4430 25600
rect 4366 25540 4370 25596
rect 4370 25540 4426 25596
rect 4426 25540 4430 25596
rect 4366 25536 4430 25540
rect 10474 25596 10538 25600
rect 10474 25540 10478 25596
rect 10478 25540 10534 25596
rect 10534 25540 10538 25596
rect 10474 25536 10538 25540
rect 10554 25596 10618 25600
rect 10554 25540 10558 25596
rect 10558 25540 10614 25596
rect 10614 25540 10618 25596
rect 10554 25536 10618 25540
rect 10634 25596 10698 25600
rect 10634 25540 10638 25596
rect 10638 25540 10694 25596
rect 10694 25540 10698 25596
rect 10634 25536 10698 25540
rect 10714 25596 10778 25600
rect 10714 25540 10718 25596
rect 10718 25540 10774 25596
rect 10774 25540 10778 25596
rect 10714 25536 10778 25540
rect 16822 25596 16886 25600
rect 16822 25540 16826 25596
rect 16826 25540 16882 25596
rect 16882 25540 16886 25596
rect 16822 25536 16886 25540
rect 16902 25596 16966 25600
rect 16902 25540 16906 25596
rect 16906 25540 16962 25596
rect 16962 25540 16966 25596
rect 16902 25536 16966 25540
rect 16982 25596 17046 25600
rect 16982 25540 16986 25596
rect 16986 25540 17042 25596
rect 17042 25540 17046 25596
rect 16982 25536 17046 25540
rect 17062 25596 17126 25600
rect 17062 25540 17066 25596
rect 17066 25540 17122 25596
rect 17122 25540 17126 25596
rect 17062 25536 17126 25540
rect 23170 25596 23234 25600
rect 23170 25540 23174 25596
rect 23174 25540 23230 25596
rect 23230 25540 23234 25596
rect 23170 25536 23234 25540
rect 23250 25596 23314 25600
rect 23250 25540 23254 25596
rect 23254 25540 23310 25596
rect 23310 25540 23314 25596
rect 23250 25536 23314 25540
rect 23330 25596 23394 25600
rect 23330 25540 23334 25596
rect 23334 25540 23390 25596
rect 23390 25540 23394 25596
rect 23330 25536 23394 25540
rect 23410 25596 23474 25600
rect 23410 25540 23414 25596
rect 23414 25540 23470 25596
rect 23470 25540 23474 25596
rect 23410 25536 23474 25540
rect 7300 25052 7364 25056
rect 7300 24996 7304 25052
rect 7304 24996 7360 25052
rect 7360 24996 7364 25052
rect 7300 24992 7364 24996
rect 7380 25052 7444 25056
rect 7380 24996 7384 25052
rect 7384 24996 7440 25052
rect 7440 24996 7444 25052
rect 7380 24992 7444 24996
rect 7460 25052 7524 25056
rect 7460 24996 7464 25052
rect 7464 24996 7520 25052
rect 7520 24996 7524 25052
rect 7460 24992 7524 24996
rect 7540 25052 7604 25056
rect 7540 24996 7544 25052
rect 7544 24996 7600 25052
rect 7600 24996 7604 25052
rect 7540 24992 7604 24996
rect 13648 25052 13712 25056
rect 13648 24996 13652 25052
rect 13652 24996 13708 25052
rect 13708 24996 13712 25052
rect 13648 24992 13712 24996
rect 13728 25052 13792 25056
rect 13728 24996 13732 25052
rect 13732 24996 13788 25052
rect 13788 24996 13792 25052
rect 13728 24992 13792 24996
rect 13808 25052 13872 25056
rect 13808 24996 13812 25052
rect 13812 24996 13868 25052
rect 13868 24996 13872 25052
rect 13808 24992 13872 24996
rect 13888 25052 13952 25056
rect 13888 24996 13892 25052
rect 13892 24996 13948 25052
rect 13948 24996 13952 25052
rect 13888 24992 13952 24996
rect 19996 25052 20060 25056
rect 19996 24996 20000 25052
rect 20000 24996 20056 25052
rect 20056 24996 20060 25052
rect 19996 24992 20060 24996
rect 20076 25052 20140 25056
rect 20076 24996 20080 25052
rect 20080 24996 20136 25052
rect 20136 24996 20140 25052
rect 20076 24992 20140 24996
rect 20156 25052 20220 25056
rect 20156 24996 20160 25052
rect 20160 24996 20216 25052
rect 20216 24996 20220 25052
rect 20156 24992 20220 24996
rect 20236 25052 20300 25056
rect 20236 24996 20240 25052
rect 20240 24996 20296 25052
rect 20296 24996 20300 25052
rect 20236 24992 20300 24996
rect 26344 25052 26408 25056
rect 26344 24996 26348 25052
rect 26348 24996 26404 25052
rect 26404 24996 26408 25052
rect 26344 24992 26408 24996
rect 26424 25052 26488 25056
rect 26424 24996 26428 25052
rect 26428 24996 26484 25052
rect 26484 24996 26488 25052
rect 26424 24992 26488 24996
rect 26504 25052 26568 25056
rect 26504 24996 26508 25052
rect 26508 24996 26564 25052
rect 26564 24996 26568 25052
rect 26504 24992 26568 24996
rect 26584 25052 26648 25056
rect 26584 24996 26588 25052
rect 26588 24996 26644 25052
rect 26644 24996 26648 25052
rect 26584 24992 26648 24996
rect 4126 24508 4190 24512
rect 4126 24452 4130 24508
rect 4130 24452 4186 24508
rect 4186 24452 4190 24508
rect 4126 24448 4190 24452
rect 4206 24508 4270 24512
rect 4206 24452 4210 24508
rect 4210 24452 4266 24508
rect 4266 24452 4270 24508
rect 4206 24448 4270 24452
rect 4286 24508 4350 24512
rect 4286 24452 4290 24508
rect 4290 24452 4346 24508
rect 4346 24452 4350 24508
rect 4286 24448 4350 24452
rect 4366 24508 4430 24512
rect 4366 24452 4370 24508
rect 4370 24452 4426 24508
rect 4426 24452 4430 24508
rect 4366 24448 4430 24452
rect 10474 24508 10538 24512
rect 10474 24452 10478 24508
rect 10478 24452 10534 24508
rect 10534 24452 10538 24508
rect 10474 24448 10538 24452
rect 10554 24508 10618 24512
rect 10554 24452 10558 24508
rect 10558 24452 10614 24508
rect 10614 24452 10618 24508
rect 10554 24448 10618 24452
rect 10634 24508 10698 24512
rect 10634 24452 10638 24508
rect 10638 24452 10694 24508
rect 10694 24452 10698 24508
rect 10634 24448 10698 24452
rect 10714 24508 10778 24512
rect 10714 24452 10718 24508
rect 10718 24452 10774 24508
rect 10774 24452 10778 24508
rect 10714 24448 10778 24452
rect 16822 24508 16886 24512
rect 16822 24452 16826 24508
rect 16826 24452 16882 24508
rect 16882 24452 16886 24508
rect 16822 24448 16886 24452
rect 16902 24508 16966 24512
rect 16902 24452 16906 24508
rect 16906 24452 16962 24508
rect 16962 24452 16966 24508
rect 16902 24448 16966 24452
rect 16982 24508 17046 24512
rect 16982 24452 16986 24508
rect 16986 24452 17042 24508
rect 17042 24452 17046 24508
rect 16982 24448 17046 24452
rect 17062 24508 17126 24512
rect 17062 24452 17066 24508
rect 17066 24452 17122 24508
rect 17122 24452 17126 24508
rect 17062 24448 17126 24452
rect 23170 24508 23234 24512
rect 23170 24452 23174 24508
rect 23174 24452 23230 24508
rect 23230 24452 23234 24508
rect 23170 24448 23234 24452
rect 23250 24508 23314 24512
rect 23250 24452 23254 24508
rect 23254 24452 23310 24508
rect 23310 24452 23314 24508
rect 23250 24448 23314 24452
rect 23330 24508 23394 24512
rect 23330 24452 23334 24508
rect 23334 24452 23390 24508
rect 23390 24452 23394 24508
rect 23330 24448 23394 24452
rect 23410 24508 23474 24512
rect 23410 24452 23414 24508
rect 23414 24452 23470 24508
rect 23470 24452 23474 24508
rect 23410 24448 23474 24452
rect 7300 23964 7364 23968
rect 7300 23908 7304 23964
rect 7304 23908 7360 23964
rect 7360 23908 7364 23964
rect 7300 23904 7364 23908
rect 7380 23964 7444 23968
rect 7380 23908 7384 23964
rect 7384 23908 7440 23964
rect 7440 23908 7444 23964
rect 7380 23904 7444 23908
rect 7460 23964 7524 23968
rect 7460 23908 7464 23964
rect 7464 23908 7520 23964
rect 7520 23908 7524 23964
rect 7460 23904 7524 23908
rect 7540 23964 7604 23968
rect 7540 23908 7544 23964
rect 7544 23908 7600 23964
rect 7600 23908 7604 23964
rect 7540 23904 7604 23908
rect 13648 23964 13712 23968
rect 13648 23908 13652 23964
rect 13652 23908 13708 23964
rect 13708 23908 13712 23964
rect 13648 23904 13712 23908
rect 13728 23964 13792 23968
rect 13728 23908 13732 23964
rect 13732 23908 13788 23964
rect 13788 23908 13792 23964
rect 13728 23904 13792 23908
rect 13808 23964 13872 23968
rect 13808 23908 13812 23964
rect 13812 23908 13868 23964
rect 13868 23908 13872 23964
rect 13808 23904 13872 23908
rect 13888 23964 13952 23968
rect 13888 23908 13892 23964
rect 13892 23908 13948 23964
rect 13948 23908 13952 23964
rect 13888 23904 13952 23908
rect 19996 23964 20060 23968
rect 19996 23908 20000 23964
rect 20000 23908 20056 23964
rect 20056 23908 20060 23964
rect 19996 23904 20060 23908
rect 20076 23964 20140 23968
rect 20076 23908 20080 23964
rect 20080 23908 20136 23964
rect 20136 23908 20140 23964
rect 20076 23904 20140 23908
rect 20156 23964 20220 23968
rect 20156 23908 20160 23964
rect 20160 23908 20216 23964
rect 20216 23908 20220 23964
rect 20156 23904 20220 23908
rect 20236 23964 20300 23968
rect 20236 23908 20240 23964
rect 20240 23908 20296 23964
rect 20296 23908 20300 23964
rect 20236 23904 20300 23908
rect 26344 23964 26408 23968
rect 26344 23908 26348 23964
rect 26348 23908 26404 23964
rect 26404 23908 26408 23964
rect 26344 23904 26408 23908
rect 26424 23964 26488 23968
rect 26424 23908 26428 23964
rect 26428 23908 26484 23964
rect 26484 23908 26488 23964
rect 26424 23904 26488 23908
rect 26504 23964 26568 23968
rect 26504 23908 26508 23964
rect 26508 23908 26564 23964
rect 26564 23908 26568 23964
rect 26504 23904 26568 23908
rect 26584 23964 26648 23968
rect 26584 23908 26588 23964
rect 26588 23908 26644 23964
rect 26644 23908 26648 23964
rect 26584 23904 26648 23908
rect 4126 23420 4190 23424
rect 4126 23364 4130 23420
rect 4130 23364 4186 23420
rect 4186 23364 4190 23420
rect 4126 23360 4190 23364
rect 4206 23420 4270 23424
rect 4206 23364 4210 23420
rect 4210 23364 4266 23420
rect 4266 23364 4270 23420
rect 4206 23360 4270 23364
rect 4286 23420 4350 23424
rect 4286 23364 4290 23420
rect 4290 23364 4346 23420
rect 4346 23364 4350 23420
rect 4286 23360 4350 23364
rect 4366 23420 4430 23424
rect 4366 23364 4370 23420
rect 4370 23364 4426 23420
rect 4426 23364 4430 23420
rect 4366 23360 4430 23364
rect 10474 23420 10538 23424
rect 10474 23364 10478 23420
rect 10478 23364 10534 23420
rect 10534 23364 10538 23420
rect 10474 23360 10538 23364
rect 10554 23420 10618 23424
rect 10554 23364 10558 23420
rect 10558 23364 10614 23420
rect 10614 23364 10618 23420
rect 10554 23360 10618 23364
rect 10634 23420 10698 23424
rect 10634 23364 10638 23420
rect 10638 23364 10694 23420
rect 10694 23364 10698 23420
rect 10634 23360 10698 23364
rect 10714 23420 10778 23424
rect 10714 23364 10718 23420
rect 10718 23364 10774 23420
rect 10774 23364 10778 23420
rect 10714 23360 10778 23364
rect 16822 23420 16886 23424
rect 16822 23364 16826 23420
rect 16826 23364 16882 23420
rect 16882 23364 16886 23420
rect 16822 23360 16886 23364
rect 16902 23420 16966 23424
rect 16902 23364 16906 23420
rect 16906 23364 16962 23420
rect 16962 23364 16966 23420
rect 16902 23360 16966 23364
rect 16982 23420 17046 23424
rect 16982 23364 16986 23420
rect 16986 23364 17042 23420
rect 17042 23364 17046 23420
rect 16982 23360 17046 23364
rect 17062 23420 17126 23424
rect 17062 23364 17066 23420
rect 17066 23364 17122 23420
rect 17122 23364 17126 23420
rect 17062 23360 17126 23364
rect 23170 23420 23234 23424
rect 23170 23364 23174 23420
rect 23174 23364 23230 23420
rect 23230 23364 23234 23420
rect 23170 23360 23234 23364
rect 23250 23420 23314 23424
rect 23250 23364 23254 23420
rect 23254 23364 23310 23420
rect 23310 23364 23314 23420
rect 23250 23360 23314 23364
rect 23330 23420 23394 23424
rect 23330 23364 23334 23420
rect 23334 23364 23390 23420
rect 23390 23364 23394 23420
rect 23330 23360 23394 23364
rect 23410 23420 23474 23424
rect 23410 23364 23414 23420
rect 23414 23364 23470 23420
rect 23470 23364 23474 23420
rect 23410 23360 23474 23364
rect 7300 22876 7364 22880
rect 7300 22820 7304 22876
rect 7304 22820 7360 22876
rect 7360 22820 7364 22876
rect 7300 22816 7364 22820
rect 7380 22876 7444 22880
rect 7380 22820 7384 22876
rect 7384 22820 7440 22876
rect 7440 22820 7444 22876
rect 7380 22816 7444 22820
rect 7460 22876 7524 22880
rect 7460 22820 7464 22876
rect 7464 22820 7520 22876
rect 7520 22820 7524 22876
rect 7460 22816 7524 22820
rect 7540 22876 7604 22880
rect 7540 22820 7544 22876
rect 7544 22820 7600 22876
rect 7600 22820 7604 22876
rect 7540 22816 7604 22820
rect 13648 22876 13712 22880
rect 13648 22820 13652 22876
rect 13652 22820 13708 22876
rect 13708 22820 13712 22876
rect 13648 22816 13712 22820
rect 13728 22876 13792 22880
rect 13728 22820 13732 22876
rect 13732 22820 13788 22876
rect 13788 22820 13792 22876
rect 13728 22816 13792 22820
rect 13808 22876 13872 22880
rect 13808 22820 13812 22876
rect 13812 22820 13868 22876
rect 13868 22820 13872 22876
rect 13808 22816 13872 22820
rect 13888 22876 13952 22880
rect 13888 22820 13892 22876
rect 13892 22820 13948 22876
rect 13948 22820 13952 22876
rect 13888 22816 13952 22820
rect 19996 22876 20060 22880
rect 19996 22820 20000 22876
rect 20000 22820 20056 22876
rect 20056 22820 20060 22876
rect 19996 22816 20060 22820
rect 20076 22876 20140 22880
rect 20076 22820 20080 22876
rect 20080 22820 20136 22876
rect 20136 22820 20140 22876
rect 20076 22816 20140 22820
rect 20156 22876 20220 22880
rect 20156 22820 20160 22876
rect 20160 22820 20216 22876
rect 20216 22820 20220 22876
rect 20156 22816 20220 22820
rect 20236 22876 20300 22880
rect 20236 22820 20240 22876
rect 20240 22820 20296 22876
rect 20296 22820 20300 22876
rect 20236 22816 20300 22820
rect 26344 22876 26408 22880
rect 26344 22820 26348 22876
rect 26348 22820 26404 22876
rect 26404 22820 26408 22876
rect 26344 22816 26408 22820
rect 26424 22876 26488 22880
rect 26424 22820 26428 22876
rect 26428 22820 26484 22876
rect 26484 22820 26488 22876
rect 26424 22816 26488 22820
rect 26504 22876 26568 22880
rect 26504 22820 26508 22876
rect 26508 22820 26564 22876
rect 26564 22820 26568 22876
rect 26504 22816 26568 22820
rect 26584 22876 26648 22880
rect 26584 22820 26588 22876
rect 26588 22820 26644 22876
rect 26644 22820 26648 22876
rect 26584 22816 26648 22820
rect 4126 22332 4190 22336
rect 4126 22276 4130 22332
rect 4130 22276 4186 22332
rect 4186 22276 4190 22332
rect 4126 22272 4190 22276
rect 4206 22332 4270 22336
rect 4206 22276 4210 22332
rect 4210 22276 4266 22332
rect 4266 22276 4270 22332
rect 4206 22272 4270 22276
rect 4286 22332 4350 22336
rect 4286 22276 4290 22332
rect 4290 22276 4346 22332
rect 4346 22276 4350 22332
rect 4286 22272 4350 22276
rect 4366 22332 4430 22336
rect 4366 22276 4370 22332
rect 4370 22276 4426 22332
rect 4426 22276 4430 22332
rect 4366 22272 4430 22276
rect 10474 22332 10538 22336
rect 10474 22276 10478 22332
rect 10478 22276 10534 22332
rect 10534 22276 10538 22332
rect 10474 22272 10538 22276
rect 10554 22332 10618 22336
rect 10554 22276 10558 22332
rect 10558 22276 10614 22332
rect 10614 22276 10618 22332
rect 10554 22272 10618 22276
rect 10634 22332 10698 22336
rect 10634 22276 10638 22332
rect 10638 22276 10694 22332
rect 10694 22276 10698 22332
rect 10634 22272 10698 22276
rect 10714 22332 10778 22336
rect 10714 22276 10718 22332
rect 10718 22276 10774 22332
rect 10774 22276 10778 22332
rect 10714 22272 10778 22276
rect 16822 22332 16886 22336
rect 16822 22276 16826 22332
rect 16826 22276 16882 22332
rect 16882 22276 16886 22332
rect 16822 22272 16886 22276
rect 16902 22332 16966 22336
rect 16902 22276 16906 22332
rect 16906 22276 16962 22332
rect 16962 22276 16966 22332
rect 16902 22272 16966 22276
rect 16982 22332 17046 22336
rect 16982 22276 16986 22332
rect 16986 22276 17042 22332
rect 17042 22276 17046 22332
rect 16982 22272 17046 22276
rect 17062 22332 17126 22336
rect 17062 22276 17066 22332
rect 17066 22276 17122 22332
rect 17122 22276 17126 22332
rect 17062 22272 17126 22276
rect 23170 22332 23234 22336
rect 23170 22276 23174 22332
rect 23174 22276 23230 22332
rect 23230 22276 23234 22332
rect 23170 22272 23234 22276
rect 23250 22332 23314 22336
rect 23250 22276 23254 22332
rect 23254 22276 23310 22332
rect 23310 22276 23314 22332
rect 23250 22272 23314 22276
rect 23330 22332 23394 22336
rect 23330 22276 23334 22332
rect 23334 22276 23390 22332
rect 23390 22276 23394 22332
rect 23330 22272 23394 22276
rect 23410 22332 23474 22336
rect 23410 22276 23414 22332
rect 23414 22276 23470 22332
rect 23470 22276 23474 22332
rect 23410 22272 23474 22276
rect 7300 21788 7364 21792
rect 7300 21732 7304 21788
rect 7304 21732 7360 21788
rect 7360 21732 7364 21788
rect 7300 21728 7364 21732
rect 7380 21788 7444 21792
rect 7380 21732 7384 21788
rect 7384 21732 7440 21788
rect 7440 21732 7444 21788
rect 7380 21728 7444 21732
rect 7460 21788 7524 21792
rect 7460 21732 7464 21788
rect 7464 21732 7520 21788
rect 7520 21732 7524 21788
rect 7460 21728 7524 21732
rect 7540 21788 7604 21792
rect 7540 21732 7544 21788
rect 7544 21732 7600 21788
rect 7600 21732 7604 21788
rect 7540 21728 7604 21732
rect 13648 21788 13712 21792
rect 13648 21732 13652 21788
rect 13652 21732 13708 21788
rect 13708 21732 13712 21788
rect 13648 21728 13712 21732
rect 13728 21788 13792 21792
rect 13728 21732 13732 21788
rect 13732 21732 13788 21788
rect 13788 21732 13792 21788
rect 13728 21728 13792 21732
rect 13808 21788 13872 21792
rect 13808 21732 13812 21788
rect 13812 21732 13868 21788
rect 13868 21732 13872 21788
rect 13808 21728 13872 21732
rect 13888 21788 13952 21792
rect 13888 21732 13892 21788
rect 13892 21732 13948 21788
rect 13948 21732 13952 21788
rect 13888 21728 13952 21732
rect 19996 21788 20060 21792
rect 19996 21732 20000 21788
rect 20000 21732 20056 21788
rect 20056 21732 20060 21788
rect 19996 21728 20060 21732
rect 20076 21788 20140 21792
rect 20076 21732 20080 21788
rect 20080 21732 20136 21788
rect 20136 21732 20140 21788
rect 20076 21728 20140 21732
rect 20156 21788 20220 21792
rect 20156 21732 20160 21788
rect 20160 21732 20216 21788
rect 20216 21732 20220 21788
rect 20156 21728 20220 21732
rect 20236 21788 20300 21792
rect 20236 21732 20240 21788
rect 20240 21732 20296 21788
rect 20296 21732 20300 21788
rect 20236 21728 20300 21732
rect 26344 21788 26408 21792
rect 26344 21732 26348 21788
rect 26348 21732 26404 21788
rect 26404 21732 26408 21788
rect 26344 21728 26408 21732
rect 26424 21788 26488 21792
rect 26424 21732 26428 21788
rect 26428 21732 26484 21788
rect 26484 21732 26488 21788
rect 26424 21728 26488 21732
rect 26504 21788 26568 21792
rect 26504 21732 26508 21788
rect 26508 21732 26564 21788
rect 26564 21732 26568 21788
rect 26504 21728 26568 21732
rect 26584 21788 26648 21792
rect 26584 21732 26588 21788
rect 26588 21732 26644 21788
rect 26644 21732 26648 21788
rect 26584 21728 26648 21732
rect 4126 21244 4190 21248
rect 4126 21188 4130 21244
rect 4130 21188 4186 21244
rect 4186 21188 4190 21244
rect 4126 21184 4190 21188
rect 4206 21244 4270 21248
rect 4206 21188 4210 21244
rect 4210 21188 4266 21244
rect 4266 21188 4270 21244
rect 4206 21184 4270 21188
rect 4286 21244 4350 21248
rect 4286 21188 4290 21244
rect 4290 21188 4346 21244
rect 4346 21188 4350 21244
rect 4286 21184 4350 21188
rect 4366 21244 4430 21248
rect 4366 21188 4370 21244
rect 4370 21188 4426 21244
rect 4426 21188 4430 21244
rect 4366 21184 4430 21188
rect 10474 21244 10538 21248
rect 10474 21188 10478 21244
rect 10478 21188 10534 21244
rect 10534 21188 10538 21244
rect 10474 21184 10538 21188
rect 10554 21244 10618 21248
rect 10554 21188 10558 21244
rect 10558 21188 10614 21244
rect 10614 21188 10618 21244
rect 10554 21184 10618 21188
rect 10634 21244 10698 21248
rect 10634 21188 10638 21244
rect 10638 21188 10694 21244
rect 10694 21188 10698 21244
rect 10634 21184 10698 21188
rect 10714 21244 10778 21248
rect 10714 21188 10718 21244
rect 10718 21188 10774 21244
rect 10774 21188 10778 21244
rect 10714 21184 10778 21188
rect 16822 21244 16886 21248
rect 16822 21188 16826 21244
rect 16826 21188 16882 21244
rect 16882 21188 16886 21244
rect 16822 21184 16886 21188
rect 16902 21244 16966 21248
rect 16902 21188 16906 21244
rect 16906 21188 16962 21244
rect 16962 21188 16966 21244
rect 16902 21184 16966 21188
rect 16982 21244 17046 21248
rect 16982 21188 16986 21244
rect 16986 21188 17042 21244
rect 17042 21188 17046 21244
rect 16982 21184 17046 21188
rect 17062 21244 17126 21248
rect 17062 21188 17066 21244
rect 17066 21188 17122 21244
rect 17122 21188 17126 21244
rect 17062 21184 17126 21188
rect 23170 21244 23234 21248
rect 23170 21188 23174 21244
rect 23174 21188 23230 21244
rect 23230 21188 23234 21244
rect 23170 21184 23234 21188
rect 23250 21244 23314 21248
rect 23250 21188 23254 21244
rect 23254 21188 23310 21244
rect 23310 21188 23314 21244
rect 23250 21184 23314 21188
rect 23330 21244 23394 21248
rect 23330 21188 23334 21244
rect 23334 21188 23390 21244
rect 23390 21188 23394 21244
rect 23330 21184 23394 21188
rect 23410 21244 23474 21248
rect 23410 21188 23414 21244
rect 23414 21188 23470 21244
rect 23470 21188 23474 21244
rect 23410 21184 23474 21188
rect 7300 20700 7364 20704
rect 7300 20644 7304 20700
rect 7304 20644 7360 20700
rect 7360 20644 7364 20700
rect 7300 20640 7364 20644
rect 7380 20700 7444 20704
rect 7380 20644 7384 20700
rect 7384 20644 7440 20700
rect 7440 20644 7444 20700
rect 7380 20640 7444 20644
rect 7460 20700 7524 20704
rect 7460 20644 7464 20700
rect 7464 20644 7520 20700
rect 7520 20644 7524 20700
rect 7460 20640 7524 20644
rect 7540 20700 7604 20704
rect 7540 20644 7544 20700
rect 7544 20644 7600 20700
rect 7600 20644 7604 20700
rect 7540 20640 7604 20644
rect 13648 20700 13712 20704
rect 13648 20644 13652 20700
rect 13652 20644 13708 20700
rect 13708 20644 13712 20700
rect 13648 20640 13712 20644
rect 13728 20700 13792 20704
rect 13728 20644 13732 20700
rect 13732 20644 13788 20700
rect 13788 20644 13792 20700
rect 13728 20640 13792 20644
rect 13808 20700 13872 20704
rect 13808 20644 13812 20700
rect 13812 20644 13868 20700
rect 13868 20644 13872 20700
rect 13808 20640 13872 20644
rect 13888 20700 13952 20704
rect 13888 20644 13892 20700
rect 13892 20644 13948 20700
rect 13948 20644 13952 20700
rect 13888 20640 13952 20644
rect 19996 20700 20060 20704
rect 19996 20644 20000 20700
rect 20000 20644 20056 20700
rect 20056 20644 20060 20700
rect 19996 20640 20060 20644
rect 20076 20700 20140 20704
rect 20076 20644 20080 20700
rect 20080 20644 20136 20700
rect 20136 20644 20140 20700
rect 20076 20640 20140 20644
rect 20156 20700 20220 20704
rect 20156 20644 20160 20700
rect 20160 20644 20216 20700
rect 20216 20644 20220 20700
rect 20156 20640 20220 20644
rect 20236 20700 20300 20704
rect 20236 20644 20240 20700
rect 20240 20644 20296 20700
rect 20296 20644 20300 20700
rect 20236 20640 20300 20644
rect 26344 20700 26408 20704
rect 26344 20644 26348 20700
rect 26348 20644 26404 20700
rect 26404 20644 26408 20700
rect 26344 20640 26408 20644
rect 26424 20700 26488 20704
rect 26424 20644 26428 20700
rect 26428 20644 26484 20700
rect 26484 20644 26488 20700
rect 26424 20640 26488 20644
rect 26504 20700 26568 20704
rect 26504 20644 26508 20700
rect 26508 20644 26564 20700
rect 26564 20644 26568 20700
rect 26504 20640 26568 20644
rect 26584 20700 26648 20704
rect 26584 20644 26588 20700
rect 26588 20644 26644 20700
rect 26644 20644 26648 20700
rect 26584 20640 26648 20644
rect 4126 20156 4190 20160
rect 4126 20100 4130 20156
rect 4130 20100 4186 20156
rect 4186 20100 4190 20156
rect 4126 20096 4190 20100
rect 4206 20156 4270 20160
rect 4206 20100 4210 20156
rect 4210 20100 4266 20156
rect 4266 20100 4270 20156
rect 4206 20096 4270 20100
rect 4286 20156 4350 20160
rect 4286 20100 4290 20156
rect 4290 20100 4346 20156
rect 4346 20100 4350 20156
rect 4286 20096 4350 20100
rect 4366 20156 4430 20160
rect 4366 20100 4370 20156
rect 4370 20100 4426 20156
rect 4426 20100 4430 20156
rect 4366 20096 4430 20100
rect 10474 20156 10538 20160
rect 10474 20100 10478 20156
rect 10478 20100 10534 20156
rect 10534 20100 10538 20156
rect 10474 20096 10538 20100
rect 10554 20156 10618 20160
rect 10554 20100 10558 20156
rect 10558 20100 10614 20156
rect 10614 20100 10618 20156
rect 10554 20096 10618 20100
rect 10634 20156 10698 20160
rect 10634 20100 10638 20156
rect 10638 20100 10694 20156
rect 10694 20100 10698 20156
rect 10634 20096 10698 20100
rect 10714 20156 10778 20160
rect 10714 20100 10718 20156
rect 10718 20100 10774 20156
rect 10774 20100 10778 20156
rect 10714 20096 10778 20100
rect 16822 20156 16886 20160
rect 16822 20100 16826 20156
rect 16826 20100 16882 20156
rect 16882 20100 16886 20156
rect 16822 20096 16886 20100
rect 16902 20156 16966 20160
rect 16902 20100 16906 20156
rect 16906 20100 16962 20156
rect 16962 20100 16966 20156
rect 16902 20096 16966 20100
rect 16982 20156 17046 20160
rect 16982 20100 16986 20156
rect 16986 20100 17042 20156
rect 17042 20100 17046 20156
rect 16982 20096 17046 20100
rect 17062 20156 17126 20160
rect 17062 20100 17066 20156
rect 17066 20100 17122 20156
rect 17122 20100 17126 20156
rect 17062 20096 17126 20100
rect 23170 20156 23234 20160
rect 23170 20100 23174 20156
rect 23174 20100 23230 20156
rect 23230 20100 23234 20156
rect 23170 20096 23234 20100
rect 23250 20156 23314 20160
rect 23250 20100 23254 20156
rect 23254 20100 23310 20156
rect 23310 20100 23314 20156
rect 23250 20096 23314 20100
rect 23330 20156 23394 20160
rect 23330 20100 23334 20156
rect 23334 20100 23390 20156
rect 23390 20100 23394 20156
rect 23330 20096 23394 20100
rect 23410 20156 23474 20160
rect 23410 20100 23414 20156
rect 23414 20100 23470 20156
rect 23470 20100 23474 20156
rect 23410 20096 23474 20100
rect 7300 19612 7364 19616
rect 7300 19556 7304 19612
rect 7304 19556 7360 19612
rect 7360 19556 7364 19612
rect 7300 19552 7364 19556
rect 7380 19612 7444 19616
rect 7380 19556 7384 19612
rect 7384 19556 7440 19612
rect 7440 19556 7444 19612
rect 7380 19552 7444 19556
rect 7460 19612 7524 19616
rect 7460 19556 7464 19612
rect 7464 19556 7520 19612
rect 7520 19556 7524 19612
rect 7460 19552 7524 19556
rect 7540 19612 7604 19616
rect 7540 19556 7544 19612
rect 7544 19556 7600 19612
rect 7600 19556 7604 19612
rect 7540 19552 7604 19556
rect 13648 19612 13712 19616
rect 13648 19556 13652 19612
rect 13652 19556 13708 19612
rect 13708 19556 13712 19612
rect 13648 19552 13712 19556
rect 13728 19612 13792 19616
rect 13728 19556 13732 19612
rect 13732 19556 13788 19612
rect 13788 19556 13792 19612
rect 13728 19552 13792 19556
rect 13808 19612 13872 19616
rect 13808 19556 13812 19612
rect 13812 19556 13868 19612
rect 13868 19556 13872 19612
rect 13808 19552 13872 19556
rect 13888 19612 13952 19616
rect 13888 19556 13892 19612
rect 13892 19556 13948 19612
rect 13948 19556 13952 19612
rect 13888 19552 13952 19556
rect 19996 19612 20060 19616
rect 19996 19556 20000 19612
rect 20000 19556 20056 19612
rect 20056 19556 20060 19612
rect 19996 19552 20060 19556
rect 20076 19612 20140 19616
rect 20076 19556 20080 19612
rect 20080 19556 20136 19612
rect 20136 19556 20140 19612
rect 20076 19552 20140 19556
rect 20156 19612 20220 19616
rect 20156 19556 20160 19612
rect 20160 19556 20216 19612
rect 20216 19556 20220 19612
rect 20156 19552 20220 19556
rect 20236 19612 20300 19616
rect 20236 19556 20240 19612
rect 20240 19556 20296 19612
rect 20296 19556 20300 19612
rect 20236 19552 20300 19556
rect 26344 19612 26408 19616
rect 26344 19556 26348 19612
rect 26348 19556 26404 19612
rect 26404 19556 26408 19612
rect 26344 19552 26408 19556
rect 26424 19612 26488 19616
rect 26424 19556 26428 19612
rect 26428 19556 26484 19612
rect 26484 19556 26488 19612
rect 26424 19552 26488 19556
rect 26504 19612 26568 19616
rect 26504 19556 26508 19612
rect 26508 19556 26564 19612
rect 26564 19556 26568 19612
rect 26504 19552 26568 19556
rect 26584 19612 26648 19616
rect 26584 19556 26588 19612
rect 26588 19556 26644 19612
rect 26644 19556 26648 19612
rect 26584 19552 26648 19556
rect 4126 19068 4190 19072
rect 4126 19012 4130 19068
rect 4130 19012 4186 19068
rect 4186 19012 4190 19068
rect 4126 19008 4190 19012
rect 4206 19068 4270 19072
rect 4206 19012 4210 19068
rect 4210 19012 4266 19068
rect 4266 19012 4270 19068
rect 4206 19008 4270 19012
rect 4286 19068 4350 19072
rect 4286 19012 4290 19068
rect 4290 19012 4346 19068
rect 4346 19012 4350 19068
rect 4286 19008 4350 19012
rect 4366 19068 4430 19072
rect 4366 19012 4370 19068
rect 4370 19012 4426 19068
rect 4426 19012 4430 19068
rect 4366 19008 4430 19012
rect 10474 19068 10538 19072
rect 10474 19012 10478 19068
rect 10478 19012 10534 19068
rect 10534 19012 10538 19068
rect 10474 19008 10538 19012
rect 10554 19068 10618 19072
rect 10554 19012 10558 19068
rect 10558 19012 10614 19068
rect 10614 19012 10618 19068
rect 10554 19008 10618 19012
rect 10634 19068 10698 19072
rect 10634 19012 10638 19068
rect 10638 19012 10694 19068
rect 10694 19012 10698 19068
rect 10634 19008 10698 19012
rect 10714 19068 10778 19072
rect 10714 19012 10718 19068
rect 10718 19012 10774 19068
rect 10774 19012 10778 19068
rect 10714 19008 10778 19012
rect 16822 19068 16886 19072
rect 16822 19012 16826 19068
rect 16826 19012 16882 19068
rect 16882 19012 16886 19068
rect 16822 19008 16886 19012
rect 16902 19068 16966 19072
rect 16902 19012 16906 19068
rect 16906 19012 16962 19068
rect 16962 19012 16966 19068
rect 16902 19008 16966 19012
rect 16982 19068 17046 19072
rect 16982 19012 16986 19068
rect 16986 19012 17042 19068
rect 17042 19012 17046 19068
rect 16982 19008 17046 19012
rect 17062 19068 17126 19072
rect 17062 19012 17066 19068
rect 17066 19012 17122 19068
rect 17122 19012 17126 19068
rect 17062 19008 17126 19012
rect 23170 19068 23234 19072
rect 23170 19012 23174 19068
rect 23174 19012 23230 19068
rect 23230 19012 23234 19068
rect 23170 19008 23234 19012
rect 23250 19068 23314 19072
rect 23250 19012 23254 19068
rect 23254 19012 23310 19068
rect 23310 19012 23314 19068
rect 23250 19008 23314 19012
rect 23330 19068 23394 19072
rect 23330 19012 23334 19068
rect 23334 19012 23390 19068
rect 23390 19012 23394 19068
rect 23330 19008 23394 19012
rect 23410 19068 23474 19072
rect 23410 19012 23414 19068
rect 23414 19012 23470 19068
rect 23470 19012 23474 19068
rect 23410 19008 23474 19012
rect 7300 18524 7364 18528
rect 7300 18468 7304 18524
rect 7304 18468 7360 18524
rect 7360 18468 7364 18524
rect 7300 18464 7364 18468
rect 7380 18524 7444 18528
rect 7380 18468 7384 18524
rect 7384 18468 7440 18524
rect 7440 18468 7444 18524
rect 7380 18464 7444 18468
rect 7460 18524 7524 18528
rect 7460 18468 7464 18524
rect 7464 18468 7520 18524
rect 7520 18468 7524 18524
rect 7460 18464 7524 18468
rect 7540 18524 7604 18528
rect 7540 18468 7544 18524
rect 7544 18468 7600 18524
rect 7600 18468 7604 18524
rect 7540 18464 7604 18468
rect 13648 18524 13712 18528
rect 13648 18468 13652 18524
rect 13652 18468 13708 18524
rect 13708 18468 13712 18524
rect 13648 18464 13712 18468
rect 13728 18524 13792 18528
rect 13728 18468 13732 18524
rect 13732 18468 13788 18524
rect 13788 18468 13792 18524
rect 13728 18464 13792 18468
rect 13808 18524 13872 18528
rect 13808 18468 13812 18524
rect 13812 18468 13868 18524
rect 13868 18468 13872 18524
rect 13808 18464 13872 18468
rect 13888 18524 13952 18528
rect 13888 18468 13892 18524
rect 13892 18468 13948 18524
rect 13948 18468 13952 18524
rect 13888 18464 13952 18468
rect 19996 18524 20060 18528
rect 19996 18468 20000 18524
rect 20000 18468 20056 18524
rect 20056 18468 20060 18524
rect 19996 18464 20060 18468
rect 20076 18524 20140 18528
rect 20076 18468 20080 18524
rect 20080 18468 20136 18524
rect 20136 18468 20140 18524
rect 20076 18464 20140 18468
rect 20156 18524 20220 18528
rect 20156 18468 20160 18524
rect 20160 18468 20216 18524
rect 20216 18468 20220 18524
rect 20156 18464 20220 18468
rect 20236 18524 20300 18528
rect 20236 18468 20240 18524
rect 20240 18468 20296 18524
rect 20296 18468 20300 18524
rect 20236 18464 20300 18468
rect 26344 18524 26408 18528
rect 26344 18468 26348 18524
rect 26348 18468 26404 18524
rect 26404 18468 26408 18524
rect 26344 18464 26408 18468
rect 26424 18524 26488 18528
rect 26424 18468 26428 18524
rect 26428 18468 26484 18524
rect 26484 18468 26488 18524
rect 26424 18464 26488 18468
rect 26504 18524 26568 18528
rect 26504 18468 26508 18524
rect 26508 18468 26564 18524
rect 26564 18468 26568 18524
rect 26504 18464 26568 18468
rect 26584 18524 26648 18528
rect 26584 18468 26588 18524
rect 26588 18468 26644 18524
rect 26644 18468 26648 18524
rect 26584 18464 26648 18468
rect 4126 17980 4190 17984
rect 4126 17924 4130 17980
rect 4130 17924 4186 17980
rect 4186 17924 4190 17980
rect 4126 17920 4190 17924
rect 4206 17980 4270 17984
rect 4206 17924 4210 17980
rect 4210 17924 4266 17980
rect 4266 17924 4270 17980
rect 4206 17920 4270 17924
rect 4286 17980 4350 17984
rect 4286 17924 4290 17980
rect 4290 17924 4346 17980
rect 4346 17924 4350 17980
rect 4286 17920 4350 17924
rect 4366 17980 4430 17984
rect 4366 17924 4370 17980
rect 4370 17924 4426 17980
rect 4426 17924 4430 17980
rect 4366 17920 4430 17924
rect 10474 17980 10538 17984
rect 10474 17924 10478 17980
rect 10478 17924 10534 17980
rect 10534 17924 10538 17980
rect 10474 17920 10538 17924
rect 10554 17980 10618 17984
rect 10554 17924 10558 17980
rect 10558 17924 10614 17980
rect 10614 17924 10618 17980
rect 10554 17920 10618 17924
rect 10634 17980 10698 17984
rect 10634 17924 10638 17980
rect 10638 17924 10694 17980
rect 10694 17924 10698 17980
rect 10634 17920 10698 17924
rect 10714 17980 10778 17984
rect 10714 17924 10718 17980
rect 10718 17924 10774 17980
rect 10774 17924 10778 17980
rect 10714 17920 10778 17924
rect 16822 17980 16886 17984
rect 16822 17924 16826 17980
rect 16826 17924 16882 17980
rect 16882 17924 16886 17980
rect 16822 17920 16886 17924
rect 16902 17980 16966 17984
rect 16902 17924 16906 17980
rect 16906 17924 16962 17980
rect 16962 17924 16966 17980
rect 16902 17920 16966 17924
rect 16982 17980 17046 17984
rect 16982 17924 16986 17980
rect 16986 17924 17042 17980
rect 17042 17924 17046 17980
rect 16982 17920 17046 17924
rect 17062 17980 17126 17984
rect 17062 17924 17066 17980
rect 17066 17924 17122 17980
rect 17122 17924 17126 17980
rect 17062 17920 17126 17924
rect 23170 17980 23234 17984
rect 23170 17924 23174 17980
rect 23174 17924 23230 17980
rect 23230 17924 23234 17980
rect 23170 17920 23234 17924
rect 23250 17980 23314 17984
rect 23250 17924 23254 17980
rect 23254 17924 23310 17980
rect 23310 17924 23314 17980
rect 23250 17920 23314 17924
rect 23330 17980 23394 17984
rect 23330 17924 23334 17980
rect 23334 17924 23390 17980
rect 23390 17924 23394 17980
rect 23330 17920 23394 17924
rect 23410 17980 23474 17984
rect 23410 17924 23414 17980
rect 23414 17924 23470 17980
rect 23470 17924 23474 17980
rect 23410 17920 23474 17924
rect 7300 17436 7364 17440
rect 7300 17380 7304 17436
rect 7304 17380 7360 17436
rect 7360 17380 7364 17436
rect 7300 17376 7364 17380
rect 7380 17436 7444 17440
rect 7380 17380 7384 17436
rect 7384 17380 7440 17436
rect 7440 17380 7444 17436
rect 7380 17376 7444 17380
rect 7460 17436 7524 17440
rect 7460 17380 7464 17436
rect 7464 17380 7520 17436
rect 7520 17380 7524 17436
rect 7460 17376 7524 17380
rect 7540 17436 7604 17440
rect 7540 17380 7544 17436
rect 7544 17380 7600 17436
rect 7600 17380 7604 17436
rect 7540 17376 7604 17380
rect 13648 17436 13712 17440
rect 13648 17380 13652 17436
rect 13652 17380 13708 17436
rect 13708 17380 13712 17436
rect 13648 17376 13712 17380
rect 13728 17436 13792 17440
rect 13728 17380 13732 17436
rect 13732 17380 13788 17436
rect 13788 17380 13792 17436
rect 13728 17376 13792 17380
rect 13808 17436 13872 17440
rect 13808 17380 13812 17436
rect 13812 17380 13868 17436
rect 13868 17380 13872 17436
rect 13808 17376 13872 17380
rect 13888 17436 13952 17440
rect 13888 17380 13892 17436
rect 13892 17380 13948 17436
rect 13948 17380 13952 17436
rect 13888 17376 13952 17380
rect 19996 17436 20060 17440
rect 19996 17380 20000 17436
rect 20000 17380 20056 17436
rect 20056 17380 20060 17436
rect 19996 17376 20060 17380
rect 20076 17436 20140 17440
rect 20076 17380 20080 17436
rect 20080 17380 20136 17436
rect 20136 17380 20140 17436
rect 20076 17376 20140 17380
rect 20156 17436 20220 17440
rect 20156 17380 20160 17436
rect 20160 17380 20216 17436
rect 20216 17380 20220 17436
rect 20156 17376 20220 17380
rect 20236 17436 20300 17440
rect 20236 17380 20240 17436
rect 20240 17380 20296 17436
rect 20296 17380 20300 17436
rect 20236 17376 20300 17380
rect 26344 17436 26408 17440
rect 26344 17380 26348 17436
rect 26348 17380 26404 17436
rect 26404 17380 26408 17436
rect 26344 17376 26408 17380
rect 26424 17436 26488 17440
rect 26424 17380 26428 17436
rect 26428 17380 26484 17436
rect 26484 17380 26488 17436
rect 26424 17376 26488 17380
rect 26504 17436 26568 17440
rect 26504 17380 26508 17436
rect 26508 17380 26564 17436
rect 26564 17380 26568 17436
rect 26504 17376 26568 17380
rect 26584 17436 26648 17440
rect 26584 17380 26588 17436
rect 26588 17380 26644 17436
rect 26644 17380 26648 17436
rect 26584 17376 26648 17380
rect 4126 16892 4190 16896
rect 4126 16836 4130 16892
rect 4130 16836 4186 16892
rect 4186 16836 4190 16892
rect 4126 16832 4190 16836
rect 4206 16892 4270 16896
rect 4206 16836 4210 16892
rect 4210 16836 4266 16892
rect 4266 16836 4270 16892
rect 4206 16832 4270 16836
rect 4286 16892 4350 16896
rect 4286 16836 4290 16892
rect 4290 16836 4346 16892
rect 4346 16836 4350 16892
rect 4286 16832 4350 16836
rect 4366 16892 4430 16896
rect 4366 16836 4370 16892
rect 4370 16836 4426 16892
rect 4426 16836 4430 16892
rect 4366 16832 4430 16836
rect 10474 16892 10538 16896
rect 10474 16836 10478 16892
rect 10478 16836 10534 16892
rect 10534 16836 10538 16892
rect 10474 16832 10538 16836
rect 10554 16892 10618 16896
rect 10554 16836 10558 16892
rect 10558 16836 10614 16892
rect 10614 16836 10618 16892
rect 10554 16832 10618 16836
rect 10634 16892 10698 16896
rect 10634 16836 10638 16892
rect 10638 16836 10694 16892
rect 10694 16836 10698 16892
rect 10634 16832 10698 16836
rect 10714 16892 10778 16896
rect 10714 16836 10718 16892
rect 10718 16836 10774 16892
rect 10774 16836 10778 16892
rect 10714 16832 10778 16836
rect 16822 16892 16886 16896
rect 16822 16836 16826 16892
rect 16826 16836 16882 16892
rect 16882 16836 16886 16892
rect 16822 16832 16886 16836
rect 16902 16892 16966 16896
rect 16902 16836 16906 16892
rect 16906 16836 16962 16892
rect 16962 16836 16966 16892
rect 16902 16832 16966 16836
rect 16982 16892 17046 16896
rect 16982 16836 16986 16892
rect 16986 16836 17042 16892
rect 17042 16836 17046 16892
rect 16982 16832 17046 16836
rect 17062 16892 17126 16896
rect 17062 16836 17066 16892
rect 17066 16836 17122 16892
rect 17122 16836 17126 16892
rect 17062 16832 17126 16836
rect 23170 16892 23234 16896
rect 23170 16836 23174 16892
rect 23174 16836 23230 16892
rect 23230 16836 23234 16892
rect 23170 16832 23234 16836
rect 23250 16892 23314 16896
rect 23250 16836 23254 16892
rect 23254 16836 23310 16892
rect 23310 16836 23314 16892
rect 23250 16832 23314 16836
rect 23330 16892 23394 16896
rect 23330 16836 23334 16892
rect 23334 16836 23390 16892
rect 23390 16836 23394 16892
rect 23330 16832 23394 16836
rect 23410 16892 23474 16896
rect 23410 16836 23414 16892
rect 23414 16836 23470 16892
rect 23470 16836 23474 16892
rect 23410 16832 23474 16836
rect 7300 16348 7364 16352
rect 7300 16292 7304 16348
rect 7304 16292 7360 16348
rect 7360 16292 7364 16348
rect 7300 16288 7364 16292
rect 7380 16348 7444 16352
rect 7380 16292 7384 16348
rect 7384 16292 7440 16348
rect 7440 16292 7444 16348
rect 7380 16288 7444 16292
rect 7460 16348 7524 16352
rect 7460 16292 7464 16348
rect 7464 16292 7520 16348
rect 7520 16292 7524 16348
rect 7460 16288 7524 16292
rect 7540 16348 7604 16352
rect 7540 16292 7544 16348
rect 7544 16292 7600 16348
rect 7600 16292 7604 16348
rect 7540 16288 7604 16292
rect 13648 16348 13712 16352
rect 13648 16292 13652 16348
rect 13652 16292 13708 16348
rect 13708 16292 13712 16348
rect 13648 16288 13712 16292
rect 13728 16348 13792 16352
rect 13728 16292 13732 16348
rect 13732 16292 13788 16348
rect 13788 16292 13792 16348
rect 13728 16288 13792 16292
rect 13808 16348 13872 16352
rect 13808 16292 13812 16348
rect 13812 16292 13868 16348
rect 13868 16292 13872 16348
rect 13808 16288 13872 16292
rect 13888 16348 13952 16352
rect 13888 16292 13892 16348
rect 13892 16292 13948 16348
rect 13948 16292 13952 16348
rect 13888 16288 13952 16292
rect 19996 16348 20060 16352
rect 19996 16292 20000 16348
rect 20000 16292 20056 16348
rect 20056 16292 20060 16348
rect 19996 16288 20060 16292
rect 20076 16348 20140 16352
rect 20076 16292 20080 16348
rect 20080 16292 20136 16348
rect 20136 16292 20140 16348
rect 20076 16288 20140 16292
rect 20156 16348 20220 16352
rect 20156 16292 20160 16348
rect 20160 16292 20216 16348
rect 20216 16292 20220 16348
rect 20156 16288 20220 16292
rect 20236 16348 20300 16352
rect 20236 16292 20240 16348
rect 20240 16292 20296 16348
rect 20296 16292 20300 16348
rect 20236 16288 20300 16292
rect 26344 16348 26408 16352
rect 26344 16292 26348 16348
rect 26348 16292 26404 16348
rect 26404 16292 26408 16348
rect 26344 16288 26408 16292
rect 26424 16348 26488 16352
rect 26424 16292 26428 16348
rect 26428 16292 26484 16348
rect 26484 16292 26488 16348
rect 26424 16288 26488 16292
rect 26504 16348 26568 16352
rect 26504 16292 26508 16348
rect 26508 16292 26564 16348
rect 26564 16292 26568 16348
rect 26504 16288 26568 16292
rect 26584 16348 26648 16352
rect 26584 16292 26588 16348
rect 26588 16292 26644 16348
rect 26644 16292 26648 16348
rect 26584 16288 26648 16292
rect 4126 15804 4190 15808
rect 4126 15748 4130 15804
rect 4130 15748 4186 15804
rect 4186 15748 4190 15804
rect 4126 15744 4190 15748
rect 4206 15804 4270 15808
rect 4206 15748 4210 15804
rect 4210 15748 4266 15804
rect 4266 15748 4270 15804
rect 4206 15744 4270 15748
rect 4286 15804 4350 15808
rect 4286 15748 4290 15804
rect 4290 15748 4346 15804
rect 4346 15748 4350 15804
rect 4286 15744 4350 15748
rect 4366 15804 4430 15808
rect 4366 15748 4370 15804
rect 4370 15748 4426 15804
rect 4426 15748 4430 15804
rect 4366 15744 4430 15748
rect 10474 15804 10538 15808
rect 10474 15748 10478 15804
rect 10478 15748 10534 15804
rect 10534 15748 10538 15804
rect 10474 15744 10538 15748
rect 10554 15804 10618 15808
rect 10554 15748 10558 15804
rect 10558 15748 10614 15804
rect 10614 15748 10618 15804
rect 10554 15744 10618 15748
rect 10634 15804 10698 15808
rect 10634 15748 10638 15804
rect 10638 15748 10694 15804
rect 10694 15748 10698 15804
rect 10634 15744 10698 15748
rect 10714 15804 10778 15808
rect 10714 15748 10718 15804
rect 10718 15748 10774 15804
rect 10774 15748 10778 15804
rect 10714 15744 10778 15748
rect 16822 15804 16886 15808
rect 16822 15748 16826 15804
rect 16826 15748 16882 15804
rect 16882 15748 16886 15804
rect 16822 15744 16886 15748
rect 16902 15804 16966 15808
rect 16902 15748 16906 15804
rect 16906 15748 16962 15804
rect 16962 15748 16966 15804
rect 16902 15744 16966 15748
rect 16982 15804 17046 15808
rect 16982 15748 16986 15804
rect 16986 15748 17042 15804
rect 17042 15748 17046 15804
rect 16982 15744 17046 15748
rect 17062 15804 17126 15808
rect 17062 15748 17066 15804
rect 17066 15748 17122 15804
rect 17122 15748 17126 15804
rect 17062 15744 17126 15748
rect 23170 15804 23234 15808
rect 23170 15748 23174 15804
rect 23174 15748 23230 15804
rect 23230 15748 23234 15804
rect 23170 15744 23234 15748
rect 23250 15804 23314 15808
rect 23250 15748 23254 15804
rect 23254 15748 23310 15804
rect 23310 15748 23314 15804
rect 23250 15744 23314 15748
rect 23330 15804 23394 15808
rect 23330 15748 23334 15804
rect 23334 15748 23390 15804
rect 23390 15748 23394 15804
rect 23330 15744 23394 15748
rect 23410 15804 23474 15808
rect 23410 15748 23414 15804
rect 23414 15748 23470 15804
rect 23470 15748 23474 15804
rect 23410 15744 23474 15748
rect 7300 15260 7364 15264
rect 7300 15204 7304 15260
rect 7304 15204 7360 15260
rect 7360 15204 7364 15260
rect 7300 15200 7364 15204
rect 7380 15260 7444 15264
rect 7380 15204 7384 15260
rect 7384 15204 7440 15260
rect 7440 15204 7444 15260
rect 7380 15200 7444 15204
rect 7460 15260 7524 15264
rect 7460 15204 7464 15260
rect 7464 15204 7520 15260
rect 7520 15204 7524 15260
rect 7460 15200 7524 15204
rect 7540 15260 7604 15264
rect 7540 15204 7544 15260
rect 7544 15204 7600 15260
rect 7600 15204 7604 15260
rect 7540 15200 7604 15204
rect 13648 15260 13712 15264
rect 13648 15204 13652 15260
rect 13652 15204 13708 15260
rect 13708 15204 13712 15260
rect 13648 15200 13712 15204
rect 13728 15260 13792 15264
rect 13728 15204 13732 15260
rect 13732 15204 13788 15260
rect 13788 15204 13792 15260
rect 13728 15200 13792 15204
rect 13808 15260 13872 15264
rect 13808 15204 13812 15260
rect 13812 15204 13868 15260
rect 13868 15204 13872 15260
rect 13808 15200 13872 15204
rect 13888 15260 13952 15264
rect 13888 15204 13892 15260
rect 13892 15204 13948 15260
rect 13948 15204 13952 15260
rect 13888 15200 13952 15204
rect 19996 15260 20060 15264
rect 19996 15204 20000 15260
rect 20000 15204 20056 15260
rect 20056 15204 20060 15260
rect 19996 15200 20060 15204
rect 20076 15260 20140 15264
rect 20076 15204 20080 15260
rect 20080 15204 20136 15260
rect 20136 15204 20140 15260
rect 20076 15200 20140 15204
rect 20156 15260 20220 15264
rect 20156 15204 20160 15260
rect 20160 15204 20216 15260
rect 20216 15204 20220 15260
rect 20156 15200 20220 15204
rect 20236 15260 20300 15264
rect 20236 15204 20240 15260
rect 20240 15204 20296 15260
rect 20296 15204 20300 15260
rect 20236 15200 20300 15204
rect 26344 15260 26408 15264
rect 26344 15204 26348 15260
rect 26348 15204 26404 15260
rect 26404 15204 26408 15260
rect 26344 15200 26408 15204
rect 26424 15260 26488 15264
rect 26424 15204 26428 15260
rect 26428 15204 26484 15260
rect 26484 15204 26488 15260
rect 26424 15200 26488 15204
rect 26504 15260 26568 15264
rect 26504 15204 26508 15260
rect 26508 15204 26564 15260
rect 26564 15204 26568 15260
rect 26504 15200 26568 15204
rect 26584 15260 26648 15264
rect 26584 15204 26588 15260
rect 26588 15204 26644 15260
rect 26644 15204 26648 15260
rect 26584 15200 26648 15204
rect 4126 14716 4190 14720
rect 4126 14660 4130 14716
rect 4130 14660 4186 14716
rect 4186 14660 4190 14716
rect 4126 14656 4190 14660
rect 4206 14716 4270 14720
rect 4206 14660 4210 14716
rect 4210 14660 4266 14716
rect 4266 14660 4270 14716
rect 4206 14656 4270 14660
rect 4286 14716 4350 14720
rect 4286 14660 4290 14716
rect 4290 14660 4346 14716
rect 4346 14660 4350 14716
rect 4286 14656 4350 14660
rect 4366 14716 4430 14720
rect 4366 14660 4370 14716
rect 4370 14660 4426 14716
rect 4426 14660 4430 14716
rect 4366 14656 4430 14660
rect 10474 14716 10538 14720
rect 10474 14660 10478 14716
rect 10478 14660 10534 14716
rect 10534 14660 10538 14716
rect 10474 14656 10538 14660
rect 10554 14716 10618 14720
rect 10554 14660 10558 14716
rect 10558 14660 10614 14716
rect 10614 14660 10618 14716
rect 10554 14656 10618 14660
rect 10634 14716 10698 14720
rect 10634 14660 10638 14716
rect 10638 14660 10694 14716
rect 10694 14660 10698 14716
rect 10634 14656 10698 14660
rect 10714 14716 10778 14720
rect 10714 14660 10718 14716
rect 10718 14660 10774 14716
rect 10774 14660 10778 14716
rect 10714 14656 10778 14660
rect 16822 14716 16886 14720
rect 16822 14660 16826 14716
rect 16826 14660 16882 14716
rect 16882 14660 16886 14716
rect 16822 14656 16886 14660
rect 16902 14716 16966 14720
rect 16902 14660 16906 14716
rect 16906 14660 16962 14716
rect 16962 14660 16966 14716
rect 16902 14656 16966 14660
rect 16982 14716 17046 14720
rect 16982 14660 16986 14716
rect 16986 14660 17042 14716
rect 17042 14660 17046 14716
rect 16982 14656 17046 14660
rect 17062 14716 17126 14720
rect 17062 14660 17066 14716
rect 17066 14660 17122 14716
rect 17122 14660 17126 14716
rect 17062 14656 17126 14660
rect 23170 14716 23234 14720
rect 23170 14660 23174 14716
rect 23174 14660 23230 14716
rect 23230 14660 23234 14716
rect 23170 14656 23234 14660
rect 23250 14716 23314 14720
rect 23250 14660 23254 14716
rect 23254 14660 23310 14716
rect 23310 14660 23314 14716
rect 23250 14656 23314 14660
rect 23330 14716 23394 14720
rect 23330 14660 23334 14716
rect 23334 14660 23390 14716
rect 23390 14660 23394 14716
rect 23330 14656 23394 14660
rect 23410 14716 23474 14720
rect 23410 14660 23414 14716
rect 23414 14660 23470 14716
rect 23470 14660 23474 14716
rect 23410 14656 23474 14660
rect 7300 14172 7364 14176
rect 7300 14116 7304 14172
rect 7304 14116 7360 14172
rect 7360 14116 7364 14172
rect 7300 14112 7364 14116
rect 7380 14172 7444 14176
rect 7380 14116 7384 14172
rect 7384 14116 7440 14172
rect 7440 14116 7444 14172
rect 7380 14112 7444 14116
rect 7460 14172 7524 14176
rect 7460 14116 7464 14172
rect 7464 14116 7520 14172
rect 7520 14116 7524 14172
rect 7460 14112 7524 14116
rect 7540 14172 7604 14176
rect 7540 14116 7544 14172
rect 7544 14116 7600 14172
rect 7600 14116 7604 14172
rect 7540 14112 7604 14116
rect 13648 14172 13712 14176
rect 13648 14116 13652 14172
rect 13652 14116 13708 14172
rect 13708 14116 13712 14172
rect 13648 14112 13712 14116
rect 13728 14172 13792 14176
rect 13728 14116 13732 14172
rect 13732 14116 13788 14172
rect 13788 14116 13792 14172
rect 13728 14112 13792 14116
rect 13808 14172 13872 14176
rect 13808 14116 13812 14172
rect 13812 14116 13868 14172
rect 13868 14116 13872 14172
rect 13808 14112 13872 14116
rect 13888 14172 13952 14176
rect 13888 14116 13892 14172
rect 13892 14116 13948 14172
rect 13948 14116 13952 14172
rect 13888 14112 13952 14116
rect 19996 14172 20060 14176
rect 19996 14116 20000 14172
rect 20000 14116 20056 14172
rect 20056 14116 20060 14172
rect 19996 14112 20060 14116
rect 20076 14172 20140 14176
rect 20076 14116 20080 14172
rect 20080 14116 20136 14172
rect 20136 14116 20140 14172
rect 20076 14112 20140 14116
rect 20156 14172 20220 14176
rect 20156 14116 20160 14172
rect 20160 14116 20216 14172
rect 20216 14116 20220 14172
rect 20156 14112 20220 14116
rect 20236 14172 20300 14176
rect 20236 14116 20240 14172
rect 20240 14116 20296 14172
rect 20296 14116 20300 14172
rect 20236 14112 20300 14116
rect 26344 14172 26408 14176
rect 26344 14116 26348 14172
rect 26348 14116 26404 14172
rect 26404 14116 26408 14172
rect 26344 14112 26408 14116
rect 26424 14172 26488 14176
rect 26424 14116 26428 14172
rect 26428 14116 26484 14172
rect 26484 14116 26488 14172
rect 26424 14112 26488 14116
rect 26504 14172 26568 14176
rect 26504 14116 26508 14172
rect 26508 14116 26564 14172
rect 26564 14116 26568 14172
rect 26504 14112 26568 14116
rect 26584 14172 26648 14176
rect 26584 14116 26588 14172
rect 26588 14116 26644 14172
rect 26644 14116 26648 14172
rect 26584 14112 26648 14116
rect 4126 13628 4190 13632
rect 4126 13572 4130 13628
rect 4130 13572 4186 13628
rect 4186 13572 4190 13628
rect 4126 13568 4190 13572
rect 4206 13628 4270 13632
rect 4206 13572 4210 13628
rect 4210 13572 4266 13628
rect 4266 13572 4270 13628
rect 4206 13568 4270 13572
rect 4286 13628 4350 13632
rect 4286 13572 4290 13628
rect 4290 13572 4346 13628
rect 4346 13572 4350 13628
rect 4286 13568 4350 13572
rect 4366 13628 4430 13632
rect 4366 13572 4370 13628
rect 4370 13572 4426 13628
rect 4426 13572 4430 13628
rect 4366 13568 4430 13572
rect 10474 13628 10538 13632
rect 10474 13572 10478 13628
rect 10478 13572 10534 13628
rect 10534 13572 10538 13628
rect 10474 13568 10538 13572
rect 10554 13628 10618 13632
rect 10554 13572 10558 13628
rect 10558 13572 10614 13628
rect 10614 13572 10618 13628
rect 10554 13568 10618 13572
rect 10634 13628 10698 13632
rect 10634 13572 10638 13628
rect 10638 13572 10694 13628
rect 10694 13572 10698 13628
rect 10634 13568 10698 13572
rect 10714 13628 10778 13632
rect 10714 13572 10718 13628
rect 10718 13572 10774 13628
rect 10774 13572 10778 13628
rect 10714 13568 10778 13572
rect 16822 13628 16886 13632
rect 16822 13572 16826 13628
rect 16826 13572 16882 13628
rect 16882 13572 16886 13628
rect 16822 13568 16886 13572
rect 16902 13628 16966 13632
rect 16902 13572 16906 13628
rect 16906 13572 16962 13628
rect 16962 13572 16966 13628
rect 16902 13568 16966 13572
rect 16982 13628 17046 13632
rect 16982 13572 16986 13628
rect 16986 13572 17042 13628
rect 17042 13572 17046 13628
rect 16982 13568 17046 13572
rect 17062 13628 17126 13632
rect 17062 13572 17066 13628
rect 17066 13572 17122 13628
rect 17122 13572 17126 13628
rect 17062 13568 17126 13572
rect 23170 13628 23234 13632
rect 23170 13572 23174 13628
rect 23174 13572 23230 13628
rect 23230 13572 23234 13628
rect 23170 13568 23234 13572
rect 23250 13628 23314 13632
rect 23250 13572 23254 13628
rect 23254 13572 23310 13628
rect 23310 13572 23314 13628
rect 23250 13568 23314 13572
rect 23330 13628 23394 13632
rect 23330 13572 23334 13628
rect 23334 13572 23390 13628
rect 23390 13572 23394 13628
rect 23330 13568 23394 13572
rect 23410 13628 23474 13632
rect 23410 13572 23414 13628
rect 23414 13572 23470 13628
rect 23470 13572 23474 13628
rect 23410 13568 23474 13572
rect 7300 13084 7364 13088
rect 7300 13028 7304 13084
rect 7304 13028 7360 13084
rect 7360 13028 7364 13084
rect 7300 13024 7364 13028
rect 7380 13084 7444 13088
rect 7380 13028 7384 13084
rect 7384 13028 7440 13084
rect 7440 13028 7444 13084
rect 7380 13024 7444 13028
rect 7460 13084 7524 13088
rect 7460 13028 7464 13084
rect 7464 13028 7520 13084
rect 7520 13028 7524 13084
rect 7460 13024 7524 13028
rect 7540 13084 7604 13088
rect 7540 13028 7544 13084
rect 7544 13028 7600 13084
rect 7600 13028 7604 13084
rect 7540 13024 7604 13028
rect 13648 13084 13712 13088
rect 13648 13028 13652 13084
rect 13652 13028 13708 13084
rect 13708 13028 13712 13084
rect 13648 13024 13712 13028
rect 13728 13084 13792 13088
rect 13728 13028 13732 13084
rect 13732 13028 13788 13084
rect 13788 13028 13792 13084
rect 13728 13024 13792 13028
rect 13808 13084 13872 13088
rect 13808 13028 13812 13084
rect 13812 13028 13868 13084
rect 13868 13028 13872 13084
rect 13808 13024 13872 13028
rect 13888 13084 13952 13088
rect 13888 13028 13892 13084
rect 13892 13028 13948 13084
rect 13948 13028 13952 13084
rect 13888 13024 13952 13028
rect 19996 13084 20060 13088
rect 19996 13028 20000 13084
rect 20000 13028 20056 13084
rect 20056 13028 20060 13084
rect 19996 13024 20060 13028
rect 20076 13084 20140 13088
rect 20076 13028 20080 13084
rect 20080 13028 20136 13084
rect 20136 13028 20140 13084
rect 20076 13024 20140 13028
rect 20156 13084 20220 13088
rect 20156 13028 20160 13084
rect 20160 13028 20216 13084
rect 20216 13028 20220 13084
rect 20156 13024 20220 13028
rect 20236 13084 20300 13088
rect 20236 13028 20240 13084
rect 20240 13028 20296 13084
rect 20296 13028 20300 13084
rect 20236 13024 20300 13028
rect 26344 13084 26408 13088
rect 26344 13028 26348 13084
rect 26348 13028 26404 13084
rect 26404 13028 26408 13084
rect 26344 13024 26408 13028
rect 26424 13084 26488 13088
rect 26424 13028 26428 13084
rect 26428 13028 26484 13084
rect 26484 13028 26488 13084
rect 26424 13024 26488 13028
rect 26504 13084 26568 13088
rect 26504 13028 26508 13084
rect 26508 13028 26564 13084
rect 26564 13028 26568 13084
rect 26504 13024 26568 13028
rect 26584 13084 26648 13088
rect 26584 13028 26588 13084
rect 26588 13028 26644 13084
rect 26644 13028 26648 13084
rect 26584 13024 26648 13028
rect 4126 12540 4190 12544
rect 4126 12484 4130 12540
rect 4130 12484 4186 12540
rect 4186 12484 4190 12540
rect 4126 12480 4190 12484
rect 4206 12540 4270 12544
rect 4206 12484 4210 12540
rect 4210 12484 4266 12540
rect 4266 12484 4270 12540
rect 4206 12480 4270 12484
rect 4286 12540 4350 12544
rect 4286 12484 4290 12540
rect 4290 12484 4346 12540
rect 4346 12484 4350 12540
rect 4286 12480 4350 12484
rect 4366 12540 4430 12544
rect 4366 12484 4370 12540
rect 4370 12484 4426 12540
rect 4426 12484 4430 12540
rect 4366 12480 4430 12484
rect 10474 12540 10538 12544
rect 10474 12484 10478 12540
rect 10478 12484 10534 12540
rect 10534 12484 10538 12540
rect 10474 12480 10538 12484
rect 10554 12540 10618 12544
rect 10554 12484 10558 12540
rect 10558 12484 10614 12540
rect 10614 12484 10618 12540
rect 10554 12480 10618 12484
rect 10634 12540 10698 12544
rect 10634 12484 10638 12540
rect 10638 12484 10694 12540
rect 10694 12484 10698 12540
rect 10634 12480 10698 12484
rect 10714 12540 10778 12544
rect 10714 12484 10718 12540
rect 10718 12484 10774 12540
rect 10774 12484 10778 12540
rect 10714 12480 10778 12484
rect 16822 12540 16886 12544
rect 16822 12484 16826 12540
rect 16826 12484 16882 12540
rect 16882 12484 16886 12540
rect 16822 12480 16886 12484
rect 16902 12540 16966 12544
rect 16902 12484 16906 12540
rect 16906 12484 16962 12540
rect 16962 12484 16966 12540
rect 16902 12480 16966 12484
rect 16982 12540 17046 12544
rect 16982 12484 16986 12540
rect 16986 12484 17042 12540
rect 17042 12484 17046 12540
rect 16982 12480 17046 12484
rect 17062 12540 17126 12544
rect 17062 12484 17066 12540
rect 17066 12484 17122 12540
rect 17122 12484 17126 12540
rect 17062 12480 17126 12484
rect 23170 12540 23234 12544
rect 23170 12484 23174 12540
rect 23174 12484 23230 12540
rect 23230 12484 23234 12540
rect 23170 12480 23234 12484
rect 23250 12540 23314 12544
rect 23250 12484 23254 12540
rect 23254 12484 23310 12540
rect 23310 12484 23314 12540
rect 23250 12480 23314 12484
rect 23330 12540 23394 12544
rect 23330 12484 23334 12540
rect 23334 12484 23390 12540
rect 23390 12484 23394 12540
rect 23330 12480 23394 12484
rect 23410 12540 23474 12544
rect 23410 12484 23414 12540
rect 23414 12484 23470 12540
rect 23470 12484 23474 12540
rect 23410 12480 23474 12484
rect 7300 11996 7364 12000
rect 7300 11940 7304 11996
rect 7304 11940 7360 11996
rect 7360 11940 7364 11996
rect 7300 11936 7364 11940
rect 7380 11996 7444 12000
rect 7380 11940 7384 11996
rect 7384 11940 7440 11996
rect 7440 11940 7444 11996
rect 7380 11936 7444 11940
rect 7460 11996 7524 12000
rect 7460 11940 7464 11996
rect 7464 11940 7520 11996
rect 7520 11940 7524 11996
rect 7460 11936 7524 11940
rect 7540 11996 7604 12000
rect 7540 11940 7544 11996
rect 7544 11940 7600 11996
rect 7600 11940 7604 11996
rect 7540 11936 7604 11940
rect 13648 11996 13712 12000
rect 13648 11940 13652 11996
rect 13652 11940 13708 11996
rect 13708 11940 13712 11996
rect 13648 11936 13712 11940
rect 13728 11996 13792 12000
rect 13728 11940 13732 11996
rect 13732 11940 13788 11996
rect 13788 11940 13792 11996
rect 13728 11936 13792 11940
rect 13808 11996 13872 12000
rect 13808 11940 13812 11996
rect 13812 11940 13868 11996
rect 13868 11940 13872 11996
rect 13808 11936 13872 11940
rect 13888 11996 13952 12000
rect 13888 11940 13892 11996
rect 13892 11940 13948 11996
rect 13948 11940 13952 11996
rect 13888 11936 13952 11940
rect 19996 11996 20060 12000
rect 19996 11940 20000 11996
rect 20000 11940 20056 11996
rect 20056 11940 20060 11996
rect 19996 11936 20060 11940
rect 20076 11996 20140 12000
rect 20076 11940 20080 11996
rect 20080 11940 20136 11996
rect 20136 11940 20140 11996
rect 20076 11936 20140 11940
rect 20156 11996 20220 12000
rect 20156 11940 20160 11996
rect 20160 11940 20216 11996
rect 20216 11940 20220 11996
rect 20156 11936 20220 11940
rect 20236 11996 20300 12000
rect 20236 11940 20240 11996
rect 20240 11940 20296 11996
rect 20296 11940 20300 11996
rect 20236 11936 20300 11940
rect 26344 11996 26408 12000
rect 26344 11940 26348 11996
rect 26348 11940 26404 11996
rect 26404 11940 26408 11996
rect 26344 11936 26408 11940
rect 26424 11996 26488 12000
rect 26424 11940 26428 11996
rect 26428 11940 26484 11996
rect 26484 11940 26488 11996
rect 26424 11936 26488 11940
rect 26504 11996 26568 12000
rect 26504 11940 26508 11996
rect 26508 11940 26564 11996
rect 26564 11940 26568 11996
rect 26504 11936 26568 11940
rect 26584 11996 26648 12000
rect 26584 11940 26588 11996
rect 26588 11940 26644 11996
rect 26644 11940 26648 11996
rect 26584 11936 26648 11940
rect 4126 11452 4190 11456
rect 4126 11396 4130 11452
rect 4130 11396 4186 11452
rect 4186 11396 4190 11452
rect 4126 11392 4190 11396
rect 4206 11452 4270 11456
rect 4206 11396 4210 11452
rect 4210 11396 4266 11452
rect 4266 11396 4270 11452
rect 4206 11392 4270 11396
rect 4286 11452 4350 11456
rect 4286 11396 4290 11452
rect 4290 11396 4346 11452
rect 4346 11396 4350 11452
rect 4286 11392 4350 11396
rect 4366 11452 4430 11456
rect 4366 11396 4370 11452
rect 4370 11396 4426 11452
rect 4426 11396 4430 11452
rect 4366 11392 4430 11396
rect 10474 11452 10538 11456
rect 10474 11396 10478 11452
rect 10478 11396 10534 11452
rect 10534 11396 10538 11452
rect 10474 11392 10538 11396
rect 10554 11452 10618 11456
rect 10554 11396 10558 11452
rect 10558 11396 10614 11452
rect 10614 11396 10618 11452
rect 10554 11392 10618 11396
rect 10634 11452 10698 11456
rect 10634 11396 10638 11452
rect 10638 11396 10694 11452
rect 10694 11396 10698 11452
rect 10634 11392 10698 11396
rect 10714 11452 10778 11456
rect 10714 11396 10718 11452
rect 10718 11396 10774 11452
rect 10774 11396 10778 11452
rect 10714 11392 10778 11396
rect 16822 11452 16886 11456
rect 16822 11396 16826 11452
rect 16826 11396 16882 11452
rect 16882 11396 16886 11452
rect 16822 11392 16886 11396
rect 16902 11452 16966 11456
rect 16902 11396 16906 11452
rect 16906 11396 16962 11452
rect 16962 11396 16966 11452
rect 16902 11392 16966 11396
rect 16982 11452 17046 11456
rect 16982 11396 16986 11452
rect 16986 11396 17042 11452
rect 17042 11396 17046 11452
rect 16982 11392 17046 11396
rect 17062 11452 17126 11456
rect 17062 11396 17066 11452
rect 17066 11396 17122 11452
rect 17122 11396 17126 11452
rect 17062 11392 17126 11396
rect 23170 11452 23234 11456
rect 23170 11396 23174 11452
rect 23174 11396 23230 11452
rect 23230 11396 23234 11452
rect 23170 11392 23234 11396
rect 23250 11452 23314 11456
rect 23250 11396 23254 11452
rect 23254 11396 23310 11452
rect 23310 11396 23314 11452
rect 23250 11392 23314 11396
rect 23330 11452 23394 11456
rect 23330 11396 23334 11452
rect 23334 11396 23390 11452
rect 23390 11396 23394 11452
rect 23330 11392 23394 11396
rect 23410 11452 23474 11456
rect 23410 11396 23414 11452
rect 23414 11396 23470 11452
rect 23470 11396 23474 11452
rect 23410 11392 23474 11396
rect 7300 10908 7364 10912
rect 7300 10852 7304 10908
rect 7304 10852 7360 10908
rect 7360 10852 7364 10908
rect 7300 10848 7364 10852
rect 7380 10908 7444 10912
rect 7380 10852 7384 10908
rect 7384 10852 7440 10908
rect 7440 10852 7444 10908
rect 7380 10848 7444 10852
rect 7460 10908 7524 10912
rect 7460 10852 7464 10908
rect 7464 10852 7520 10908
rect 7520 10852 7524 10908
rect 7460 10848 7524 10852
rect 7540 10908 7604 10912
rect 7540 10852 7544 10908
rect 7544 10852 7600 10908
rect 7600 10852 7604 10908
rect 7540 10848 7604 10852
rect 13648 10908 13712 10912
rect 13648 10852 13652 10908
rect 13652 10852 13708 10908
rect 13708 10852 13712 10908
rect 13648 10848 13712 10852
rect 13728 10908 13792 10912
rect 13728 10852 13732 10908
rect 13732 10852 13788 10908
rect 13788 10852 13792 10908
rect 13728 10848 13792 10852
rect 13808 10908 13872 10912
rect 13808 10852 13812 10908
rect 13812 10852 13868 10908
rect 13868 10852 13872 10908
rect 13808 10848 13872 10852
rect 13888 10908 13952 10912
rect 13888 10852 13892 10908
rect 13892 10852 13948 10908
rect 13948 10852 13952 10908
rect 13888 10848 13952 10852
rect 19996 10908 20060 10912
rect 19996 10852 20000 10908
rect 20000 10852 20056 10908
rect 20056 10852 20060 10908
rect 19996 10848 20060 10852
rect 20076 10908 20140 10912
rect 20076 10852 20080 10908
rect 20080 10852 20136 10908
rect 20136 10852 20140 10908
rect 20076 10848 20140 10852
rect 20156 10908 20220 10912
rect 20156 10852 20160 10908
rect 20160 10852 20216 10908
rect 20216 10852 20220 10908
rect 20156 10848 20220 10852
rect 20236 10908 20300 10912
rect 20236 10852 20240 10908
rect 20240 10852 20296 10908
rect 20296 10852 20300 10908
rect 20236 10848 20300 10852
rect 26344 10908 26408 10912
rect 26344 10852 26348 10908
rect 26348 10852 26404 10908
rect 26404 10852 26408 10908
rect 26344 10848 26408 10852
rect 26424 10908 26488 10912
rect 26424 10852 26428 10908
rect 26428 10852 26484 10908
rect 26484 10852 26488 10908
rect 26424 10848 26488 10852
rect 26504 10908 26568 10912
rect 26504 10852 26508 10908
rect 26508 10852 26564 10908
rect 26564 10852 26568 10908
rect 26504 10848 26568 10852
rect 26584 10908 26648 10912
rect 26584 10852 26588 10908
rect 26588 10852 26644 10908
rect 26644 10852 26648 10908
rect 26584 10848 26648 10852
rect 4126 10364 4190 10368
rect 4126 10308 4130 10364
rect 4130 10308 4186 10364
rect 4186 10308 4190 10364
rect 4126 10304 4190 10308
rect 4206 10364 4270 10368
rect 4206 10308 4210 10364
rect 4210 10308 4266 10364
rect 4266 10308 4270 10364
rect 4206 10304 4270 10308
rect 4286 10364 4350 10368
rect 4286 10308 4290 10364
rect 4290 10308 4346 10364
rect 4346 10308 4350 10364
rect 4286 10304 4350 10308
rect 4366 10364 4430 10368
rect 4366 10308 4370 10364
rect 4370 10308 4426 10364
rect 4426 10308 4430 10364
rect 4366 10304 4430 10308
rect 10474 10364 10538 10368
rect 10474 10308 10478 10364
rect 10478 10308 10534 10364
rect 10534 10308 10538 10364
rect 10474 10304 10538 10308
rect 10554 10364 10618 10368
rect 10554 10308 10558 10364
rect 10558 10308 10614 10364
rect 10614 10308 10618 10364
rect 10554 10304 10618 10308
rect 10634 10364 10698 10368
rect 10634 10308 10638 10364
rect 10638 10308 10694 10364
rect 10694 10308 10698 10364
rect 10634 10304 10698 10308
rect 10714 10364 10778 10368
rect 10714 10308 10718 10364
rect 10718 10308 10774 10364
rect 10774 10308 10778 10364
rect 10714 10304 10778 10308
rect 16822 10364 16886 10368
rect 16822 10308 16826 10364
rect 16826 10308 16882 10364
rect 16882 10308 16886 10364
rect 16822 10304 16886 10308
rect 16902 10364 16966 10368
rect 16902 10308 16906 10364
rect 16906 10308 16962 10364
rect 16962 10308 16966 10364
rect 16902 10304 16966 10308
rect 16982 10364 17046 10368
rect 16982 10308 16986 10364
rect 16986 10308 17042 10364
rect 17042 10308 17046 10364
rect 16982 10304 17046 10308
rect 17062 10364 17126 10368
rect 17062 10308 17066 10364
rect 17066 10308 17122 10364
rect 17122 10308 17126 10364
rect 17062 10304 17126 10308
rect 23170 10364 23234 10368
rect 23170 10308 23174 10364
rect 23174 10308 23230 10364
rect 23230 10308 23234 10364
rect 23170 10304 23234 10308
rect 23250 10364 23314 10368
rect 23250 10308 23254 10364
rect 23254 10308 23310 10364
rect 23310 10308 23314 10364
rect 23250 10304 23314 10308
rect 23330 10364 23394 10368
rect 23330 10308 23334 10364
rect 23334 10308 23390 10364
rect 23390 10308 23394 10364
rect 23330 10304 23394 10308
rect 23410 10364 23474 10368
rect 23410 10308 23414 10364
rect 23414 10308 23470 10364
rect 23470 10308 23474 10364
rect 23410 10304 23474 10308
rect 7300 9820 7364 9824
rect 7300 9764 7304 9820
rect 7304 9764 7360 9820
rect 7360 9764 7364 9820
rect 7300 9760 7364 9764
rect 7380 9820 7444 9824
rect 7380 9764 7384 9820
rect 7384 9764 7440 9820
rect 7440 9764 7444 9820
rect 7380 9760 7444 9764
rect 7460 9820 7524 9824
rect 7460 9764 7464 9820
rect 7464 9764 7520 9820
rect 7520 9764 7524 9820
rect 7460 9760 7524 9764
rect 7540 9820 7604 9824
rect 7540 9764 7544 9820
rect 7544 9764 7600 9820
rect 7600 9764 7604 9820
rect 7540 9760 7604 9764
rect 13648 9820 13712 9824
rect 13648 9764 13652 9820
rect 13652 9764 13708 9820
rect 13708 9764 13712 9820
rect 13648 9760 13712 9764
rect 13728 9820 13792 9824
rect 13728 9764 13732 9820
rect 13732 9764 13788 9820
rect 13788 9764 13792 9820
rect 13728 9760 13792 9764
rect 13808 9820 13872 9824
rect 13808 9764 13812 9820
rect 13812 9764 13868 9820
rect 13868 9764 13872 9820
rect 13808 9760 13872 9764
rect 13888 9820 13952 9824
rect 13888 9764 13892 9820
rect 13892 9764 13948 9820
rect 13948 9764 13952 9820
rect 13888 9760 13952 9764
rect 19996 9820 20060 9824
rect 19996 9764 20000 9820
rect 20000 9764 20056 9820
rect 20056 9764 20060 9820
rect 19996 9760 20060 9764
rect 20076 9820 20140 9824
rect 20076 9764 20080 9820
rect 20080 9764 20136 9820
rect 20136 9764 20140 9820
rect 20076 9760 20140 9764
rect 20156 9820 20220 9824
rect 20156 9764 20160 9820
rect 20160 9764 20216 9820
rect 20216 9764 20220 9820
rect 20156 9760 20220 9764
rect 20236 9820 20300 9824
rect 20236 9764 20240 9820
rect 20240 9764 20296 9820
rect 20296 9764 20300 9820
rect 20236 9760 20300 9764
rect 26344 9820 26408 9824
rect 26344 9764 26348 9820
rect 26348 9764 26404 9820
rect 26404 9764 26408 9820
rect 26344 9760 26408 9764
rect 26424 9820 26488 9824
rect 26424 9764 26428 9820
rect 26428 9764 26484 9820
rect 26484 9764 26488 9820
rect 26424 9760 26488 9764
rect 26504 9820 26568 9824
rect 26504 9764 26508 9820
rect 26508 9764 26564 9820
rect 26564 9764 26568 9820
rect 26504 9760 26568 9764
rect 26584 9820 26648 9824
rect 26584 9764 26588 9820
rect 26588 9764 26644 9820
rect 26644 9764 26648 9820
rect 26584 9760 26648 9764
rect 4126 9276 4190 9280
rect 4126 9220 4130 9276
rect 4130 9220 4186 9276
rect 4186 9220 4190 9276
rect 4126 9216 4190 9220
rect 4206 9276 4270 9280
rect 4206 9220 4210 9276
rect 4210 9220 4266 9276
rect 4266 9220 4270 9276
rect 4206 9216 4270 9220
rect 4286 9276 4350 9280
rect 4286 9220 4290 9276
rect 4290 9220 4346 9276
rect 4346 9220 4350 9276
rect 4286 9216 4350 9220
rect 4366 9276 4430 9280
rect 4366 9220 4370 9276
rect 4370 9220 4426 9276
rect 4426 9220 4430 9276
rect 4366 9216 4430 9220
rect 10474 9276 10538 9280
rect 10474 9220 10478 9276
rect 10478 9220 10534 9276
rect 10534 9220 10538 9276
rect 10474 9216 10538 9220
rect 10554 9276 10618 9280
rect 10554 9220 10558 9276
rect 10558 9220 10614 9276
rect 10614 9220 10618 9276
rect 10554 9216 10618 9220
rect 10634 9276 10698 9280
rect 10634 9220 10638 9276
rect 10638 9220 10694 9276
rect 10694 9220 10698 9276
rect 10634 9216 10698 9220
rect 10714 9276 10778 9280
rect 10714 9220 10718 9276
rect 10718 9220 10774 9276
rect 10774 9220 10778 9276
rect 10714 9216 10778 9220
rect 16822 9276 16886 9280
rect 16822 9220 16826 9276
rect 16826 9220 16882 9276
rect 16882 9220 16886 9276
rect 16822 9216 16886 9220
rect 16902 9276 16966 9280
rect 16902 9220 16906 9276
rect 16906 9220 16962 9276
rect 16962 9220 16966 9276
rect 16902 9216 16966 9220
rect 16982 9276 17046 9280
rect 16982 9220 16986 9276
rect 16986 9220 17042 9276
rect 17042 9220 17046 9276
rect 16982 9216 17046 9220
rect 17062 9276 17126 9280
rect 17062 9220 17066 9276
rect 17066 9220 17122 9276
rect 17122 9220 17126 9276
rect 17062 9216 17126 9220
rect 23170 9276 23234 9280
rect 23170 9220 23174 9276
rect 23174 9220 23230 9276
rect 23230 9220 23234 9276
rect 23170 9216 23234 9220
rect 23250 9276 23314 9280
rect 23250 9220 23254 9276
rect 23254 9220 23310 9276
rect 23310 9220 23314 9276
rect 23250 9216 23314 9220
rect 23330 9276 23394 9280
rect 23330 9220 23334 9276
rect 23334 9220 23390 9276
rect 23390 9220 23394 9276
rect 23330 9216 23394 9220
rect 23410 9276 23474 9280
rect 23410 9220 23414 9276
rect 23414 9220 23470 9276
rect 23470 9220 23474 9276
rect 23410 9216 23474 9220
rect 7300 8732 7364 8736
rect 7300 8676 7304 8732
rect 7304 8676 7360 8732
rect 7360 8676 7364 8732
rect 7300 8672 7364 8676
rect 7380 8732 7444 8736
rect 7380 8676 7384 8732
rect 7384 8676 7440 8732
rect 7440 8676 7444 8732
rect 7380 8672 7444 8676
rect 7460 8732 7524 8736
rect 7460 8676 7464 8732
rect 7464 8676 7520 8732
rect 7520 8676 7524 8732
rect 7460 8672 7524 8676
rect 7540 8732 7604 8736
rect 7540 8676 7544 8732
rect 7544 8676 7600 8732
rect 7600 8676 7604 8732
rect 7540 8672 7604 8676
rect 13648 8732 13712 8736
rect 13648 8676 13652 8732
rect 13652 8676 13708 8732
rect 13708 8676 13712 8732
rect 13648 8672 13712 8676
rect 13728 8732 13792 8736
rect 13728 8676 13732 8732
rect 13732 8676 13788 8732
rect 13788 8676 13792 8732
rect 13728 8672 13792 8676
rect 13808 8732 13872 8736
rect 13808 8676 13812 8732
rect 13812 8676 13868 8732
rect 13868 8676 13872 8732
rect 13808 8672 13872 8676
rect 13888 8732 13952 8736
rect 13888 8676 13892 8732
rect 13892 8676 13948 8732
rect 13948 8676 13952 8732
rect 13888 8672 13952 8676
rect 19996 8732 20060 8736
rect 19996 8676 20000 8732
rect 20000 8676 20056 8732
rect 20056 8676 20060 8732
rect 19996 8672 20060 8676
rect 20076 8732 20140 8736
rect 20076 8676 20080 8732
rect 20080 8676 20136 8732
rect 20136 8676 20140 8732
rect 20076 8672 20140 8676
rect 20156 8732 20220 8736
rect 20156 8676 20160 8732
rect 20160 8676 20216 8732
rect 20216 8676 20220 8732
rect 20156 8672 20220 8676
rect 20236 8732 20300 8736
rect 20236 8676 20240 8732
rect 20240 8676 20296 8732
rect 20296 8676 20300 8732
rect 20236 8672 20300 8676
rect 26344 8732 26408 8736
rect 26344 8676 26348 8732
rect 26348 8676 26404 8732
rect 26404 8676 26408 8732
rect 26344 8672 26408 8676
rect 26424 8732 26488 8736
rect 26424 8676 26428 8732
rect 26428 8676 26484 8732
rect 26484 8676 26488 8732
rect 26424 8672 26488 8676
rect 26504 8732 26568 8736
rect 26504 8676 26508 8732
rect 26508 8676 26564 8732
rect 26564 8676 26568 8732
rect 26504 8672 26568 8676
rect 26584 8732 26648 8736
rect 26584 8676 26588 8732
rect 26588 8676 26644 8732
rect 26644 8676 26648 8732
rect 26584 8672 26648 8676
rect 4126 8188 4190 8192
rect 4126 8132 4130 8188
rect 4130 8132 4186 8188
rect 4186 8132 4190 8188
rect 4126 8128 4190 8132
rect 4206 8188 4270 8192
rect 4206 8132 4210 8188
rect 4210 8132 4266 8188
rect 4266 8132 4270 8188
rect 4206 8128 4270 8132
rect 4286 8188 4350 8192
rect 4286 8132 4290 8188
rect 4290 8132 4346 8188
rect 4346 8132 4350 8188
rect 4286 8128 4350 8132
rect 4366 8188 4430 8192
rect 4366 8132 4370 8188
rect 4370 8132 4426 8188
rect 4426 8132 4430 8188
rect 4366 8128 4430 8132
rect 10474 8188 10538 8192
rect 10474 8132 10478 8188
rect 10478 8132 10534 8188
rect 10534 8132 10538 8188
rect 10474 8128 10538 8132
rect 10554 8188 10618 8192
rect 10554 8132 10558 8188
rect 10558 8132 10614 8188
rect 10614 8132 10618 8188
rect 10554 8128 10618 8132
rect 10634 8188 10698 8192
rect 10634 8132 10638 8188
rect 10638 8132 10694 8188
rect 10694 8132 10698 8188
rect 10634 8128 10698 8132
rect 10714 8188 10778 8192
rect 10714 8132 10718 8188
rect 10718 8132 10774 8188
rect 10774 8132 10778 8188
rect 10714 8128 10778 8132
rect 16822 8188 16886 8192
rect 16822 8132 16826 8188
rect 16826 8132 16882 8188
rect 16882 8132 16886 8188
rect 16822 8128 16886 8132
rect 16902 8188 16966 8192
rect 16902 8132 16906 8188
rect 16906 8132 16962 8188
rect 16962 8132 16966 8188
rect 16902 8128 16966 8132
rect 16982 8188 17046 8192
rect 16982 8132 16986 8188
rect 16986 8132 17042 8188
rect 17042 8132 17046 8188
rect 16982 8128 17046 8132
rect 17062 8188 17126 8192
rect 17062 8132 17066 8188
rect 17066 8132 17122 8188
rect 17122 8132 17126 8188
rect 17062 8128 17126 8132
rect 23170 8188 23234 8192
rect 23170 8132 23174 8188
rect 23174 8132 23230 8188
rect 23230 8132 23234 8188
rect 23170 8128 23234 8132
rect 23250 8188 23314 8192
rect 23250 8132 23254 8188
rect 23254 8132 23310 8188
rect 23310 8132 23314 8188
rect 23250 8128 23314 8132
rect 23330 8188 23394 8192
rect 23330 8132 23334 8188
rect 23334 8132 23390 8188
rect 23390 8132 23394 8188
rect 23330 8128 23394 8132
rect 23410 8188 23474 8192
rect 23410 8132 23414 8188
rect 23414 8132 23470 8188
rect 23470 8132 23474 8188
rect 23410 8128 23474 8132
rect 7300 7644 7364 7648
rect 7300 7588 7304 7644
rect 7304 7588 7360 7644
rect 7360 7588 7364 7644
rect 7300 7584 7364 7588
rect 7380 7644 7444 7648
rect 7380 7588 7384 7644
rect 7384 7588 7440 7644
rect 7440 7588 7444 7644
rect 7380 7584 7444 7588
rect 7460 7644 7524 7648
rect 7460 7588 7464 7644
rect 7464 7588 7520 7644
rect 7520 7588 7524 7644
rect 7460 7584 7524 7588
rect 7540 7644 7604 7648
rect 7540 7588 7544 7644
rect 7544 7588 7600 7644
rect 7600 7588 7604 7644
rect 7540 7584 7604 7588
rect 13648 7644 13712 7648
rect 13648 7588 13652 7644
rect 13652 7588 13708 7644
rect 13708 7588 13712 7644
rect 13648 7584 13712 7588
rect 13728 7644 13792 7648
rect 13728 7588 13732 7644
rect 13732 7588 13788 7644
rect 13788 7588 13792 7644
rect 13728 7584 13792 7588
rect 13808 7644 13872 7648
rect 13808 7588 13812 7644
rect 13812 7588 13868 7644
rect 13868 7588 13872 7644
rect 13808 7584 13872 7588
rect 13888 7644 13952 7648
rect 13888 7588 13892 7644
rect 13892 7588 13948 7644
rect 13948 7588 13952 7644
rect 13888 7584 13952 7588
rect 19996 7644 20060 7648
rect 19996 7588 20000 7644
rect 20000 7588 20056 7644
rect 20056 7588 20060 7644
rect 19996 7584 20060 7588
rect 20076 7644 20140 7648
rect 20076 7588 20080 7644
rect 20080 7588 20136 7644
rect 20136 7588 20140 7644
rect 20076 7584 20140 7588
rect 20156 7644 20220 7648
rect 20156 7588 20160 7644
rect 20160 7588 20216 7644
rect 20216 7588 20220 7644
rect 20156 7584 20220 7588
rect 20236 7644 20300 7648
rect 20236 7588 20240 7644
rect 20240 7588 20296 7644
rect 20296 7588 20300 7644
rect 20236 7584 20300 7588
rect 26344 7644 26408 7648
rect 26344 7588 26348 7644
rect 26348 7588 26404 7644
rect 26404 7588 26408 7644
rect 26344 7584 26408 7588
rect 26424 7644 26488 7648
rect 26424 7588 26428 7644
rect 26428 7588 26484 7644
rect 26484 7588 26488 7644
rect 26424 7584 26488 7588
rect 26504 7644 26568 7648
rect 26504 7588 26508 7644
rect 26508 7588 26564 7644
rect 26564 7588 26568 7644
rect 26504 7584 26568 7588
rect 26584 7644 26648 7648
rect 26584 7588 26588 7644
rect 26588 7588 26644 7644
rect 26644 7588 26648 7644
rect 26584 7584 26648 7588
rect 4126 7100 4190 7104
rect 4126 7044 4130 7100
rect 4130 7044 4186 7100
rect 4186 7044 4190 7100
rect 4126 7040 4190 7044
rect 4206 7100 4270 7104
rect 4206 7044 4210 7100
rect 4210 7044 4266 7100
rect 4266 7044 4270 7100
rect 4206 7040 4270 7044
rect 4286 7100 4350 7104
rect 4286 7044 4290 7100
rect 4290 7044 4346 7100
rect 4346 7044 4350 7100
rect 4286 7040 4350 7044
rect 4366 7100 4430 7104
rect 4366 7044 4370 7100
rect 4370 7044 4426 7100
rect 4426 7044 4430 7100
rect 4366 7040 4430 7044
rect 10474 7100 10538 7104
rect 10474 7044 10478 7100
rect 10478 7044 10534 7100
rect 10534 7044 10538 7100
rect 10474 7040 10538 7044
rect 10554 7100 10618 7104
rect 10554 7044 10558 7100
rect 10558 7044 10614 7100
rect 10614 7044 10618 7100
rect 10554 7040 10618 7044
rect 10634 7100 10698 7104
rect 10634 7044 10638 7100
rect 10638 7044 10694 7100
rect 10694 7044 10698 7100
rect 10634 7040 10698 7044
rect 10714 7100 10778 7104
rect 10714 7044 10718 7100
rect 10718 7044 10774 7100
rect 10774 7044 10778 7100
rect 10714 7040 10778 7044
rect 16822 7100 16886 7104
rect 16822 7044 16826 7100
rect 16826 7044 16882 7100
rect 16882 7044 16886 7100
rect 16822 7040 16886 7044
rect 16902 7100 16966 7104
rect 16902 7044 16906 7100
rect 16906 7044 16962 7100
rect 16962 7044 16966 7100
rect 16902 7040 16966 7044
rect 16982 7100 17046 7104
rect 16982 7044 16986 7100
rect 16986 7044 17042 7100
rect 17042 7044 17046 7100
rect 16982 7040 17046 7044
rect 17062 7100 17126 7104
rect 17062 7044 17066 7100
rect 17066 7044 17122 7100
rect 17122 7044 17126 7100
rect 17062 7040 17126 7044
rect 23170 7100 23234 7104
rect 23170 7044 23174 7100
rect 23174 7044 23230 7100
rect 23230 7044 23234 7100
rect 23170 7040 23234 7044
rect 23250 7100 23314 7104
rect 23250 7044 23254 7100
rect 23254 7044 23310 7100
rect 23310 7044 23314 7100
rect 23250 7040 23314 7044
rect 23330 7100 23394 7104
rect 23330 7044 23334 7100
rect 23334 7044 23390 7100
rect 23390 7044 23394 7100
rect 23330 7040 23394 7044
rect 23410 7100 23474 7104
rect 23410 7044 23414 7100
rect 23414 7044 23470 7100
rect 23470 7044 23474 7100
rect 23410 7040 23474 7044
rect 7300 6556 7364 6560
rect 7300 6500 7304 6556
rect 7304 6500 7360 6556
rect 7360 6500 7364 6556
rect 7300 6496 7364 6500
rect 7380 6556 7444 6560
rect 7380 6500 7384 6556
rect 7384 6500 7440 6556
rect 7440 6500 7444 6556
rect 7380 6496 7444 6500
rect 7460 6556 7524 6560
rect 7460 6500 7464 6556
rect 7464 6500 7520 6556
rect 7520 6500 7524 6556
rect 7460 6496 7524 6500
rect 7540 6556 7604 6560
rect 7540 6500 7544 6556
rect 7544 6500 7600 6556
rect 7600 6500 7604 6556
rect 7540 6496 7604 6500
rect 13648 6556 13712 6560
rect 13648 6500 13652 6556
rect 13652 6500 13708 6556
rect 13708 6500 13712 6556
rect 13648 6496 13712 6500
rect 13728 6556 13792 6560
rect 13728 6500 13732 6556
rect 13732 6500 13788 6556
rect 13788 6500 13792 6556
rect 13728 6496 13792 6500
rect 13808 6556 13872 6560
rect 13808 6500 13812 6556
rect 13812 6500 13868 6556
rect 13868 6500 13872 6556
rect 13808 6496 13872 6500
rect 13888 6556 13952 6560
rect 13888 6500 13892 6556
rect 13892 6500 13948 6556
rect 13948 6500 13952 6556
rect 13888 6496 13952 6500
rect 19996 6556 20060 6560
rect 19996 6500 20000 6556
rect 20000 6500 20056 6556
rect 20056 6500 20060 6556
rect 19996 6496 20060 6500
rect 20076 6556 20140 6560
rect 20076 6500 20080 6556
rect 20080 6500 20136 6556
rect 20136 6500 20140 6556
rect 20076 6496 20140 6500
rect 20156 6556 20220 6560
rect 20156 6500 20160 6556
rect 20160 6500 20216 6556
rect 20216 6500 20220 6556
rect 20156 6496 20220 6500
rect 20236 6556 20300 6560
rect 20236 6500 20240 6556
rect 20240 6500 20296 6556
rect 20296 6500 20300 6556
rect 20236 6496 20300 6500
rect 26344 6556 26408 6560
rect 26344 6500 26348 6556
rect 26348 6500 26404 6556
rect 26404 6500 26408 6556
rect 26344 6496 26408 6500
rect 26424 6556 26488 6560
rect 26424 6500 26428 6556
rect 26428 6500 26484 6556
rect 26484 6500 26488 6556
rect 26424 6496 26488 6500
rect 26504 6556 26568 6560
rect 26504 6500 26508 6556
rect 26508 6500 26564 6556
rect 26564 6500 26568 6556
rect 26504 6496 26568 6500
rect 26584 6556 26648 6560
rect 26584 6500 26588 6556
rect 26588 6500 26644 6556
rect 26644 6500 26648 6556
rect 26584 6496 26648 6500
rect 4126 6012 4190 6016
rect 4126 5956 4130 6012
rect 4130 5956 4186 6012
rect 4186 5956 4190 6012
rect 4126 5952 4190 5956
rect 4206 6012 4270 6016
rect 4206 5956 4210 6012
rect 4210 5956 4266 6012
rect 4266 5956 4270 6012
rect 4206 5952 4270 5956
rect 4286 6012 4350 6016
rect 4286 5956 4290 6012
rect 4290 5956 4346 6012
rect 4346 5956 4350 6012
rect 4286 5952 4350 5956
rect 4366 6012 4430 6016
rect 4366 5956 4370 6012
rect 4370 5956 4426 6012
rect 4426 5956 4430 6012
rect 4366 5952 4430 5956
rect 10474 6012 10538 6016
rect 10474 5956 10478 6012
rect 10478 5956 10534 6012
rect 10534 5956 10538 6012
rect 10474 5952 10538 5956
rect 10554 6012 10618 6016
rect 10554 5956 10558 6012
rect 10558 5956 10614 6012
rect 10614 5956 10618 6012
rect 10554 5952 10618 5956
rect 10634 6012 10698 6016
rect 10634 5956 10638 6012
rect 10638 5956 10694 6012
rect 10694 5956 10698 6012
rect 10634 5952 10698 5956
rect 10714 6012 10778 6016
rect 10714 5956 10718 6012
rect 10718 5956 10774 6012
rect 10774 5956 10778 6012
rect 10714 5952 10778 5956
rect 16822 6012 16886 6016
rect 16822 5956 16826 6012
rect 16826 5956 16882 6012
rect 16882 5956 16886 6012
rect 16822 5952 16886 5956
rect 16902 6012 16966 6016
rect 16902 5956 16906 6012
rect 16906 5956 16962 6012
rect 16962 5956 16966 6012
rect 16902 5952 16966 5956
rect 16982 6012 17046 6016
rect 16982 5956 16986 6012
rect 16986 5956 17042 6012
rect 17042 5956 17046 6012
rect 16982 5952 17046 5956
rect 17062 6012 17126 6016
rect 17062 5956 17066 6012
rect 17066 5956 17122 6012
rect 17122 5956 17126 6012
rect 17062 5952 17126 5956
rect 23170 6012 23234 6016
rect 23170 5956 23174 6012
rect 23174 5956 23230 6012
rect 23230 5956 23234 6012
rect 23170 5952 23234 5956
rect 23250 6012 23314 6016
rect 23250 5956 23254 6012
rect 23254 5956 23310 6012
rect 23310 5956 23314 6012
rect 23250 5952 23314 5956
rect 23330 6012 23394 6016
rect 23330 5956 23334 6012
rect 23334 5956 23390 6012
rect 23390 5956 23394 6012
rect 23330 5952 23394 5956
rect 23410 6012 23474 6016
rect 23410 5956 23414 6012
rect 23414 5956 23470 6012
rect 23470 5956 23474 6012
rect 23410 5952 23474 5956
rect 7300 5468 7364 5472
rect 7300 5412 7304 5468
rect 7304 5412 7360 5468
rect 7360 5412 7364 5468
rect 7300 5408 7364 5412
rect 7380 5468 7444 5472
rect 7380 5412 7384 5468
rect 7384 5412 7440 5468
rect 7440 5412 7444 5468
rect 7380 5408 7444 5412
rect 7460 5468 7524 5472
rect 7460 5412 7464 5468
rect 7464 5412 7520 5468
rect 7520 5412 7524 5468
rect 7460 5408 7524 5412
rect 7540 5468 7604 5472
rect 7540 5412 7544 5468
rect 7544 5412 7600 5468
rect 7600 5412 7604 5468
rect 7540 5408 7604 5412
rect 13648 5468 13712 5472
rect 13648 5412 13652 5468
rect 13652 5412 13708 5468
rect 13708 5412 13712 5468
rect 13648 5408 13712 5412
rect 13728 5468 13792 5472
rect 13728 5412 13732 5468
rect 13732 5412 13788 5468
rect 13788 5412 13792 5468
rect 13728 5408 13792 5412
rect 13808 5468 13872 5472
rect 13808 5412 13812 5468
rect 13812 5412 13868 5468
rect 13868 5412 13872 5468
rect 13808 5408 13872 5412
rect 13888 5468 13952 5472
rect 13888 5412 13892 5468
rect 13892 5412 13948 5468
rect 13948 5412 13952 5468
rect 13888 5408 13952 5412
rect 19996 5468 20060 5472
rect 19996 5412 20000 5468
rect 20000 5412 20056 5468
rect 20056 5412 20060 5468
rect 19996 5408 20060 5412
rect 20076 5468 20140 5472
rect 20076 5412 20080 5468
rect 20080 5412 20136 5468
rect 20136 5412 20140 5468
rect 20076 5408 20140 5412
rect 20156 5468 20220 5472
rect 20156 5412 20160 5468
rect 20160 5412 20216 5468
rect 20216 5412 20220 5468
rect 20156 5408 20220 5412
rect 20236 5468 20300 5472
rect 20236 5412 20240 5468
rect 20240 5412 20296 5468
rect 20296 5412 20300 5468
rect 20236 5408 20300 5412
rect 26344 5468 26408 5472
rect 26344 5412 26348 5468
rect 26348 5412 26404 5468
rect 26404 5412 26408 5468
rect 26344 5408 26408 5412
rect 26424 5468 26488 5472
rect 26424 5412 26428 5468
rect 26428 5412 26484 5468
rect 26484 5412 26488 5468
rect 26424 5408 26488 5412
rect 26504 5468 26568 5472
rect 26504 5412 26508 5468
rect 26508 5412 26564 5468
rect 26564 5412 26568 5468
rect 26504 5408 26568 5412
rect 26584 5468 26648 5472
rect 26584 5412 26588 5468
rect 26588 5412 26644 5468
rect 26644 5412 26648 5468
rect 26584 5408 26648 5412
rect 4126 4924 4190 4928
rect 4126 4868 4130 4924
rect 4130 4868 4186 4924
rect 4186 4868 4190 4924
rect 4126 4864 4190 4868
rect 4206 4924 4270 4928
rect 4206 4868 4210 4924
rect 4210 4868 4266 4924
rect 4266 4868 4270 4924
rect 4206 4864 4270 4868
rect 4286 4924 4350 4928
rect 4286 4868 4290 4924
rect 4290 4868 4346 4924
rect 4346 4868 4350 4924
rect 4286 4864 4350 4868
rect 4366 4924 4430 4928
rect 4366 4868 4370 4924
rect 4370 4868 4426 4924
rect 4426 4868 4430 4924
rect 4366 4864 4430 4868
rect 10474 4924 10538 4928
rect 10474 4868 10478 4924
rect 10478 4868 10534 4924
rect 10534 4868 10538 4924
rect 10474 4864 10538 4868
rect 10554 4924 10618 4928
rect 10554 4868 10558 4924
rect 10558 4868 10614 4924
rect 10614 4868 10618 4924
rect 10554 4864 10618 4868
rect 10634 4924 10698 4928
rect 10634 4868 10638 4924
rect 10638 4868 10694 4924
rect 10694 4868 10698 4924
rect 10634 4864 10698 4868
rect 10714 4924 10778 4928
rect 10714 4868 10718 4924
rect 10718 4868 10774 4924
rect 10774 4868 10778 4924
rect 10714 4864 10778 4868
rect 16822 4924 16886 4928
rect 16822 4868 16826 4924
rect 16826 4868 16882 4924
rect 16882 4868 16886 4924
rect 16822 4864 16886 4868
rect 16902 4924 16966 4928
rect 16902 4868 16906 4924
rect 16906 4868 16962 4924
rect 16962 4868 16966 4924
rect 16902 4864 16966 4868
rect 16982 4924 17046 4928
rect 16982 4868 16986 4924
rect 16986 4868 17042 4924
rect 17042 4868 17046 4924
rect 16982 4864 17046 4868
rect 17062 4924 17126 4928
rect 17062 4868 17066 4924
rect 17066 4868 17122 4924
rect 17122 4868 17126 4924
rect 17062 4864 17126 4868
rect 23170 4924 23234 4928
rect 23170 4868 23174 4924
rect 23174 4868 23230 4924
rect 23230 4868 23234 4924
rect 23170 4864 23234 4868
rect 23250 4924 23314 4928
rect 23250 4868 23254 4924
rect 23254 4868 23310 4924
rect 23310 4868 23314 4924
rect 23250 4864 23314 4868
rect 23330 4924 23394 4928
rect 23330 4868 23334 4924
rect 23334 4868 23390 4924
rect 23390 4868 23394 4924
rect 23330 4864 23394 4868
rect 23410 4924 23474 4928
rect 23410 4868 23414 4924
rect 23414 4868 23470 4924
rect 23470 4868 23474 4924
rect 23410 4864 23474 4868
rect 7300 4380 7364 4384
rect 7300 4324 7304 4380
rect 7304 4324 7360 4380
rect 7360 4324 7364 4380
rect 7300 4320 7364 4324
rect 7380 4380 7444 4384
rect 7380 4324 7384 4380
rect 7384 4324 7440 4380
rect 7440 4324 7444 4380
rect 7380 4320 7444 4324
rect 7460 4380 7524 4384
rect 7460 4324 7464 4380
rect 7464 4324 7520 4380
rect 7520 4324 7524 4380
rect 7460 4320 7524 4324
rect 7540 4380 7604 4384
rect 7540 4324 7544 4380
rect 7544 4324 7600 4380
rect 7600 4324 7604 4380
rect 7540 4320 7604 4324
rect 13648 4380 13712 4384
rect 13648 4324 13652 4380
rect 13652 4324 13708 4380
rect 13708 4324 13712 4380
rect 13648 4320 13712 4324
rect 13728 4380 13792 4384
rect 13728 4324 13732 4380
rect 13732 4324 13788 4380
rect 13788 4324 13792 4380
rect 13728 4320 13792 4324
rect 13808 4380 13872 4384
rect 13808 4324 13812 4380
rect 13812 4324 13868 4380
rect 13868 4324 13872 4380
rect 13808 4320 13872 4324
rect 13888 4380 13952 4384
rect 13888 4324 13892 4380
rect 13892 4324 13948 4380
rect 13948 4324 13952 4380
rect 13888 4320 13952 4324
rect 19996 4380 20060 4384
rect 19996 4324 20000 4380
rect 20000 4324 20056 4380
rect 20056 4324 20060 4380
rect 19996 4320 20060 4324
rect 20076 4380 20140 4384
rect 20076 4324 20080 4380
rect 20080 4324 20136 4380
rect 20136 4324 20140 4380
rect 20076 4320 20140 4324
rect 20156 4380 20220 4384
rect 20156 4324 20160 4380
rect 20160 4324 20216 4380
rect 20216 4324 20220 4380
rect 20156 4320 20220 4324
rect 20236 4380 20300 4384
rect 20236 4324 20240 4380
rect 20240 4324 20296 4380
rect 20296 4324 20300 4380
rect 20236 4320 20300 4324
rect 26344 4380 26408 4384
rect 26344 4324 26348 4380
rect 26348 4324 26404 4380
rect 26404 4324 26408 4380
rect 26344 4320 26408 4324
rect 26424 4380 26488 4384
rect 26424 4324 26428 4380
rect 26428 4324 26484 4380
rect 26484 4324 26488 4380
rect 26424 4320 26488 4324
rect 26504 4380 26568 4384
rect 26504 4324 26508 4380
rect 26508 4324 26564 4380
rect 26564 4324 26568 4380
rect 26504 4320 26568 4324
rect 26584 4380 26648 4384
rect 26584 4324 26588 4380
rect 26588 4324 26644 4380
rect 26644 4324 26648 4380
rect 26584 4320 26648 4324
rect 4126 3836 4190 3840
rect 4126 3780 4130 3836
rect 4130 3780 4186 3836
rect 4186 3780 4190 3836
rect 4126 3776 4190 3780
rect 4206 3836 4270 3840
rect 4206 3780 4210 3836
rect 4210 3780 4266 3836
rect 4266 3780 4270 3836
rect 4206 3776 4270 3780
rect 4286 3836 4350 3840
rect 4286 3780 4290 3836
rect 4290 3780 4346 3836
rect 4346 3780 4350 3836
rect 4286 3776 4350 3780
rect 4366 3836 4430 3840
rect 4366 3780 4370 3836
rect 4370 3780 4426 3836
rect 4426 3780 4430 3836
rect 4366 3776 4430 3780
rect 10474 3836 10538 3840
rect 10474 3780 10478 3836
rect 10478 3780 10534 3836
rect 10534 3780 10538 3836
rect 10474 3776 10538 3780
rect 10554 3836 10618 3840
rect 10554 3780 10558 3836
rect 10558 3780 10614 3836
rect 10614 3780 10618 3836
rect 10554 3776 10618 3780
rect 10634 3836 10698 3840
rect 10634 3780 10638 3836
rect 10638 3780 10694 3836
rect 10694 3780 10698 3836
rect 10634 3776 10698 3780
rect 10714 3836 10778 3840
rect 10714 3780 10718 3836
rect 10718 3780 10774 3836
rect 10774 3780 10778 3836
rect 10714 3776 10778 3780
rect 16822 3836 16886 3840
rect 16822 3780 16826 3836
rect 16826 3780 16882 3836
rect 16882 3780 16886 3836
rect 16822 3776 16886 3780
rect 16902 3836 16966 3840
rect 16902 3780 16906 3836
rect 16906 3780 16962 3836
rect 16962 3780 16966 3836
rect 16902 3776 16966 3780
rect 16982 3836 17046 3840
rect 16982 3780 16986 3836
rect 16986 3780 17042 3836
rect 17042 3780 17046 3836
rect 16982 3776 17046 3780
rect 17062 3836 17126 3840
rect 17062 3780 17066 3836
rect 17066 3780 17122 3836
rect 17122 3780 17126 3836
rect 17062 3776 17126 3780
rect 23170 3836 23234 3840
rect 23170 3780 23174 3836
rect 23174 3780 23230 3836
rect 23230 3780 23234 3836
rect 23170 3776 23234 3780
rect 23250 3836 23314 3840
rect 23250 3780 23254 3836
rect 23254 3780 23310 3836
rect 23310 3780 23314 3836
rect 23250 3776 23314 3780
rect 23330 3836 23394 3840
rect 23330 3780 23334 3836
rect 23334 3780 23390 3836
rect 23390 3780 23394 3836
rect 23330 3776 23394 3780
rect 23410 3836 23474 3840
rect 23410 3780 23414 3836
rect 23414 3780 23470 3836
rect 23470 3780 23474 3836
rect 23410 3776 23474 3780
rect 7300 3292 7364 3296
rect 7300 3236 7304 3292
rect 7304 3236 7360 3292
rect 7360 3236 7364 3292
rect 7300 3232 7364 3236
rect 7380 3292 7444 3296
rect 7380 3236 7384 3292
rect 7384 3236 7440 3292
rect 7440 3236 7444 3292
rect 7380 3232 7444 3236
rect 7460 3292 7524 3296
rect 7460 3236 7464 3292
rect 7464 3236 7520 3292
rect 7520 3236 7524 3292
rect 7460 3232 7524 3236
rect 7540 3292 7604 3296
rect 7540 3236 7544 3292
rect 7544 3236 7600 3292
rect 7600 3236 7604 3292
rect 7540 3232 7604 3236
rect 13648 3292 13712 3296
rect 13648 3236 13652 3292
rect 13652 3236 13708 3292
rect 13708 3236 13712 3292
rect 13648 3232 13712 3236
rect 13728 3292 13792 3296
rect 13728 3236 13732 3292
rect 13732 3236 13788 3292
rect 13788 3236 13792 3292
rect 13728 3232 13792 3236
rect 13808 3292 13872 3296
rect 13808 3236 13812 3292
rect 13812 3236 13868 3292
rect 13868 3236 13872 3292
rect 13808 3232 13872 3236
rect 13888 3292 13952 3296
rect 13888 3236 13892 3292
rect 13892 3236 13948 3292
rect 13948 3236 13952 3292
rect 13888 3232 13952 3236
rect 19996 3292 20060 3296
rect 19996 3236 20000 3292
rect 20000 3236 20056 3292
rect 20056 3236 20060 3292
rect 19996 3232 20060 3236
rect 20076 3292 20140 3296
rect 20076 3236 20080 3292
rect 20080 3236 20136 3292
rect 20136 3236 20140 3292
rect 20076 3232 20140 3236
rect 20156 3292 20220 3296
rect 20156 3236 20160 3292
rect 20160 3236 20216 3292
rect 20216 3236 20220 3292
rect 20156 3232 20220 3236
rect 20236 3292 20300 3296
rect 20236 3236 20240 3292
rect 20240 3236 20296 3292
rect 20296 3236 20300 3292
rect 20236 3232 20300 3236
rect 26344 3292 26408 3296
rect 26344 3236 26348 3292
rect 26348 3236 26404 3292
rect 26404 3236 26408 3292
rect 26344 3232 26408 3236
rect 26424 3292 26488 3296
rect 26424 3236 26428 3292
rect 26428 3236 26484 3292
rect 26484 3236 26488 3292
rect 26424 3232 26488 3236
rect 26504 3292 26568 3296
rect 26504 3236 26508 3292
rect 26508 3236 26564 3292
rect 26564 3236 26568 3292
rect 26504 3232 26568 3236
rect 26584 3292 26648 3296
rect 26584 3236 26588 3292
rect 26588 3236 26644 3292
rect 26644 3236 26648 3292
rect 26584 3232 26648 3236
rect 4126 2748 4190 2752
rect 4126 2692 4130 2748
rect 4130 2692 4186 2748
rect 4186 2692 4190 2748
rect 4126 2688 4190 2692
rect 4206 2748 4270 2752
rect 4206 2692 4210 2748
rect 4210 2692 4266 2748
rect 4266 2692 4270 2748
rect 4206 2688 4270 2692
rect 4286 2748 4350 2752
rect 4286 2692 4290 2748
rect 4290 2692 4346 2748
rect 4346 2692 4350 2748
rect 4286 2688 4350 2692
rect 4366 2748 4430 2752
rect 4366 2692 4370 2748
rect 4370 2692 4426 2748
rect 4426 2692 4430 2748
rect 4366 2688 4430 2692
rect 10474 2748 10538 2752
rect 10474 2692 10478 2748
rect 10478 2692 10534 2748
rect 10534 2692 10538 2748
rect 10474 2688 10538 2692
rect 10554 2748 10618 2752
rect 10554 2692 10558 2748
rect 10558 2692 10614 2748
rect 10614 2692 10618 2748
rect 10554 2688 10618 2692
rect 10634 2748 10698 2752
rect 10634 2692 10638 2748
rect 10638 2692 10694 2748
rect 10694 2692 10698 2748
rect 10634 2688 10698 2692
rect 10714 2748 10778 2752
rect 10714 2692 10718 2748
rect 10718 2692 10774 2748
rect 10774 2692 10778 2748
rect 10714 2688 10778 2692
rect 16822 2748 16886 2752
rect 16822 2692 16826 2748
rect 16826 2692 16882 2748
rect 16882 2692 16886 2748
rect 16822 2688 16886 2692
rect 16902 2748 16966 2752
rect 16902 2692 16906 2748
rect 16906 2692 16962 2748
rect 16962 2692 16966 2748
rect 16902 2688 16966 2692
rect 16982 2748 17046 2752
rect 16982 2692 16986 2748
rect 16986 2692 17042 2748
rect 17042 2692 17046 2748
rect 16982 2688 17046 2692
rect 17062 2748 17126 2752
rect 17062 2692 17066 2748
rect 17066 2692 17122 2748
rect 17122 2692 17126 2748
rect 17062 2688 17126 2692
rect 23170 2748 23234 2752
rect 23170 2692 23174 2748
rect 23174 2692 23230 2748
rect 23230 2692 23234 2748
rect 23170 2688 23234 2692
rect 23250 2748 23314 2752
rect 23250 2692 23254 2748
rect 23254 2692 23310 2748
rect 23310 2692 23314 2748
rect 23250 2688 23314 2692
rect 23330 2748 23394 2752
rect 23330 2692 23334 2748
rect 23334 2692 23390 2748
rect 23390 2692 23394 2748
rect 23330 2688 23394 2692
rect 23410 2748 23474 2752
rect 23410 2692 23414 2748
rect 23414 2692 23470 2748
rect 23470 2692 23474 2748
rect 23410 2688 23474 2692
rect 7300 2204 7364 2208
rect 7300 2148 7304 2204
rect 7304 2148 7360 2204
rect 7360 2148 7364 2204
rect 7300 2144 7364 2148
rect 7380 2204 7444 2208
rect 7380 2148 7384 2204
rect 7384 2148 7440 2204
rect 7440 2148 7444 2204
rect 7380 2144 7444 2148
rect 7460 2204 7524 2208
rect 7460 2148 7464 2204
rect 7464 2148 7520 2204
rect 7520 2148 7524 2204
rect 7460 2144 7524 2148
rect 7540 2204 7604 2208
rect 7540 2148 7544 2204
rect 7544 2148 7600 2204
rect 7600 2148 7604 2204
rect 7540 2144 7604 2148
rect 13648 2204 13712 2208
rect 13648 2148 13652 2204
rect 13652 2148 13708 2204
rect 13708 2148 13712 2204
rect 13648 2144 13712 2148
rect 13728 2204 13792 2208
rect 13728 2148 13732 2204
rect 13732 2148 13788 2204
rect 13788 2148 13792 2204
rect 13728 2144 13792 2148
rect 13808 2204 13872 2208
rect 13808 2148 13812 2204
rect 13812 2148 13868 2204
rect 13868 2148 13872 2204
rect 13808 2144 13872 2148
rect 13888 2204 13952 2208
rect 13888 2148 13892 2204
rect 13892 2148 13948 2204
rect 13948 2148 13952 2204
rect 13888 2144 13952 2148
rect 19996 2204 20060 2208
rect 19996 2148 20000 2204
rect 20000 2148 20056 2204
rect 20056 2148 20060 2204
rect 19996 2144 20060 2148
rect 20076 2204 20140 2208
rect 20076 2148 20080 2204
rect 20080 2148 20136 2204
rect 20136 2148 20140 2204
rect 20076 2144 20140 2148
rect 20156 2204 20220 2208
rect 20156 2148 20160 2204
rect 20160 2148 20216 2204
rect 20216 2148 20220 2204
rect 20156 2144 20220 2148
rect 20236 2204 20300 2208
rect 20236 2148 20240 2204
rect 20240 2148 20296 2204
rect 20296 2148 20300 2204
rect 20236 2144 20300 2148
rect 26344 2204 26408 2208
rect 26344 2148 26348 2204
rect 26348 2148 26404 2204
rect 26404 2148 26408 2204
rect 26344 2144 26408 2148
rect 26424 2204 26488 2208
rect 26424 2148 26428 2204
rect 26428 2148 26484 2204
rect 26484 2148 26488 2204
rect 26424 2144 26488 2148
rect 26504 2204 26568 2208
rect 26504 2148 26508 2204
rect 26508 2148 26564 2204
rect 26564 2148 26568 2204
rect 26504 2144 26568 2148
rect 26584 2204 26648 2208
rect 26584 2148 26588 2204
rect 26588 2148 26644 2204
rect 26644 2148 26648 2204
rect 26584 2144 26648 2148
<< metal4 >>
rect 4118 26688 4438 27248
rect 4118 26624 4126 26688
rect 4190 26624 4206 26688
rect 4270 26624 4286 26688
rect 4350 26624 4366 26688
rect 4430 26624 4438 26688
rect 4118 25600 4438 26624
rect 4118 25536 4126 25600
rect 4190 25536 4206 25600
rect 4270 25536 4286 25600
rect 4350 25536 4366 25600
rect 4430 25536 4438 25600
rect 4118 24512 4438 25536
rect 4118 24448 4126 24512
rect 4190 24448 4206 24512
rect 4270 24448 4286 24512
rect 4350 24448 4366 24512
rect 4430 24448 4438 24512
rect 4118 23424 4438 24448
rect 4118 23360 4126 23424
rect 4190 23360 4206 23424
rect 4270 23360 4286 23424
rect 4350 23360 4366 23424
rect 4430 23360 4438 23424
rect 4118 22336 4438 23360
rect 4118 22272 4126 22336
rect 4190 22272 4206 22336
rect 4270 22272 4286 22336
rect 4350 22272 4366 22336
rect 4430 22272 4438 22336
rect 4118 21248 4438 22272
rect 4118 21184 4126 21248
rect 4190 21184 4206 21248
rect 4270 21184 4286 21248
rect 4350 21184 4366 21248
rect 4430 21184 4438 21248
rect 4118 20160 4438 21184
rect 4118 20096 4126 20160
rect 4190 20096 4206 20160
rect 4270 20096 4286 20160
rect 4350 20096 4366 20160
rect 4430 20096 4438 20160
rect 4118 19072 4438 20096
rect 4118 19008 4126 19072
rect 4190 19008 4206 19072
rect 4270 19008 4286 19072
rect 4350 19008 4366 19072
rect 4430 19008 4438 19072
rect 4118 17984 4438 19008
rect 4118 17920 4126 17984
rect 4190 17920 4206 17984
rect 4270 17920 4286 17984
rect 4350 17920 4366 17984
rect 4430 17920 4438 17984
rect 4118 16896 4438 17920
rect 4118 16832 4126 16896
rect 4190 16832 4206 16896
rect 4270 16832 4286 16896
rect 4350 16832 4366 16896
rect 4430 16832 4438 16896
rect 4118 15808 4438 16832
rect 4118 15744 4126 15808
rect 4190 15744 4206 15808
rect 4270 15744 4286 15808
rect 4350 15744 4366 15808
rect 4430 15744 4438 15808
rect 4118 14720 4438 15744
rect 4118 14656 4126 14720
rect 4190 14656 4206 14720
rect 4270 14656 4286 14720
rect 4350 14656 4366 14720
rect 4430 14656 4438 14720
rect 4118 13632 4438 14656
rect 4118 13568 4126 13632
rect 4190 13568 4206 13632
rect 4270 13568 4286 13632
rect 4350 13568 4366 13632
rect 4430 13568 4438 13632
rect 4118 12544 4438 13568
rect 4118 12480 4126 12544
rect 4190 12480 4206 12544
rect 4270 12480 4286 12544
rect 4350 12480 4366 12544
rect 4430 12480 4438 12544
rect 4118 11456 4438 12480
rect 4118 11392 4126 11456
rect 4190 11392 4206 11456
rect 4270 11392 4286 11456
rect 4350 11392 4366 11456
rect 4430 11392 4438 11456
rect 4118 10368 4438 11392
rect 4118 10304 4126 10368
rect 4190 10304 4206 10368
rect 4270 10304 4286 10368
rect 4350 10304 4366 10368
rect 4430 10304 4438 10368
rect 4118 9280 4438 10304
rect 4118 9216 4126 9280
rect 4190 9216 4206 9280
rect 4270 9216 4286 9280
rect 4350 9216 4366 9280
rect 4430 9216 4438 9280
rect 4118 8192 4438 9216
rect 4118 8128 4126 8192
rect 4190 8128 4206 8192
rect 4270 8128 4286 8192
rect 4350 8128 4366 8192
rect 4430 8128 4438 8192
rect 4118 7104 4438 8128
rect 4118 7040 4126 7104
rect 4190 7040 4206 7104
rect 4270 7040 4286 7104
rect 4350 7040 4366 7104
rect 4430 7040 4438 7104
rect 4118 6016 4438 7040
rect 4118 5952 4126 6016
rect 4190 5952 4206 6016
rect 4270 5952 4286 6016
rect 4350 5952 4366 6016
rect 4430 5952 4438 6016
rect 4118 4928 4438 5952
rect 4118 4864 4126 4928
rect 4190 4864 4206 4928
rect 4270 4864 4286 4928
rect 4350 4864 4366 4928
rect 4430 4864 4438 4928
rect 4118 3840 4438 4864
rect 4118 3776 4126 3840
rect 4190 3776 4206 3840
rect 4270 3776 4286 3840
rect 4350 3776 4366 3840
rect 4430 3776 4438 3840
rect 4118 2752 4438 3776
rect 4118 2688 4126 2752
rect 4190 2688 4206 2752
rect 4270 2688 4286 2752
rect 4350 2688 4366 2752
rect 4430 2688 4438 2752
rect 4118 2128 4438 2688
rect 7292 27232 7612 27248
rect 7292 27168 7300 27232
rect 7364 27168 7380 27232
rect 7444 27168 7460 27232
rect 7524 27168 7540 27232
rect 7604 27168 7612 27232
rect 7292 26144 7612 27168
rect 7292 26080 7300 26144
rect 7364 26080 7380 26144
rect 7444 26080 7460 26144
rect 7524 26080 7540 26144
rect 7604 26080 7612 26144
rect 7292 25056 7612 26080
rect 7292 24992 7300 25056
rect 7364 24992 7380 25056
rect 7444 24992 7460 25056
rect 7524 24992 7540 25056
rect 7604 24992 7612 25056
rect 7292 23968 7612 24992
rect 7292 23904 7300 23968
rect 7364 23904 7380 23968
rect 7444 23904 7460 23968
rect 7524 23904 7540 23968
rect 7604 23904 7612 23968
rect 7292 22880 7612 23904
rect 7292 22816 7300 22880
rect 7364 22816 7380 22880
rect 7444 22816 7460 22880
rect 7524 22816 7540 22880
rect 7604 22816 7612 22880
rect 7292 21792 7612 22816
rect 7292 21728 7300 21792
rect 7364 21728 7380 21792
rect 7444 21728 7460 21792
rect 7524 21728 7540 21792
rect 7604 21728 7612 21792
rect 7292 20704 7612 21728
rect 7292 20640 7300 20704
rect 7364 20640 7380 20704
rect 7444 20640 7460 20704
rect 7524 20640 7540 20704
rect 7604 20640 7612 20704
rect 7292 19616 7612 20640
rect 7292 19552 7300 19616
rect 7364 19552 7380 19616
rect 7444 19552 7460 19616
rect 7524 19552 7540 19616
rect 7604 19552 7612 19616
rect 7292 18528 7612 19552
rect 7292 18464 7300 18528
rect 7364 18464 7380 18528
rect 7444 18464 7460 18528
rect 7524 18464 7540 18528
rect 7604 18464 7612 18528
rect 7292 17440 7612 18464
rect 7292 17376 7300 17440
rect 7364 17376 7380 17440
rect 7444 17376 7460 17440
rect 7524 17376 7540 17440
rect 7604 17376 7612 17440
rect 7292 16352 7612 17376
rect 7292 16288 7300 16352
rect 7364 16288 7380 16352
rect 7444 16288 7460 16352
rect 7524 16288 7540 16352
rect 7604 16288 7612 16352
rect 7292 15264 7612 16288
rect 7292 15200 7300 15264
rect 7364 15200 7380 15264
rect 7444 15200 7460 15264
rect 7524 15200 7540 15264
rect 7604 15200 7612 15264
rect 7292 14176 7612 15200
rect 7292 14112 7300 14176
rect 7364 14112 7380 14176
rect 7444 14112 7460 14176
rect 7524 14112 7540 14176
rect 7604 14112 7612 14176
rect 7292 13088 7612 14112
rect 7292 13024 7300 13088
rect 7364 13024 7380 13088
rect 7444 13024 7460 13088
rect 7524 13024 7540 13088
rect 7604 13024 7612 13088
rect 7292 12000 7612 13024
rect 7292 11936 7300 12000
rect 7364 11936 7380 12000
rect 7444 11936 7460 12000
rect 7524 11936 7540 12000
rect 7604 11936 7612 12000
rect 7292 10912 7612 11936
rect 7292 10848 7300 10912
rect 7364 10848 7380 10912
rect 7444 10848 7460 10912
rect 7524 10848 7540 10912
rect 7604 10848 7612 10912
rect 7292 9824 7612 10848
rect 7292 9760 7300 9824
rect 7364 9760 7380 9824
rect 7444 9760 7460 9824
rect 7524 9760 7540 9824
rect 7604 9760 7612 9824
rect 7292 8736 7612 9760
rect 7292 8672 7300 8736
rect 7364 8672 7380 8736
rect 7444 8672 7460 8736
rect 7524 8672 7540 8736
rect 7604 8672 7612 8736
rect 7292 7648 7612 8672
rect 7292 7584 7300 7648
rect 7364 7584 7380 7648
rect 7444 7584 7460 7648
rect 7524 7584 7540 7648
rect 7604 7584 7612 7648
rect 7292 6560 7612 7584
rect 7292 6496 7300 6560
rect 7364 6496 7380 6560
rect 7444 6496 7460 6560
rect 7524 6496 7540 6560
rect 7604 6496 7612 6560
rect 7292 5472 7612 6496
rect 7292 5408 7300 5472
rect 7364 5408 7380 5472
rect 7444 5408 7460 5472
rect 7524 5408 7540 5472
rect 7604 5408 7612 5472
rect 7292 4384 7612 5408
rect 7292 4320 7300 4384
rect 7364 4320 7380 4384
rect 7444 4320 7460 4384
rect 7524 4320 7540 4384
rect 7604 4320 7612 4384
rect 7292 3296 7612 4320
rect 7292 3232 7300 3296
rect 7364 3232 7380 3296
rect 7444 3232 7460 3296
rect 7524 3232 7540 3296
rect 7604 3232 7612 3296
rect 7292 2208 7612 3232
rect 7292 2144 7300 2208
rect 7364 2144 7380 2208
rect 7444 2144 7460 2208
rect 7524 2144 7540 2208
rect 7604 2144 7612 2208
rect 7292 2128 7612 2144
rect 10466 26688 10786 27248
rect 10466 26624 10474 26688
rect 10538 26624 10554 26688
rect 10618 26624 10634 26688
rect 10698 26624 10714 26688
rect 10778 26624 10786 26688
rect 10466 25600 10786 26624
rect 10466 25536 10474 25600
rect 10538 25536 10554 25600
rect 10618 25536 10634 25600
rect 10698 25536 10714 25600
rect 10778 25536 10786 25600
rect 10466 24512 10786 25536
rect 10466 24448 10474 24512
rect 10538 24448 10554 24512
rect 10618 24448 10634 24512
rect 10698 24448 10714 24512
rect 10778 24448 10786 24512
rect 10466 23424 10786 24448
rect 10466 23360 10474 23424
rect 10538 23360 10554 23424
rect 10618 23360 10634 23424
rect 10698 23360 10714 23424
rect 10778 23360 10786 23424
rect 10466 22336 10786 23360
rect 10466 22272 10474 22336
rect 10538 22272 10554 22336
rect 10618 22272 10634 22336
rect 10698 22272 10714 22336
rect 10778 22272 10786 22336
rect 10466 21248 10786 22272
rect 10466 21184 10474 21248
rect 10538 21184 10554 21248
rect 10618 21184 10634 21248
rect 10698 21184 10714 21248
rect 10778 21184 10786 21248
rect 10466 20160 10786 21184
rect 10466 20096 10474 20160
rect 10538 20096 10554 20160
rect 10618 20096 10634 20160
rect 10698 20096 10714 20160
rect 10778 20096 10786 20160
rect 10466 19072 10786 20096
rect 10466 19008 10474 19072
rect 10538 19008 10554 19072
rect 10618 19008 10634 19072
rect 10698 19008 10714 19072
rect 10778 19008 10786 19072
rect 10466 17984 10786 19008
rect 10466 17920 10474 17984
rect 10538 17920 10554 17984
rect 10618 17920 10634 17984
rect 10698 17920 10714 17984
rect 10778 17920 10786 17984
rect 10466 16896 10786 17920
rect 10466 16832 10474 16896
rect 10538 16832 10554 16896
rect 10618 16832 10634 16896
rect 10698 16832 10714 16896
rect 10778 16832 10786 16896
rect 10466 15808 10786 16832
rect 10466 15744 10474 15808
rect 10538 15744 10554 15808
rect 10618 15744 10634 15808
rect 10698 15744 10714 15808
rect 10778 15744 10786 15808
rect 10466 14720 10786 15744
rect 10466 14656 10474 14720
rect 10538 14656 10554 14720
rect 10618 14656 10634 14720
rect 10698 14656 10714 14720
rect 10778 14656 10786 14720
rect 10466 13632 10786 14656
rect 10466 13568 10474 13632
rect 10538 13568 10554 13632
rect 10618 13568 10634 13632
rect 10698 13568 10714 13632
rect 10778 13568 10786 13632
rect 10466 12544 10786 13568
rect 10466 12480 10474 12544
rect 10538 12480 10554 12544
rect 10618 12480 10634 12544
rect 10698 12480 10714 12544
rect 10778 12480 10786 12544
rect 10466 11456 10786 12480
rect 10466 11392 10474 11456
rect 10538 11392 10554 11456
rect 10618 11392 10634 11456
rect 10698 11392 10714 11456
rect 10778 11392 10786 11456
rect 10466 10368 10786 11392
rect 10466 10304 10474 10368
rect 10538 10304 10554 10368
rect 10618 10304 10634 10368
rect 10698 10304 10714 10368
rect 10778 10304 10786 10368
rect 10466 9280 10786 10304
rect 10466 9216 10474 9280
rect 10538 9216 10554 9280
rect 10618 9216 10634 9280
rect 10698 9216 10714 9280
rect 10778 9216 10786 9280
rect 10466 8192 10786 9216
rect 10466 8128 10474 8192
rect 10538 8128 10554 8192
rect 10618 8128 10634 8192
rect 10698 8128 10714 8192
rect 10778 8128 10786 8192
rect 10466 7104 10786 8128
rect 10466 7040 10474 7104
rect 10538 7040 10554 7104
rect 10618 7040 10634 7104
rect 10698 7040 10714 7104
rect 10778 7040 10786 7104
rect 10466 6016 10786 7040
rect 10466 5952 10474 6016
rect 10538 5952 10554 6016
rect 10618 5952 10634 6016
rect 10698 5952 10714 6016
rect 10778 5952 10786 6016
rect 10466 4928 10786 5952
rect 10466 4864 10474 4928
rect 10538 4864 10554 4928
rect 10618 4864 10634 4928
rect 10698 4864 10714 4928
rect 10778 4864 10786 4928
rect 10466 3840 10786 4864
rect 10466 3776 10474 3840
rect 10538 3776 10554 3840
rect 10618 3776 10634 3840
rect 10698 3776 10714 3840
rect 10778 3776 10786 3840
rect 10466 2752 10786 3776
rect 10466 2688 10474 2752
rect 10538 2688 10554 2752
rect 10618 2688 10634 2752
rect 10698 2688 10714 2752
rect 10778 2688 10786 2752
rect 10466 2128 10786 2688
rect 13640 27232 13960 27248
rect 13640 27168 13648 27232
rect 13712 27168 13728 27232
rect 13792 27168 13808 27232
rect 13872 27168 13888 27232
rect 13952 27168 13960 27232
rect 13640 26144 13960 27168
rect 13640 26080 13648 26144
rect 13712 26080 13728 26144
rect 13792 26080 13808 26144
rect 13872 26080 13888 26144
rect 13952 26080 13960 26144
rect 13640 25056 13960 26080
rect 13640 24992 13648 25056
rect 13712 24992 13728 25056
rect 13792 24992 13808 25056
rect 13872 24992 13888 25056
rect 13952 24992 13960 25056
rect 13640 23968 13960 24992
rect 13640 23904 13648 23968
rect 13712 23904 13728 23968
rect 13792 23904 13808 23968
rect 13872 23904 13888 23968
rect 13952 23904 13960 23968
rect 13640 22880 13960 23904
rect 13640 22816 13648 22880
rect 13712 22816 13728 22880
rect 13792 22816 13808 22880
rect 13872 22816 13888 22880
rect 13952 22816 13960 22880
rect 13640 21792 13960 22816
rect 13640 21728 13648 21792
rect 13712 21728 13728 21792
rect 13792 21728 13808 21792
rect 13872 21728 13888 21792
rect 13952 21728 13960 21792
rect 13640 20704 13960 21728
rect 13640 20640 13648 20704
rect 13712 20640 13728 20704
rect 13792 20640 13808 20704
rect 13872 20640 13888 20704
rect 13952 20640 13960 20704
rect 13640 19616 13960 20640
rect 13640 19552 13648 19616
rect 13712 19552 13728 19616
rect 13792 19552 13808 19616
rect 13872 19552 13888 19616
rect 13952 19552 13960 19616
rect 13640 18528 13960 19552
rect 13640 18464 13648 18528
rect 13712 18464 13728 18528
rect 13792 18464 13808 18528
rect 13872 18464 13888 18528
rect 13952 18464 13960 18528
rect 13640 17440 13960 18464
rect 13640 17376 13648 17440
rect 13712 17376 13728 17440
rect 13792 17376 13808 17440
rect 13872 17376 13888 17440
rect 13952 17376 13960 17440
rect 13640 16352 13960 17376
rect 13640 16288 13648 16352
rect 13712 16288 13728 16352
rect 13792 16288 13808 16352
rect 13872 16288 13888 16352
rect 13952 16288 13960 16352
rect 13640 15264 13960 16288
rect 13640 15200 13648 15264
rect 13712 15200 13728 15264
rect 13792 15200 13808 15264
rect 13872 15200 13888 15264
rect 13952 15200 13960 15264
rect 13640 14176 13960 15200
rect 13640 14112 13648 14176
rect 13712 14112 13728 14176
rect 13792 14112 13808 14176
rect 13872 14112 13888 14176
rect 13952 14112 13960 14176
rect 13640 13088 13960 14112
rect 13640 13024 13648 13088
rect 13712 13024 13728 13088
rect 13792 13024 13808 13088
rect 13872 13024 13888 13088
rect 13952 13024 13960 13088
rect 13640 12000 13960 13024
rect 13640 11936 13648 12000
rect 13712 11936 13728 12000
rect 13792 11936 13808 12000
rect 13872 11936 13888 12000
rect 13952 11936 13960 12000
rect 13640 10912 13960 11936
rect 13640 10848 13648 10912
rect 13712 10848 13728 10912
rect 13792 10848 13808 10912
rect 13872 10848 13888 10912
rect 13952 10848 13960 10912
rect 13640 9824 13960 10848
rect 13640 9760 13648 9824
rect 13712 9760 13728 9824
rect 13792 9760 13808 9824
rect 13872 9760 13888 9824
rect 13952 9760 13960 9824
rect 13640 8736 13960 9760
rect 13640 8672 13648 8736
rect 13712 8672 13728 8736
rect 13792 8672 13808 8736
rect 13872 8672 13888 8736
rect 13952 8672 13960 8736
rect 13640 7648 13960 8672
rect 13640 7584 13648 7648
rect 13712 7584 13728 7648
rect 13792 7584 13808 7648
rect 13872 7584 13888 7648
rect 13952 7584 13960 7648
rect 13640 6560 13960 7584
rect 13640 6496 13648 6560
rect 13712 6496 13728 6560
rect 13792 6496 13808 6560
rect 13872 6496 13888 6560
rect 13952 6496 13960 6560
rect 13640 5472 13960 6496
rect 13640 5408 13648 5472
rect 13712 5408 13728 5472
rect 13792 5408 13808 5472
rect 13872 5408 13888 5472
rect 13952 5408 13960 5472
rect 13640 4384 13960 5408
rect 13640 4320 13648 4384
rect 13712 4320 13728 4384
rect 13792 4320 13808 4384
rect 13872 4320 13888 4384
rect 13952 4320 13960 4384
rect 13640 3296 13960 4320
rect 13640 3232 13648 3296
rect 13712 3232 13728 3296
rect 13792 3232 13808 3296
rect 13872 3232 13888 3296
rect 13952 3232 13960 3296
rect 13640 2208 13960 3232
rect 13640 2144 13648 2208
rect 13712 2144 13728 2208
rect 13792 2144 13808 2208
rect 13872 2144 13888 2208
rect 13952 2144 13960 2208
rect 13640 2128 13960 2144
rect 16814 26688 17134 27248
rect 16814 26624 16822 26688
rect 16886 26624 16902 26688
rect 16966 26624 16982 26688
rect 17046 26624 17062 26688
rect 17126 26624 17134 26688
rect 16814 25600 17134 26624
rect 16814 25536 16822 25600
rect 16886 25536 16902 25600
rect 16966 25536 16982 25600
rect 17046 25536 17062 25600
rect 17126 25536 17134 25600
rect 16814 24512 17134 25536
rect 16814 24448 16822 24512
rect 16886 24448 16902 24512
rect 16966 24448 16982 24512
rect 17046 24448 17062 24512
rect 17126 24448 17134 24512
rect 16814 23424 17134 24448
rect 16814 23360 16822 23424
rect 16886 23360 16902 23424
rect 16966 23360 16982 23424
rect 17046 23360 17062 23424
rect 17126 23360 17134 23424
rect 16814 22336 17134 23360
rect 16814 22272 16822 22336
rect 16886 22272 16902 22336
rect 16966 22272 16982 22336
rect 17046 22272 17062 22336
rect 17126 22272 17134 22336
rect 16814 21248 17134 22272
rect 16814 21184 16822 21248
rect 16886 21184 16902 21248
rect 16966 21184 16982 21248
rect 17046 21184 17062 21248
rect 17126 21184 17134 21248
rect 16814 20160 17134 21184
rect 16814 20096 16822 20160
rect 16886 20096 16902 20160
rect 16966 20096 16982 20160
rect 17046 20096 17062 20160
rect 17126 20096 17134 20160
rect 16814 19072 17134 20096
rect 16814 19008 16822 19072
rect 16886 19008 16902 19072
rect 16966 19008 16982 19072
rect 17046 19008 17062 19072
rect 17126 19008 17134 19072
rect 16814 17984 17134 19008
rect 16814 17920 16822 17984
rect 16886 17920 16902 17984
rect 16966 17920 16982 17984
rect 17046 17920 17062 17984
rect 17126 17920 17134 17984
rect 16814 16896 17134 17920
rect 16814 16832 16822 16896
rect 16886 16832 16902 16896
rect 16966 16832 16982 16896
rect 17046 16832 17062 16896
rect 17126 16832 17134 16896
rect 16814 15808 17134 16832
rect 16814 15744 16822 15808
rect 16886 15744 16902 15808
rect 16966 15744 16982 15808
rect 17046 15744 17062 15808
rect 17126 15744 17134 15808
rect 16814 14720 17134 15744
rect 16814 14656 16822 14720
rect 16886 14656 16902 14720
rect 16966 14656 16982 14720
rect 17046 14656 17062 14720
rect 17126 14656 17134 14720
rect 16814 13632 17134 14656
rect 16814 13568 16822 13632
rect 16886 13568 16902 13632
rect 16966 13568 16982 13632
rect 17046 13568 17062 13632
rect 17126 13568 17134 13632
rect 16814 12544 17134 13568
rect 16814 12480 16822 12544
rect 16886 12480 16902 12544
rect 16966 12480 16982 12544
rect 17046 12480 17062 12544
rect 17126 12480 17134 12544
rect 16814 11456 17134 12480
rect 16814 11392 16822 11456
rect 16886 11392 16902 11456
rect 16966 11392 16982 11456
rect 17046 11392 17062 11456
rect 17126 11392 17134 11456
rect 16814 10368 17134 11392
rect 16814 10304 16822 10368
rect 16886 10304 16902 10368
rect 16966 10304 16982 10368
rect 17046 10304 17062 10368
rect 17126 10304 17134 10368
rect 16814 9280 17134 10304
rect 16814 9216 16822 9280
rect 16886 9216 16902 9280
rect 16966 9216 16982 9280
rect 17046 9216 17062 9280
rect 17126 9216 17134 9280
rect 16814 8192 17134 9216
rect 16814 8128 16822 8192
rect 16886 8128 16902 8192
rect 16966 8128 16982 8192
rect 17046 8128 17062 8192
rect 17126 8128 17134 8192
rect 16814 7104 17134 8128
rect 16814 7040 16822 7104
rect 16886 7040 16902 7104
rect 16966 7040 16982 7104
rect 17046 7040 17062 7104
rect 17126 7040 17134 7104
rect 16814 6016 17134 7040
rect 16814 5952 16822 6016
rect 16886 5952 16902 6016
rect 16966 5952 16982 6016
rect 17046 5952 17062 6016
rect 17126 5952 17134 6016
rect 16814 4928 17134 5952
rect 16814 4864 16822 4928
rect 16886 4864 16902 4928
rect 16966 4864 16982 4928
rect 17046 4864 17062 4928
rect 17126 4864 17134 4928
rect 16814 3840 17134 4864
rect 16814 3776 16822 3840
rect 16886 3776 16902 3840
rect 16966 3776 16982 3840
rect 17046 3776 17062 3840
rect 17126 3776 17134 3840
rect 16814 2752 17134 3776
rect 16814 2688 16822 2752
rect 16886 2688 16902 2752
rect 16966 2688 16982 2752
rect 17046 2688 17062 2752
rect 17126 2688 17134 2752
rect 16814 2128 17134 2688
rect 19988 27232 20308 27248
rect 19988 27168 19996 27232
rect 20060 27168 20076 27232
rect 20140 27168 20156 27232
rect 20220 27168 20236 27232
rect 20300 27168 20308 27232
rect 19988 26144 20308 27168
rect 19988 26080 19996 26144
rect 20060 26080 20076 26144
rect 20140 26080 20156 26144
rect 20220 26080 20236 26144
rect 20300 26080 20308 26144
rect 19988 25056 20308 26080
rect 19988 24992 19996 25056
rect 20060 24992 20076 25056
rect 20140 24992 20156 25056
rect 20220 24992 20236 25056
rect 20300 24992 20308 25056
rect 19988 23968 20308 24992
rect 19988 23904 19996 23968
rect 20060 23904 20076 23968
rect 20140 23904 20156 23968
rect 20220 23904 20236 23968
rect 20300 23904 20308 23968
rect 19988 22880 20308 23904
rect 19988 22816 19996 22880
rect 20060 22816 20076 22880
rect 20140 22816 20156 22880
rect 20220 22816 20236 22880
rect 20300 22816 20308 22880
rect 19988 21792 20308 22816
rect 19988 21728 19996 21792
rect 20060 21728 20076 21792
rect 20140 21728 20156 21792
rect 20220 21728 20236 21792
rect 20300 21728 20308 21792
rect 19988 20704 20308 21728
rect 19988 20640 19996 20704
rect 20060 20640 20076 20704
rect 20140 20640 20156 20704
rect 20220 20640 20236 20704
rect 20300 20640 20308 20704
rect 19988 19616 20308 20640
rect 19988 19552 19996 19616
rect 20060 19552 20076 19616
rect 20140 19552 20156 19616
rect 20220 19552 20236 19616
rect 20300 19552 20308 19616
rect 19988 18528 20308 19552
rect 19988 18464 19996 18528
rect 20060 18464 20076 18528
rect 20140 18464 20156 18528
rect 20220 18464 20236 18528
rect 20300 18464 20308 18528
rect 19988 17440 20308 18464
rect 19988 17376 19996 17440
rect 20060 17376 20076 17440
rect 20140 17376 20156 17440
rect 20220 17376 20236 17440
rect 20300 17376 20308 17440
rect 19988 16352 20308 17376
rect 19988 16288 19996 16352
rect 20060 16288 20076 16352
rect 20140 16288 20156 16352
rect 20220 16288 20236 16352
rect 20300 16288 20308 16352
rect 19988 15264 20308 16288
rect 19988 15200 19996 15264
rect 20060 15200 20076 15264
rect 20140 15200 20156 15264
rect 20220 15200 20236 15264
rect 20300 15200 20308 15264
rect 19988 14176 20308 15200
rect 19988 14112 19996 14176
rect 20060 14112 20076 14176
rect 20140 14112 20156 14176
rect 20220 14112 20236 14176
rect 20300 14112 20308 14176
rect 19988 13088 20308 14112
rect 19988 13024 19996 13088
rect 20060 13024 20076 13088
rect 20140 13024 20156 13088
rect 20220 13024 20236 13088
rect 20300 13024 20308 13088
rect 19988 12000 20308 13024
rect 19988 11936 19996 12000
rect 20060 11936 20076 12000
rect 20140 11936 20156 12000
rect 20220 11936 20236 12000
rect 20300 11936 20308 12000
rect 19988 10912 20308 11936
rect 19988 10848 19996 10912
rect 20060 10848 20076 10912
rect 20140 10848 20156 10912
rect 20220 10848 20236 10912
rect 20300 10848 20308 10912
rect 19988 9824 20308 10848
rect 19988 9760 19996 9824
rect 20060 9760 20076 9824
rect 20140 9760 20156 9824
rect 20220 9760 20236 9824
rect 20300 9760 20308 9824
rect 19988 8736 20308 9760
rect 19988 8672 19996 8736
rect 20060 8672 20076 8736
rect 20140 8672 20156 8736
rect 20220 8672 20236 8736
rect 20300 8672 20308 8736
rect 19988 7648 20308 8672
rect 19988 7584 19996 7648
rect 20060 7584 20076 7648
rect 20140 7584 20156 7648
rect 20220 7584 20236 7648
rect 20300 7584 20308 7648
rect 19988 6560 20308 7584
rect 19988 6496 19996 6560
rect 20060 6496 20076 6560
rect 20140 6496 20156 6560
rect 20220 6496 20236 6560
rect 20300 6496 20308 6560
rect 19988 5472 20308 6496
rect 19988 5408 19996 5472
rect 20060 5408 20076 5472
rect 20140 5408 20156 5472
rect 20220 5408 20236 5472
rect 20300 5408 20308 5472
rect 19988 4384 20308 5408
rect 19988 4320 19996 4384
rect 20060 4320 20076 4384
rect 20140 4320 20156 4384
rect 20220 4320 20236 4384
rect 20300 4320 20308 4384
rect 19988 3296 20308 4320
rect 19988 3232 19996 3296
rect 20060 3232 20076 3296
rect 20140 3232 20156 3296
rect 20220 3232 20236 3296
rect 20300 3232 20308 3296
rect 19988 2208 20308 3232
rect 19988 2144 19996 2208
rect 20060 2144 20076 2208
rect 20140 2144 20156 2208
rect 20220 2144 20236 2208
rect 20300 2144 20308 2208
rect 19988 2128 20308 2144
rect 23162 26688 23482 27248
rect 23162 26624 23170 26688
rect 23234 26624 23250 26688
rect 23314 26624 23330 26688
rect 23394 26624 23410 26688
rect 23474 26624 23482 26688
rect 23162 25600 23482 26624
rect 23162 25536 23170 25600
rect 23234 25536 23250 25600
rect 23314 25536 23330 25600
rect 23394 25536 23410 25600
rect 23474 25536 23482 25600
rect 23162 24512 23482 25536
rect 23162 24448 23170 24512
rect 23234 24448 23250 24512
rect 23314 24448 23330 24512
rect 23394 24448 23410 24512
rect 23474 24448 23482 24512
rect 23162 23424 23482 24448
rect 23162 23360 23170 23424
rect 23234 23360 23250 23424
rect 23314 23360 23330 23424
rect 23394 23360 23410 23424
rect 23474 23360 23482 23424
rect 23162 22336 23482 23360
rect 23162 22272 23170 22336
rect 23234 22272 23250 22336
rect 23314 22272 23330 22336
rect 23394 22272 23410 22336
rect 23474 22272 23482 22336
rect 23162 21248 23482 22272
rect 23162 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23482 21248
rect 23162 20160 23482 21184
rect 23162 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23482 20160
rect 23162 19072 23482 20096
rect 23162 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23482 19072
rect 23162 17984 23482 19008
rect 23162 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23482 17984
rect 23162 16896 23482 17920
rect 23162 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23482 16896
rect 23162 15808 23482 16832
rect 23162 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23482 15808
rect 23162 14720 23482 15744
rect 23162 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23482 14720
rect 23162 13632 23482 14656
rect 23162 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23482 13632
rect 23162 12544 23482 13568
rect 23162 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23482 12544
rect 23162 11456 23482 12480
rect 23162 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23482 11456
rect 23162 10368 23482 11392
rect 23162 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23482 10368
rect 23162 9280 23482 10304
rect 23162 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23482 9280
rect 23162 8192 23482 9216
rect 23162 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23482 8192
rect 23162 7104 23482 8128
rect 23162 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23482 7104
rect 23162 6016 23482 7040
rect 23162 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23482 6016
rect 23162 4928 23482 5952
rect 23162 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23482 4928
rect 23162 3840 23482 4864
rect 23162 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23482 3840
rect 23162 2752 23482 3776
rect 23162 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23482 2752
rect 23162 2128 23482 2688
rect 26336 27232 26656 27248
rect 26336 27168 26344 27232
rect 26408 27168 26424 27232
rect 26488 27168 26504 27232
rect 26568 27168 26584 27232
rect 26648 27168 26656 27232
rect 26336 26144 26656 27168
rect 26336 26080 26344 26144
rect 26408 26080 26424 26144
rect 26488 26080 26504 26144
rect 26568 26080 26584 26144
rect 26648 26080 26656 26144
rect 26336 25056 26656 26080
rect 26336 24992 26344 25056
rect 26408 24992 26424 25056
rect 26488 24992 26504 25056
rect 26568 24992 26584 25056
rect 26648 24992 26656 25056
rect 26336 23968 26656 24992
rect 26336 23904 26344 23968
rect 26408 23904 26424 23968
rect 26488 23904 26504 23968
rect 26568 23904 26584 23968
rect 26648 23904 26656 23968
rect 26336 22880 26656 23904
rect 26336 22816 26344 22880
rect 26408 22816 26424 22880
rect 26488 22816 26504 22880
rect 26568 22816 26584 22880
rect 26648 22816 26656 22880
rect 26336 21792 26656 22816
rect 26336 21728 26344 21792
rect 26408 21728 26424 21792
rect 26488 21728 26504 21792
rect 26568 21728 26584 21792
rect 26648 21728 26656 21792
rect 26336 20704 26656 21728
rect 26336 20640 26344 20704
rect 26408 20640 26424 20704
rect 26488 20640 26504 20704
rect 26568 20640 26584 20704
rect 26648 20640 26656 20704
rect 26336 19616 26656 20640
rect 26336 19552 26344 19616
rect 26408 19552 26424 19616
rect 26488 19552 26504 19616
rect 26568 19552 26584 19616
rect 26648 19552 26656 19616
rect 26336 18528 26656 19552
rect 26336 18464 26344 18528
rect 26408 18464 26424 18528
rect 26488 18464 26504 18528
rect 26568 18464 26584 18528
rect 26648 18464 26656 18528
rect 26336 17440 26656 18464
rect 26336 17376 26344 17440
rect 26408 17376 26424 17440
rect 26488 17376 26504 17440
rect 26568 17376 26584 17440
rect 26648 17376 26656 17440
rect 26336 16352 26656 17376
rect 26336 16288 26344 16352
rect 26408 16288 26424 16352
rect 26488 16288 26504 16352
rect 26568 16288 26584 16352
rect 26648 16288 26656 16352
rect 26336 15264 26656 16288
rect 26336 15200 26344 15264
rect 26408 15200 26424 15264
rect 26488 15200 26504 15264
rect 26568 15200 26584 15264
rect 26648 15200 26656 15264
rect 26336 14176 26656 15200
rect 26336 14112 26344 14176
rect 26408 14112 26424 14176
rect 26488 14112 26504 14176
rect 26568 14112 26584 14176
rect 26648 14112 26656 14176
rect 26336 13088 26656 14112
rect 26336 13024 26344 13088
rect 26408 13024 26424 13088
rect 26488 13024 26504 13088
rect 26568 13024 26584 13088
rect 26648 13024 26656 13088
rect 26336 12000 26656 13024
rect 26336 11936 26344 12000
rect 26408 11936 26424 12000
rect 26488 11936 26504 12000
rect 26568 11936 26584 12000
rect 26648 11936 26656 12000
rect 26336 10912 26656 11936
rect 26336 10848 26344 10912
rect 26408 10848 26424 10912
rect 26488 10848 26504 10912
rect 26568 10848 26584 10912
rect 26648 10848 26656 10912
rect 26336 9824 26656 10848
rect 26336 9760 26344 9824
rect 26408 9760 26424 9824
rect 26488 9760 26504 9824
rect 26568 9760 26584 9824
rect 26648 9760 26656 9824
rect 26336 8736 26656 9760
rect 26336 8672 26344 8736
rect 26408 8672 26424 8736
rect 26488 8672 26504 8736
rect 26568 8672 26584 8736
rect 26648 8672 26656 8736
rect 26336 7648 26656 8672
rect 26336 7584 26344 7648
rect 26408 7584 26424 7648
rect 26488 7584 26504 7648
rect 26568 7584 26584 7648
rect 26648 7584 26656 7648
rect 26336 6560 26656 7584
rect 26336 6496 26344 6560
rect 26408 6496 26424 6560
rect 26488 6496 26504 6560
rect 26568 6496 26584 6560
rect 26648 6496 26656 6560
rect 26336 5472 26656 6496
rect 26336 5408 26344 5472
rect 26408 5408 26424 5472
rect 26488 5408 26504 5472
rect 26568 5408 26584 5472
rect 26648 5408 26656 5472
rect 26336 4384 26656 5408
rect 26336 4320 26344 4384
rect 26408 4320 26424 4384
rect 26488 4320 26504 4384
rect 26568 4320 26584 4384
rect 26648 4320 26656 4384
rect 26336 3296 26656 4320
rect 26336 3232 26344 3296
rect 26408 3232 26424 3296
rect 26488 3232 26504 3296
rect 26568 3232 26584 3296
rect 26648 3232 26656 3296
rect 26336 2208 26656 3232
rect 26336 2144 26344 2208
rect 26408 2144 26424 2208
rect 26488 2144 26504 2208
rect 26568 2144 26584 2208
rect 26648 2144 26656 2208
rect 26336 2128 26656 2144
use sky130_fd_sc_hd__or3_1  _0521_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14996 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0522_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16468 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0523_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16468 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0524_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15456 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0525_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0526_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1688980957
transform 1 0 10488 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0528_
timestamp 1688980957
transform -1 0 12144 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0529_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14076 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1688980957
transform -1 0 11408 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0531_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11132 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_4  _0532_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10396 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _0533_
timestamp 1688980957
transform 1 0 12972 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1688980957
transform -1 0 15548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0535_
timestamp 1688980957
transform 1 0 12880 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0536_
timestamp 1688980957
transform 1 0 19228 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0537_
timestamp 1688980957
transform -1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1688980957
transform 1 0 3864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0539_
timestamp 1688980957
transform 1 0 4692 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0540_
timestamp 1688980957
transform 1 0 6808 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0541_
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0542_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0543_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0544_
timestamp 1688980957
transform 1 0 6532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0545_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0546_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14628 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0547_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10028 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1688980957
transform -1 0 8188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1688980957
transform -1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0550_
timestamp 1688980957
transform 1 0 5060 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0551_
timestamp 1688980957
transform -1 0 6072 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0552_
timestamp 1688980957
transform 1 0 4784 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0553_
timestamp 1688980957
transform -1 0 6440 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0554_
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0555_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0556_
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0557_
timestamp 1688980957
transform -1 0 15180 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0558_
timestamp 1688980957
transform 1 0 10120 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1688980957
transform -1 0 24288 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0560_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24196 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0561_
timestamp 1688980957
transform 1 0 22172 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0562_
timestamp 1688980957
transform -1 0 24288 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0563_
timestamp 1688980957
transform -1 0 23092 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0564_
timestamp 1688980957
transform 1 0 23092 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0565_
timestamp 1688980957
transform -1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0566_
timestamp 1688980957
transform -1 0 19872 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_2  _0567_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23920 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0568_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22264 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0569_
timestamp 1688980957
transform 1 0 21252 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0570_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0571_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24564 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0572_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25944 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0573_
timestamp 1688980957
transform -1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0574_
timestamp 1688980957
transform -1 0 21620 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0575_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20792 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0576_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21620 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1688980957
transform -1 0 16192 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0579_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0580_
timestamp 1688980957
transform -1 0 18308 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0581_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1688980957
transform -1 0 14996 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0583_
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0584_
timestamp 1688980957
transform -1 0 23920 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0585_
timestamp 1688980957
transform -1 0 22632 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0586_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0587_
timestamp 1688980957
transform -1 0 21620 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0588_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19872 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0589_
timestamp 1688980957
transform 1 0 10212 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0590_
timestamp 1688980957
transform -1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0591_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9752 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0592_
timestamp 1688980957
transform -1 0 11776 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0593_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0594_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0595_
timestamp 1688980957
transform -1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0596_
timestamp 1688980957
transform -1 0 9936 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1688980957
transform 1 0 9292 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0598_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10580 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0599_
timestamp 1688980957
transform 1 0 9936 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0600_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16284 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0601_
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0602_
timestamp 1688980957
transform 1 0 18216 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1688980957
transform 1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0604_
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0605_
timestamp 1688980957
transform -1 0 10488 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1688980957
transform -1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0607_
timestamp 1688980957
transform 1 0 11040 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0608_
timestamp 1688980957
transform -1 0 13064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0609_
timestamp 1688980957
transform -1 0 10120 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _0611_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18768 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0612_
timestamp 1688980957
transform -1 0 25116 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0613_
timestamp 1688980957
transform -1 0 23000 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0614_
timestamp 1688980957
transform -1 0 23828 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0615_
timestamp 1688980957
transform 1 0 22724 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0616_
timestamp 1688980957
transform 1 0 23184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0617_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0618_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _0619_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0620_
timestamp 1688980957
transform -1 0 16744 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0621_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1688980957
transform 1 0 16928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0623_
timestamp 1688980957
transform -1 0 15824 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _0624_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16928 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0625_
timestamp 1688980957
transform 1 0 12696 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0626_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14076 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0627_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13800 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_2  _0628_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19688 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0629_
timestamp 1688980957
transform 1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0630_
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0631_
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1688980957
transform -1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0633_
timestamp 1688980957
transform 1 0 15640 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0634_
timestamp 1688980957
transform -1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1688980957
transform 1 0 14260 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1688980957
transform -1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0637_
timestamp 1688980957
transform -1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1688980957
transform -1 0 21160 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1688980957
transform 1 0 15364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0641_
timestamp 1688980957
transform -1 0 15364 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1688980957
transform 1 0 6900 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1688980957
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0645_
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0646_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0647_
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _0648_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0649_
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0650_
timestamp 1688980957
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1688980957
transform -1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0652_
timestamp 1688980957
transform -1 0 13708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0653_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0654_
timestamp 1688980957
transform -1 0 13892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1688980957
transform 1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0656_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0657_
timestamp 1688980957
transform -1 0 17848 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0658_
timestamp 1688980957
transform 1 0 14904 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0659_
timestamp 1688980957
transform -1 0 25484 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0660_
timestamp 1688980957
transform -1 0 25300 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0661_
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _0662_
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0663_
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0664_
timestamp 1688980957
transform -1 0 23460 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0665_
timestamp 1688980957
transform 1 0 22540 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0666_
timestamp 1688980957
transform 1 0 17204 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0667_
timestamp 1688980957
transform 1 0 14904 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0668_
timestamp 1688980957
transform 1 0 12972 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0669_
timestamp 1688980957
transform 1 0 9936 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0670_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13984 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0671_
timestamp 1688980957
transform 1 0 13616 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1688980957
transform 1 0 14260 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0673_
timestamp 1688980957
transform -1 0 13616 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0674_
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0675_
timestamp 1688980957
transform 1 0 21160 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0676_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23184 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0677_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0678_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0679_
timestamp 1688980957
transform 1 0 21804 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0680_
timestamp 1688980957
transform -1 0 23644 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0681_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _0682_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0683_
timestamp 1688980957
transform 1 0 5336 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0685_
timestamp 1688980957
transform 1 0 4508 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0686_
timestamp 1688980957
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0687_
timestamp 1688980957
transform -1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0688_
timestamp 1688980957
transform 1 0 5796 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0689_
timestamp 1688980957
transform 1 0 7268 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _0690_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7360 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _0691_
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0692_
timestamp 1688980957
transform -1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 1688980957
transform -1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1688980957
transform 1 0 20148 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0696_
timestamp 1688980957
transform -1 0 19596 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0697_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0698_
timestamp 1688980957
transform 1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0699_
timestamp 1688980957
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0700_
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0701_
timestamp 1688980957
transform -1 0 17112 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0702_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0704_
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1688980957
transform -1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1688980957
transform 1 0 16192 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0708_
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1688980957
transform -1 0 13064 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0710_
timestamp 1688980957
transform 1 0 12328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1688980957
transform -1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0712_
timestamp 1688980957
transform -1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1688980957
transform 1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0714_
timestamp 1688980957
transform 1 0 10672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0715_
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1688980957
transform -1 0 19964 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0717_
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1688980957
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0719_
timestamp 1688980957
transform -1 0 19504 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0720_
timestamp 1688980957
transform -1 0 16652 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0721_
timestamp 1688980957
transform -1 0 14720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0722_
timestamp 1688980957
transform -1 0 17204 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0723_
timestamp 1688980957
transform -1 0 16560 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1688980957
transform 1 0 6900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0725_
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0726_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1688980957
transform -1 0 6716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0728_
timestamp 1688980957
transform -1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1688980957
transform 1 0 10488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0730_
timestamp 1688980957
transform -1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0731_
timestamp 1688980957
transform -1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0732_
timestamp 1688980957
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0733_
timestamp 1688980957
transform -1 0 21068 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0734_
timestamp 1688980957
transform -1 0 22264 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0735_
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0736_
timestamp 1688980957
transform -1 0 22632 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0737_
timestamp 1688980957
transform -1 0 20424 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0738_
timestamp 1688980957
transform 1 0 22908 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0739_
timestamp 1688980957
transform -1 0 22264 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0740_
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0741_
timestamp 1688980957
transform 1 0 22632 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0742_
timestamp 1688980957
transform -1 0 24104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0743_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0744_
timestamp 1688980957
transform 1 0 22356 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0745_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0746_
timestamp 1688980957
transform -1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0747_
timestamp 1688980957
transform -1 0 25208 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0748_
timestamp 1688980957
transform -1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0749_
timestamp 1688980957
transform 1 0 23276 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0750_
timestamp 1688980957
transform 1 0 23736 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0751_
timestamp 1688980957
transform -1 0 20884 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0752_
timestamp 1688980957
transform -1 0 21160 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0753_
timestamp 1688980957
transform -1 0 18584 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0754_
timestamp 1688980957
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0755_
timestamp 1688980957
transform -1 0 20516 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0756_
timestamp 1688980957
transform -1 0 19780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0757_
timestamp 1688980957
transform -1 0 19136 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0758_
timestamp 1688980957
transform 1 0 19780 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0759_
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _0760_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0761_
timestamp 1688980957
transform -1 0 21528 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0762_
timestamp 1688980957
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0763_
timestamp 1688980957
transform -1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0764_
timestamp 1688980957
transform -1 0 20884 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0765_
timestamp 1688980957
transform 1 0 20792 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0766_
timestamp 1688980957
transform -1 0 19596 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0768_
timestamp 1688980957
transform -1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0769_
timestamp 1688980957
transform -1 0 18032 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0770_
timestamp 1688980957
transform -1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0771_
timestamp 1688980957
transform 1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0772_
timestamp 1688980957
transform -1 0 17204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0773_
timestamp 1688980957
transform -1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0774_
timestamp 1688980957
transform -1 0 17388 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0775_
timestamp 1688980957
transform -1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0776_
timestamp 1688980957
transform -1 0 17848 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 1688980957
transform 1 0 11592 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0779_
timestamp 1688980957
transform -1 0 12328 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0780_
timestamp 1688980957
transform -1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 1688980957
transform -1 0 18032 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0782_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18676 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0783_
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0784_
timestamp 1688980957
transform 1 0 11592 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0785_
timestamp 1688980957
transform -1 0 14076 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0786_
timestamp 1688980957
transform 1 0 11776 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0787_
timestamp 1688980957
transform 1 0 15732 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0788_
timestamp 1688980957
transform 1 0 16192 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0789_
timestamp 1688980957
transform -1 0 14904 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0790_
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0791_
timestamp 1688980957
transform 1 0 17940 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0792_
timestamp 1688980957
transform -1 0 17204 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0793_
timestamp 1688980957
transform -1 0 17572 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0794_
timestamp 1688980957
transform -1 0 17020 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _0795_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16560 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1688980957
transform 1 0 13800 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0797_
timestamp 1688980957
transform -1 0 14720 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0798_
timestamp 1688980957
transform 1 0 15640 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0799_
timestamp 1688980957
transform 1 0 13524 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0800_
timestamp 1688980957
transform 1 0 14628 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0801_
timestamp 1688980957
transform -1 0 12972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0802_
timestamp 1688980957
transform 1 0 12420 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0803_
timestamp 1688980957
transform 1 0 12512 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0804_
timestamp 1688980957
transform 1 0 12880 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0805_
timestamp 1688980957
transform -1 0 13800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0806_
timestamp 1688980957
transform 1 0 12144 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0807_
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0808_
timestamp 1688980957
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0809_
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0810_
timestamp 1688980957
transform 1 0 9568 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0811_
timestamp 1688980957
transform -1 0 10120 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0812_
timestamp 1688980957
transform 1 0 7728 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0813_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1688980957
transform 1 0 10120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0815_
timestamp 1688980957
transform 1 0 10396 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0816_
timestamp 1688980957
transform -1 0 9752 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0817_
timestamp 1688980957
transform -1 0 10764 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1688980957
transform -1 0 9476 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0819_
timestamp 1688980957
transform 1 0 10948 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0820_
timestamp 1688980957
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0821_
timestamp 1688980957
transform -1 0 12420 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0822_
timestamp 1688980957
transform 1 0 13064 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0823_
timestamp 1688980957
transform 1 0 11960 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0824_
timestamp 1688980957
transform -1 0 16100 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 1688980957
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _0826_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16376 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0827_
timestamp 1688980957
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0828_
timestamp 1688980957
transform -1 0 8372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0829_
timestamp 1688980957
transform -1 0 4232 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0830_
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0831_
timestamp 1688980957
transform -1 0 5796 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0832_
timestamp 1688980957
transform 1 0 2668 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0833_
timestamp 1688980957
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0835_
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0836_
timestamp 1688980957
transform 1 0 4140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0837_
timestamp 1688980957
transform -1 0 4692 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1688980957
transform 1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0839_
timestamp 1688980957
transform 1 0 3496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0840_
timestamp 1688980957
transform 1 0 2944 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0841_
timestamp 1688980957
transform 1 0 2576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0842_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0843_
timestamp 1688980957
transform 1 0 3220 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0844_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0845_
timestamp 1688980957
transform -1 0 4232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0846_
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0847_
timestamp 1688980957
transform -1 0 4232 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 1688980957
transform 1 0 2668 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1688980957
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0850_
timestamp 1688980957
transform -1 0 4784 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0851_
timestamp 1688980957
transform -1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1688980957
transform -1 0 3680 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0853_
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0854_
timestamp 1688980957
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0855_
timestamp 1688980957
transform -1 0 4876 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0856_
timestamp 1688980957
transform 1 0 8004 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0857_
timestamp 1688980957
transform -1 0 3680 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0858_
timestamp 1688980957
transform -1 0 6072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0859_
timestamp 1688980957
transform -1 0 5796 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1688980957
transform 1 0 2300 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 1688980957
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0862_
timestamp 1688980957
transform -1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0863_
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0864_
timestamp 1688980957
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0865_
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0866_
timestamp 1688980957
transform 1 0 2300 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0867_
timestamp 1688980957
transform 1 0 3036 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0868_
timestamp 1688980957
transform -1 0 3680 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1688980957
transform 1 0 3772 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0870_
timestamp 1688980957
transform 1 0 2300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1688980957
transform 1 0 3220 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0872_
timestamp 1688980957
transform 1 0 3680 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1688980957
transform 1 0 3956 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0874_
timestamp 1688980957
transform -1 0 3220 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0875_
timestamp 1688980957
transform -1 0 4232 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 1688980957
transform 1 0 2576 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0877_
timestamp 1688980957
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0878_
timestamp 1688980957
transform 1 0 4416 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0879_
timestamp 1688980957
transform -1 0 5060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0880_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0881_
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0882_
timestamp 1688980957
transform 1 0 6348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1688980957
transform 1 0 4968 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1688980957
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0885_
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0886_
timestamp 1688980957
transform -1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0887_
timestamp 1688980957
transform 1 0 7360 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0888_
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0889_
timestamp 1688980957
transform 1 0 18308 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0890_
timestamp 1688980957
transform 1 0 23000 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0891_
timestamp 1688980957
transform 1 0 22172 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0892_
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 1688980957
transform 1 0 23184 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0894_
timestamp 1688980957
transform -1 0 23092 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0895_
timestamp 1688980957
transform -1 0 23184 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0896_
timestamp 1688980957
transform 1 0 21896 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0897_
timestamp 1688980957
transform 1 0 23092 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1688980957
transform 1 0 23828 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0899_
timestamp 1688980957
transform 1 0 23092 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0900_
timestamp 1688980957
transform -1 0 25116 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0901_
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1688980957
transform 1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0903_
timestamp 1688980957
transform 1 0 25116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1688980957
transform 1 0 25208 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1688980957
transform -1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0906_
timestamp 1688980957
transform -1 0 24288 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0907_
timestamp 1688980957
transform -1 0 26220 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1688980957
transform 1 0 24472 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0909_
timestamp 1688980957
transform -1 0 24288 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1688980957
transform 1 0 23276 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0912_
timestamp 1688980957
transform -1 0 25944 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0913_
timestamp 1688980957
transform -1 0 25116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0914_
timestamp 1688980957
transform 1 0 25024 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0915_
timestamp 1688980957
transform 1 0 23644 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 1688980957
transform 1 0 25208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0917_
timestamp 1688980957
transform -1 0 25024 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1688980957
transform -1 0 6440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0919_
timestamp 1688980957
transform 1 0 5704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0920_
timestamp 1688980957
transform -1 0 4416 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 1688980957
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1688980957
transform -1 0 8740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0923_
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0924_
timestamp 1688980957
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1688980957
transform -1 0 17940 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0926_
timestamp 1688980957
transform 1 0 18124 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0927_
timestamp 1688980957
transform 1 0 19688 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0928_
timestamp 1688980957
transform 1 0 17296 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0929_
timestamp 1688980957
transform -1 0 18952 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1688980957
transform 1 0 18768 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0931_
timestamp 1688980957
transform -1 0 12788 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0932_
timestamp 1688980957
transform 1 0 12052 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0933_
timestamp 1688980957
transform -1 0 12880 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1688980957
transform -1 0 12788 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0935_
timestamp 1688980957
transform 1 0 11960 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1688980957
transform -1 0 11040 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0938_
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0939_
timestamp 1688980957
transform 1 0 11960 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0940_
timestamp 1688980957
transform -1 0 11408 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0941_
timestamp 1688980957
transform -1 0 12420 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0942_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0943_
timestamp 1688980957
transform -1 0 9936 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1688980957
transform -1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1688980957
transform 1 0 9476 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0946_
timestamp 1688980957
transform 1 0 9016 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0947_
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0948_
timestamp 1688980957
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1688980957
transform 1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0950_
timestamp 1688980957
transform 1 0 7360 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 1688980957
transform -1 0 8280 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0952_
timestamp 1688980957
transform -1 0 8648 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0953_
timestamp 1688980957
transform -1 0 9476 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0954_
timestamp 1688980957
transform 1 0 8096 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0955_
timestamp 1688980957
transform -1 0 8832 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0956_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0957_
timestamp 1688980957
transform -1 0 8648 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp 1688980957
transform 1 0 7912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1688980957
transform -1 0 6624 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1688980957
transform -1 0 20516 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0961_
timestamp 1688980957
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0962_
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0963_
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0964_
timestamp 1688980957
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0965_
timestamp 1688980957
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0966_
timestamp 1688980957
transform -1 0 20700 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0967_
timestamp 1688980957
transform -1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0968_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0969_
timestamp 1688980957
transform -1 0 12696 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0970_
timestamp 1688980957
transform 1 0 12144 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0971_
timestamp 1688980957
transform -1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0972_
timestamp 1688980957
transform -1 0 11408 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 1688980957
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0974_
timestamp 1688980957
transform 1 0 17296 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2b_2  _0975_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0976_
timestamp 1688980957
transform 1 0 12328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1688980957
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0978_
timestamp 1688980957
transform -1 0 13984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0979_
timestamp 1688980957
transform -1 0 14904 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0980_
timestamp 1688980957
transform -1 0 13248 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0981_
timestamp 1688980957
transform 1 0 13432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0982_
timestamp 1688980957
transform 1 0 15640 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0983_
timestamp 1688980957
transform -1 0 15456 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1688980957
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0985_
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0986_
timestamp 1688980957
transform -1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1688980957
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0988_
timestamp 1688980957
transform 1 0 17940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0989_
timestamp 1688980957
transform 1 0 15456 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0990_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1688980957
transform -1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0992_
timestamp 1688980957
transform -1 0 17388 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0993_
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1688980957
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0995_
timestamp 1688980957
transform -1 0 18584 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0996_
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0997_
timestamp 1688980957
transform 1 0 17848 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0998_
timestamp 1688980957
transform 1 0 19504 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp 1688980957
transform -1 0 20056 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1688980957
transform 1 0 20148 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1688980957
transform 1 0 15180 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1002_
timestamp 1688980957
transform -1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1688980957
transform 1 0 15088 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1688980957
transform -1 0 15824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1005_
timestamp 1688980957
transform 1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1006_
timestamp 1688980957
transform -1 0 13248 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1007_
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1688980957
transform -1 0 19688 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1009_
timestamp 1688980957
transform -1 0 22172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1010_
timestamp 1688980957
transform -1 0 19412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1011_
timestamp 1688980957
transform 1 0 21160 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1013_
timestamp 1688980957
transform 1 0 23000 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1014_
timestamp 1688980957
transform -1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1015_
timestamp 1688980957
transform 1 0 22724 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1688980957
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1688980957
transform -1 0 23000 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1019_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1020_
timestamp 1688980957
transform 1 0 23092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1021_
timestamp 1688980957
transform -1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1022_
timestamp 1688980957
transform 1 0 22632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1023_
timestamp 1688980957
transform 1 0 25116 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1024_
timestamp 1688980957
transform -1 0 24564 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1688980957
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1026_
timestamp 1688980957
transform -1 0 24288 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1027_
timestamp 1688980957
transform -1 0 24840 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1028_
timestamp 1688980957
transform -1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1029_
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1030_
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1031_
timestamp 1688980957
transform 1 0 23276 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1032_
timestamp 1688980957
transform 1 0 23276 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1688980957
transform 1 0 23000 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1034_
timestamp 1688980957
transform -1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1035_
timestamp 1688980957
transform 1 0 23552 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1036_
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1037_
timestamp 1688980957
transform 1 0 23184 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1038_
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1039_
timestamp 1688980957
transform 1 0 22632 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1040_
timestamp 1688980957
transform -1 0 25300 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1688980957
transform 1 0 25300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1042_
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1044_
timestamp 1688980957
transform 1 0 16928 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1688980957
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1046_
timestamp 1688980957
transform 1 0 15364 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1688980957
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1688980957
transform 1 0 8004 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1688980957
transform 1 0 8004 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1688980957
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1052_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1053_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10120 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1054_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8740 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1055_
timestamp 1688980957
transform -1 0 9752 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1056_
timestamp 1688980957
transform 1 0 8924 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1057_
timestamp 1688980957
transform -1 0 10120 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1058_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22724 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1688980957
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1688980957
transform 1 0 24564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1688980957
transform 1 0 22172 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1688980957
transform 1 0 18308 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1688980957
transform 1 0 18584 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1688980957
transform -1 0 23276 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1688980957
transform 1 0 21344 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1688980957
transform 1 0 19596 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1688980957
transform 1 0 16836 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1688980957
transform 1 0 16836 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1688980957
transform 1 0 17020 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1074_
timestamp 1688980957
transform 1 0 10212 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1075_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1688980957
transform 1 0 18216 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1688980957
transform 1 0 14720 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1688980957
transform -1 0 18124 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1688980957
transform 1 0 16468 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1688980957
transform 1 0 14352 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1688980957
transform 1 0 12052 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1688980957
transform 1 0 10580 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1688980957
transform 1 0 7360 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1688980957
transform 1 0 8004 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1688980957
transform -1 0 13064 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1688980957
transform 1 0 11592 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1089_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1090_
timestamp 1688980957
transform -1 0 21344 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1688980957
transform -1 0 21344 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1093_
timestamp 1688980957
transform 1 0 9200 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1094_
timestamp 1688980957
transform 1 0 7636 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 1688980957
transform -1 0 11132 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1096_
timestamp 1688980957
transform 1 0 9108 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 1688980957
transform 1 0 6716 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1098_
timestamp 1688980957
transform -1 0 8464 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1099_
timestamp 1688980957
transform 1 0 4784 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1100_
timestamp 1688980957
transform 1 0 1472 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1101_
timestamp 1688980957
transform 1 0 4692 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1688980957
transform 1 0 2760 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1103_
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1688980957
transform 1 0 1840 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 1688980957
transform 1 0 4140 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 1688980957
transform -1 0 10396 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1110_
timestamp 1688980957
transform 1 0 13616 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1688980957
transform 1 0 14168 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1688980957
transform 1 0 12052 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 1688980957
transform -1 0 15916 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1688980957
transform 1 0 14444 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1688980957
transform 1 0 16744 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1688980957
transform 1 0 14720 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1688980957
transform 1 0 8188 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1688980957
transform -1 0 9016 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1121_
timestamp 1688980957
transform 1 0 6624 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1122_
timestamp 1688980957
transform 1 0 1564 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1123_
timestamp 1688980957
transform 1 0 4692 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1124_
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1688980957
transform 1 0 1472 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1688980957
transform 1 0 4692 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1131_
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1132_
timestamp 1688980957
transform -1 0 8188 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1133_
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 1688980957
transform 1 0 17112 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1135_
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1136_
timestamp 1688980957
transform 1 0 23092 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1137_
timestamp 1688980957
transform -1 0 22172 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1138_
timestamp 1688980957
transform 1 0 23276 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1139_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1140_
timestamp 1688980957
transform 1 0 24288 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1141_
timestamp 1688980957
transform 1 0 22448 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 1688980957
transform 1 0 22632 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1143_
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 1688980957
transform 1 0 19596 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 1688980957
transform -1 0 8372 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1147_
timestamp 1688980957
transform 1 0 2392 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1148_
timestamp 1688980957
transform 1 0 8004 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1149_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1150_
timestamp 1688980957
transform 1 0 17572 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1151_
timestamp 1688980957
transform 1 0 17572 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1688980957
transform -1 0 11408 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1153_
timestamp 1688980957
transform 1 0 11316 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 1688980957
transform 1 0 11040 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1155_
timestamp 1688980957
transform -1 0 14444 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1156_
timestamp 1688980957
transform 1 0 11040 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 1688980957
transform 1 0 8648 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1688980957
transform 1 0 8004 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1688980957
transform 1 0 7636 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1688980957
transform 1 0 6072 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1688980957
transform 1 0 10396 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 1688980957
transform 1 0 10396 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1164_
timestamp 1688980957
transform 1 0 18952 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1165_
timestamp 1688980957
transform 1 0 19136 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1166_
timestamp 1688980957
transform 1 0 20516 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1167_
timestamp 1688980957
transform -1 0 17572 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1688980957
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 1688980957
transform -1 0 19412 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1688980957
transform 1 0 16192 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1688980957
transform 1 0 11224 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1688980957
transform 1 0 9384 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1175_
timestamp 1688980957
transform 1 0 14260 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1176_
timestamp 1688980957
transform 1 0 10672 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1177_
timestamp 1688980957
transform -1 0 13616 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1178_
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 1688980957
transform 1 0 14536 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1688980957
transform -1 0 17296 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1181_
timestamp 1688980957
transform 1 0 17296 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1688980957
transform 1 0 17296 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1688980957
transform -1 0 20424 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1688980957
transform 1 0 12420 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1688980957
transform -1 0 16284 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1688980957
transform -1 0 16284 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1188_
timestamp 1688980957
transform 1 0 11592 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 1688980957
transform 1 0 19412 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1688980957
transform 1 0 19596 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1191_
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1192_
timestamp 1688980957
transform 1 0 20608 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1193_
timestamp 1688980957
transform 1 0 20608 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1194_
timestamp 1688980957
transform 1 0 22172 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1688980957
transform 1 0 23736 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1197_
timestamp 1688980957
transform 1 0 22540 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1198_
timestamp 1688980957
transform 1 0 23828 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1199_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1200_
timestamp 1688980957
transform 1 0 20608 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1688980957
transform 1 0 17848 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 1688980957
transform 1 0 17296 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1203_
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 1688980957
transform 1 0 13524 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 1688980957
transform 1 0 7360 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 1688980957
transform 1 0 6992 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13800 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7360 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform -1 0 11960 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 10396 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform -1 0 6256 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 10488 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform 1 0 9844 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform -1 0 18768 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 17940 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform 1 0 21620 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 15824 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform -1 0 16376 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform 1 0 21344 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 21344 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_23 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_24
timestamp 1688980957
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_25
timestamp 1688980957
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_26
timestamp 1688980957
transform 1 0 25944 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_27
timestamp 1688980957
transform -1 0 11316 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_28
timestamp 1688980957
transform -1 0 15180 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cnn_kws_accel_29
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout7
timestamp 1688980957
transform -1 0 4048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout8
timestamp 1688980957
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 1688980957
transform 1 0 10396 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout10
timestamp 1688980957
transform 1 0 8832 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout11
timestamp 1688980957
transform -1 0 3312 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout13
timestamp 1688980957
transform -1 0 10212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1688980957
transform -1 0 3680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout16
timestamp 1688980957
transform 1 0 23092 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1688980957
transform -1 0 22172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1688980957
transform -1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1688980957
transform 1 0 14444 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1688980957
transform -1 0 13984 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 1688980957
transform 1 0 21068 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1688980957
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_95 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_104 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_147
timestamp 1688980957
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_159
timestamp 1688980957
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_14 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_38
timestamp 1688980957
transform 1 0 4600 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_42
timestamp 1688980957
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1688980957
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_106
timestamp 1688980957
transform 1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_145
timestamp 1688980957
transform 1 0 14444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_155
timestamp 1688980957
transform 1 0 15364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_159
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_163
timestamp 1688980957
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_177
timestamp 1688980957
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_210
timestamp 1688980957
transform 1 0 20424 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_218
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_222
timestamp 1688980957
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_252
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_264
timestamp 1688980957
transform 1 0 25392 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_272
timestamp 1688980957
transform 1 0 26128 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1688980957
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_60
timestamp 1688980957
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_103
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_174
timestamp 1688980957
transform 1 0 17112 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_206
timestamp 1688980957
transform 1 0 20056 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_235
timestamp 1688980957
transform 1 0 22724 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_243
timestamp 1688980957
transform 1 0 23460 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_268
timestamp 1688980957
transform 1 0 25760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_272
timestamp 1688980957
transform 1 0 26128 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_61
timestamp 1688980957
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_107
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_136
timestamp 1688980957
transform 1 0 13616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_182
timestamp 1688980957
transform 1 0 17848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_190
timestamp 1688980957
transform 1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_210
timestamp 1688980957
transform 1 0 20424 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_222
timestamp 1688980957
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_266
timestamp 1688980957
transform 1 0 25576 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_272
timestamp 1688980957
transform 1 0 26128 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_25
timestamp 1688980957
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_39
timestamp 1688980957
transform 1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_62
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_98
timestamp 1688980957
transform 1 0 10120 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_110
timestamp 1688980957
transform 1 0 11224 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_169
timestamp 1688980957
transform 1 0 16652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_206
timestamp 1688980957
transform 1 0 20056 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_238
timestamp 1688980957
transform 1 0 23000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_266
timestamp 1688980957
transform 1 0 25576 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_272
timestamp 1688980957
transform 1 0 26128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_32
timestamp 1688980957
transform 1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_37
timestamp 1688980957
transform 1 0 4508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_50
timestamp 1688980957
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_79
timestamp 1688980957
transform 1 0 8372 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_84
timestamp 1688980957
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_96
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_108
timestamp 1688980957
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_139
timestamp 1688980957
transform 1 0 13892 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_147
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_175
timestamp 1688980957
transform 1 0 17204 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_197
timestamp 1688980957
transform 1 0 19228 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_208
timestamp 1688980957
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_220
timestamp 1688980957
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_243
timestamp 1688980957
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_247
timestamp 1688980957
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_255
timestamp 1688980957
transform 1 0 24564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_267
timestamp 1688980957
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_19
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_34
timestamp 1688980957
transform 1 0 4232 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_42
timestamp 1688980957
transform 1 0 4968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_58
timestamp 1688980957
transform 1 0 6440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_80
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_96
timestamp 1688980957
transform 1 0 9936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_108
timestamp 1688980957
transform 1 0 11040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_115
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_122
timestamp 1688980957
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_148
timestamp 1688980957
transform 1 0 14720 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_182
timestamp 1688980957
transform 1 0 17848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_227
timestamp 1688980957
transform 1 0 21988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_244
timestamp 1688980957
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_261
timestamp 1688980957
transform 1 0 25116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_29
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_45
timestamp 1688980957
transform 1 0 5244 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_61
timestamp 1688980957
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_141
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_150
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_156
timestamp 1688980957
transform 1 0 15456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_219
timestamp 1688980957
transform 1 0 21252 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_247
timestamp 1688980957
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_43
timestamp 1688980957
transform 1 0 5060 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_51
timestamp 1688980957
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_63
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_71
timestamp 1688980957
transform 1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_94
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_98
timestamp 1688980957
transform 1 0 10120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_173
timestamp 1688980957
transform 1 0 17020 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_229
timestamp 1688980957
transform 1 0 22172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_235
timestamp 1688980957
transform 1 0 22724 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_14
timestamp 1688980957
transform 1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_32
timestamp 1688980957
transform 1 0 4048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_65
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_76
timestamp 1688980957
transform 1 0 8096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_80
timestamp 1688980957
transform 1 0 8464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_107
timestamp 1688980957
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_164
timestamp 1688980957
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_208
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_233
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_243
timestamp 1688980957
transform 1 0 23460 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_263
timestamp 1688980957
transform 1 0 25300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_271
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_7
timestamp 1688980957
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_105
timestamp 1688980957
transform 1 0 10764 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_118
timestamp 1688980957
transform 1 0 11960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_130
timestamp 1688980957
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_202
timestamp 1688980957
transform 1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_243
timestamp 1688980957
transform 1 0 23460 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_23
timestamp 1688980957
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_43
timestamp 1688980957
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_94
timestamp 1688980957
transform 1 0 9752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_133
timestamp 1688980957
transform 1 0 13340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_189
timestamp 1688980957
transform 1 0 18492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_201
timestamp 1688980957
transform 1 0 19596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_206
timestamp 1688980957
transform 1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_212
timestamp 1688980957
transform 1 0 20608 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_233
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_268
timestamp 1688980957
transform 1 0 25760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_272
timestamp 1688980957
transform 1 0 26128 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_19
timestamp 1688980957
transform 1 0 2852 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_68
timestamp 1688980957
transform 1 0 7360 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_107
timestamp 1688980957
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_134
timestamp 1688980957
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_150
timestamp 1688980957
transform 1 0 14904 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_230
timestamp 1688980957
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_23
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_46
timestamp 1688980957
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1688980957
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_73
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_98
timestamp 1688980957
transform 1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_153
timestamp 1688980957
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1688980957
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_177
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_202
timestamp 1688980957
transform 1 0 19688 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_230
timestamp 1688980957
transform 1 0 22264 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_271
timestamp 1688980957
transform 1 0 26036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_24
timestamp 1688980957
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_39
timestamp 1688980957
transform 1 0 4692 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_61
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_76
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_89
timestamp 1688980957
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_149
timestamp 1688980957
transform 1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_156
timestamp 1688980957
transform 1 0 15456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_163
timestamp 1688980957
transform 1 0 16100 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_172
timestamp 1688980957
transform 1 0 16928 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_184
timestamp 1688980957
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1688980957
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_208
timestamp 1688980957
transform 1 0 20240 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_214
timestamp 1688980957
transform 1 0 20792 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_246
timestamp 1688980957
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_259
timestamp 1688980957
transform 1 0 24932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_266
timestamp 1688980957
transform 1 0 25576 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_272
timestamp 1688980957
transform 1 0 26128 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_14
timestamp 1688980957
transform 1 0 2392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_25
timestamp 1688980957
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_31
timestamp 1688980957
transform 1 0 3956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_62
timestamp 1688980957
transform 1 0 6808 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_72
timestamp 1688980957
transform 1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_96
timestamp 1688980957
transform 1 0 9936 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_104
timestamp 1688980957
transform 1 0 10672 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1688980957
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_119
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_124
timestamp 1688980957
transform 1 0 12512 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_136
timestamp 1688980957
transform 1 0 13616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_142
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_175
timestamp 1688980957
transform 1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_212
timestamp 1688980957
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_236
timestamp 1688980957
transform 1 0 22816 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_248
timestamp 1688980957
transform 1 0 23920 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_260
timestamp 1688980957
transform 1 0 25024 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_272
timestamp 1688980957
transform 1 0 26128 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_34
timestamp 1688980957
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_54
timestamp 1688980957
transform 1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_60
timestamp 1688980957
transform 1 0 6624 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_72
timestamp 1688980957
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_94
timestamp 1688980957
transform 1 0 9752 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_106
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_118
timestamp 1688980957
transform 1 0 11960 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_130
timestamp 1688980957
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_170
timestamp 1688980957
transform 1 0 16744 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_183
timestamp 1688980957
transform 1 0 17940 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_192
timestamp 1688980957
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_220
timestamp 1688980957
transform 1 0 21344 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_234
timestamp 1688980957
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_246
timestamp 1688980957
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_43
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1688980957
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_130
timestamp 1688980957
transform 1 0 13064 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 1688980957
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_177
timestamp 1688980957
transform 1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_215
timestamp 1688980957
transform 1 0 20884 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_219
timestamp 1688980957
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_233
timestamp 1688980957
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_254
timestamp 1688980957
transform 1 0 24472 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_266
timestamp 1688980957
transform 1 0 25576 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_272
timestamp 1688980957
transform 1 0 26128 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_33
timestamp 1688980957
transform 1 0 4140 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_66
timestamp 1688980957
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_78
timestamp 1688980957
transform 1 0 8280 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_117
timestamp 1688980957
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_132
timestamp 1688980957
transform 1 0 13248 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_145
timestamp 1688980957
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_205
timestamp 1688980957
transform 1 0 19964 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_11
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_28
timestamp 1688980957
transform 1 0 3680 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_32
timestamp 1688980957
transform 1 0 4048 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1688980957
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_63
timestamp 1688980957
transform 1 0 6900 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_78
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_84
timestamp 1688980957
transform 1 0 8832 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_88
timestamp 1688980957
transform 1 0 9200 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_134
timestamp 1688980957
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_157
timestamp 1688980957
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1688980957
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_191
timestamp 1688980957
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_203
timestamp 1688980957
transform 1 0 19780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_229
timestamp 1688980957
transform 1 0 22172 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_37
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_67
timestamp 1688980957
transform 1 0 7268 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_101
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_145
timestamp 1688980957
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_157
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_204
timestamp 1688980957
transform 1 0 19872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_208
timestamp 1688980957
transform 1 0 20240 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_212
timestamp 1688980957
transform 1 0 20608 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_218
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_230
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_238
timestamp 1688980957
transform 1 0 23000 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_244
timestamp 1688980957
transform 1 0 23552 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_11
timestamp 1688980957
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_28
timestamp 1688980957
transform 1 0 3680 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_36
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_65
timestamp 1688980957
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_86
timestamp 1688980957
transform 1 0 9016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_108
timestamp 1688980957
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_116
timestamp 1688980957
transform 1 0 11776 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_177
timestamp 1688980957
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_199
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_232
timestamp 1688980957
transform 1 0 22448 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_245
timestamp 1688980957
transform 1 0 23644 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_252
timestamp 1688980957
transform 1 0 24288 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_45
timestamp 1688980957
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_49
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_69
timestamp 1688980957
transform 1 0 7452 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_104
timestamp 1688980957
transform 1 0 10672 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_116
timestamp 1688980957
transform 1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1688980957
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_151
timestamp 1688980957
transform 1 0 14996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_200
timestamp 1688980957
transform 1 0 19504 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_206
timestamp 1688980957
transform 1 0 20056 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_267
timestamp 1688980957
transform 1 0 25668 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_28
timestamp 1688980957
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_40
timestamp 1688980957
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 1688980957
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_61
timestamp 1688980957
transform 1 0 6716 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_67
timestamp 1688980957
transform 1 0 7268 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_158
timestamp 1688980957
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_173
timestamp 1688980957
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_194
timestamp 1688980957
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_221
timestamp 1688980957
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_245
timestamp 1688980957
transform 1 0 23644 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_6
timestamp 1688980957
transform 1 0 1656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_10
timestamp 1688980957
transform 1 0 2024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_14
timestamp 1688980957
transform 1 0 2392 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_50
timestamp 1688980957
transform 1 0 5704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_54
timestamp 1688980957
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_135
timestamp 1688980957
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_161
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_167
timestamp 1688980957
transform 1 0 16468 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_171
timestamp 1688980957
transform 1 0 16836 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_181
timestamp 1688980957
transform 1 0 17756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_223
timestamp 1688980957
transform 1 0 21620 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_236
timestamp 1688980957
transform 1 0 22816 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_248
timestamp 1688980957
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_260
timestamp 1688980957
transform 1 0 25024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_272
timestamp 1688980957
transform 1 0 26128 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_28
timestamp 1688980957
transform 1 0 3680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_91
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_117
timestamp 1688980957
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_126
timestamp 1688980957
transform 1 0 12696 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_208
timestamp 1688980957
transform 1 0 20240 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_220
timestamp 1688980957
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_242
timestamp 1688980957
transform 1 0 23368 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_79
timestamp 1688980957
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_130
timestamp 1688980957
transform 1 0 13064 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_161
timestamp 1688980957
transform 1 0 15916 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_184
timestamp 1688980957
transform 1 0 18032 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_210
timestamp 1688980957
transform 1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_224
timestamp 1688980957
transform 1 0 21712 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_272
timestamp 1688980957
transform 1 0 26128 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_11
timestamp 1688980957
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_42
timestamp 1688980957
transform 1 0 4968 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_66
timestamp 1688980957
transform 1 0 7176 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_78
timestamp 1688980957
transform 1 0 8280 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_90
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_102
timestamp 1688980957
transform 1 0 10488 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_116
timestamp 1688980957
transform 1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_127
timestamp 1688980957
transform 1 0 12788 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_135
timestamp 1688980957
transform 1 0 13524 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_143
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_189
timestamp 1688980957
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_222
timestamp 1688980957
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_240
timestamp 1688980957
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_262
timestamp 1688980957
transform 1 0 25208 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_271
timestamp 1688980957
transform 1 0 26036 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_60
timestamp 1688980957
transform 1 0 6624 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_72
timestamp 1688980957
transform 1 0 7728 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_82
timestamp 1688980957
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_88
timestamp 1688980957
transform 1 0 9200 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_94
timestamp 1688980957
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_99
timestamp 1688980957
transform 1 0 10212 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_128
timestamp 1688980957
transform 1 0 12880 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_151
timestamp 1688980957
transform 1 0 14996 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_163
timestamp 1688980957
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_175
timestamp 1688980957
transform 1 0 17204 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 1688980957
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_205
timestamp 1688980957
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_14
timestamp 1688980957
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_26
timestamp 1688980957
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_38
timestamp 1688980957
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_50
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_123
timestamp 1688980957
transform 1 0 12420 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_141
timestamp 1688980957
transform 1 0 14076 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_156
timestamp 1688980957
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_216
timestamp 1688980957
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_262
timestamp 1688980957
transform 1 0 25208 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_270
timestamp 1688980957
transform 1 0 25944 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_113
timestamp 1688980957
transform 1 0 11500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_117
timestamp 1688980957
transform 1 0 11868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_211
timestamp 1688980957
transform 1 0 20516 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_223
timestamp 1688980957
transform 1 0 21620 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_235
timestamp 1688980957
transform 1 0 22724 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_239
timestamp 1688980957
transform 1 0 23092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_9
timestamp 1688980957
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_21
timestamp 1688980957
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_33
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_45
timestamp 1688980957
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_60
timestamp 1688980957
transform 1 0 6624 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_91
timestamp 1688980957
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_124
timestamp 1688980957
transform 1 0 12512 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_199
timestamp 1688980957
transform 1 0 19412 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_220
timestamp 1688980957
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_231
timestamp 1688980957
transform 1 0 22356 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_236
timestamp 1688980957
transform 1 0 22816 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_248
timestamp 1688980957
transform 1 0 23920 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_260
timestamp 1688980957
transform 1 0 25024 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_272
timestamp 1688980957
transform 1 0 26128 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_82
timestamp 1688980957
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_94
timestamp 1688980957
transform 1 0 9752 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_106
timestamp 1688980957
transform 1 0 10856 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_137
timestamp 1688980957
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_171
timestamp 1688980957
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_225
timestamp 1688980957
transform 1 0 21804 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_65
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_106
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_122
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_128
timestamp 1688980957
transform 1 0 12880 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_141
timestamp 1688980957
transform 1 0 14076 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_160
timestamp 1688980957
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_173
timestamp 1688980957
transform 1 0 17020 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_198
timestamp 1688980957
transform 1 0 19320 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_206
timestamp 1688980957
transform 1 0 20056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_218
timestamp 1688980957
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_262
timestamp 1688980957
transform 1 0 25208 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_270
timestamp 1688980957
transform 1 0 25944 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_73
timestamp 1688980957
transform 1 0 7820 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_101
timestamp 1688980957
transform 1 0 10396 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_128
timestamp 1688980957
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_166
timestamp 1688980957
transform 1 0 16376 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_183
timestamp 1688980957
transform 1 0 17940 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_191
timestamp 1688980957
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_217
timestamp 1688980957
transform 1 0 21068 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_248
timestamp 1688980957
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_269
timestamp 1688980957
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_91
timestamp 1688980957
transform 1 0 9476 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_103
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_119
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_123
timestamp 1688980957
transform 1 0 12420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_135
timestamp 1688980957
transform 1 0 13524 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_143
timestamp 1688980957
transform 1 0 14260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_164
timestamp 1688980957
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_172
timestamp 1688980957
transform 1 0 16928 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_191
timestamp 1688980957
transform 1 0 18676 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_203
timestamp 1688980957
transform 1 0 19780 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_210
timestamp 1688980957
transform 1 0 20424 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_218
timestamp 1688980957
transform 1 0 21160 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_254
timestamp 1688980957
transform 1 0 24472 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_270
timestamp 1688980957
transform 1 0 25944 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_91
timestamp 1688980957
transform 1 0 9476 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_103
timestamp 1688980957
transform 1 0 10580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_111
timestamp 1688980957
transform 1 0 11316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_147
timestamp 1688980957
transform 1 0 14628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_169
timestamp 1688980957
transform 1 0 16652 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_231
timestamp 1688980957
transform 1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_240
timestamp 1688980957
transform 1 0 23184 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_246
timestamp 1688980957
transform 1 0 23736 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1688980957
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_259
timestamp 1688980957
transform 1 0 24932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_270
timestamp 1688980957
transform 1 0 25944 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_162
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_271
timestamp 1688980957
transform 1 0 26036 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_108
timestamp 1688980957
transform 1 0 11040 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_116
timestamp 1688980957
transform 1 0 11776 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_126
timestamp 1688980957
transform 1 0 12696 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_147
timestamp 1688980957
transform 1 0 14628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_159
timestamp 1688980957
transform 1 0 15732 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_169
timestamp 1688980957
transform 1 0 16652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_175
timestamp 1688980957
transform 1 0 17204 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_180
timestamp 1688980957
transform 1 0 17664 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_191
timestamp 1688980957
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_205
timestamp 1688980957
transform 1 0 19964 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1688980957
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_264
timestamp 1688980957
transform 1 0 25392 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_272
timestamp 1688980957
transform 1 0 26128 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_101
timestamp 1688980957
transform 1 0 10396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_109
timestamp 1688980957
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_148
timestamp 1688980957
transform 1 0 14720 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_157
timestamp 1688980957
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_165
timestamp 1688980957
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_203
timestamp 1688980957
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_215
timestamp 1688980957
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_234
timestamp 1688980957
transform 1 0 22632 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_259
timestamp 1688980957
transform 1 0 24932 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_271
timestamp 1688980957
transform 1 0 26036 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_103
timestamp 1688980957
transform 1 0 10580 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_115
timestamp 1688980957
transform 1 0 11684 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_122
timestamp 1688980957
transform 1 0 12328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_129
timestamp 1688980957
transform 1 0 12972 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_150
timestamp 1688980957
transform 1 0 14904 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_158
timestamp 1688980957
transform 1 0 15640 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_164
timestamp 1688980957
transform 1 0 16192 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_176
timestamp 1688980957
transform 1 0 17296 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_188
timestamp 1688980957
transform 1 0 18400 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_192
timestamp 1688980957
transform 1 0 18768 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_210
timestamp 1688980957
transform 1 0 20424 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_222
timestamp 1688980957
transform 1 0 21528 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_234
timestamp 1688980957
transform 1 0 22632 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_244
timestamp 1688980957
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_269
timestamp 1688980957
transform 1 0 25852 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_106
timestamp 1688980957
transform 1 0 10856 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_141
timestamp 1688980957
transform 1 0 14076 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_179
timestamp 1688980957
transform 1 0 17572 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_234
timestamp 1688980957
transform 1 0 22632 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_246
timestamp 1688980957
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_258
timestamp 1688980957
transform 1 0 24840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_270
timestamp 1688980957
transform 1 0 25944 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_186
timestamp 1688980957
transform 1 0 18216 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_218
timestamp 1688980957
transform 1 0 21160 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_236
timestamp 1688980957
transform 1 0 22816 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_248
timestamp 1688980957
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_141
timestamp 1688980957
transform 1 0 14076 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1688980957
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_185
timestamp 1688980957
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_189
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1688980957
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_241
timestamp 1688980957
transform 1 0 23276 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_253
timestamp 1688980957
transform 1 0 24380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_265
timestamp 1688980957
transform 1 0 25484 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_92
timestamp 1688980957
transform 1 0 9568 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_104
timestamp 1688980957
transform 1 0 10672 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_113
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_127
timestamp 1688980957
transform 1 0 12788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_157
timestamp 1688980957
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_186
timestamp 1688980957
transform 1 0 18216 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1688980957
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_236
timestamp 1688980957
transform 1 0 22816 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_248
timestamp 1688980957
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_6
timestamp 1688980957
transform 1 0 1656 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_18
timestamp 1688980957
transform 1 0 2760 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_26
timestamp 1688980957
transform 1 0 3496 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_29
timestamp 1688980957
transform 1 0 3772 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_34
timestamp 1688980957
transform 1 0 4232 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_46
timestamp 1688980957
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 1688980957
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_85
timestamp 1688980957
transform 1 0 8924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_97
timestamp 1688980957
transform 1 0 10028 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_141
timestamp 1688980957
transform 1 0 14076 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_153
timestamp 1688980957
transform 1 0 15180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_165
timestamp 1688980957
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_173
timestamp 1688980957
transform 1 0 17020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_185
timestamp 1688980957
transform 1 0 18124 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_197
timestamp 1688980957
transform 1 0 19228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_209
timestamp 1688980957
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_213
timestamp 1688980957
transform 1 0 20700 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_233
timestamp 1688980957
transform 1 0 22540 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_245
timestamp 1688980957
transform 1 0 23644 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_251
timestamp 1688980957
transform 1 0 24196 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_253
timestamp 1688980957
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_265
timestamp 1688980957
transform 1 0 25484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21804 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 20148 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 21620 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 13984 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 12788 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 9844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 22448 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 12696 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 14904 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 14168 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 8096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 11500 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 22448 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 24748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 19320 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 22540 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 15916 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 15732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 10764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 9476 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 25944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 12236 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 13524 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 4784 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 3680 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 25116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 25484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 4692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 18216 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 17848 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 20516 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 16284 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform -1 0 15272 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 22540 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 19964 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 10764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 6256 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 6808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 7544 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 26220 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 15456 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 14444 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 21712 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 9108 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 5060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 19044 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 17940 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 20884 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform -1 0 22540 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 26220 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform -1 0 16284 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform -1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 3956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 24932 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 16744 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 19044 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 17572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 8096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 23736 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 17572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 9936 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 6440 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 16376 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 23092 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 22908 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 20700 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 19780 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 4968 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 6624 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform -1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 15824 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 13800 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 14076 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform -1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform -1 0 15088 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform 1 0 14168 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform -1 0 13708 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform -1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 22540 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 25300 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform -1 0 13432 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 19504 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 18492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform -1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform -1 0 19688 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform -1 0 21528 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform -1 0 13340 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 10028 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform -1 0 23184 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 8832 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 10948 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 10488 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform -1 0 10580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform -1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 17112 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 8280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform -1 0 19964 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 25116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform -1 0 4968 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform -1 0 21252 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform 1 0 25300 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform -1 0 25116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform -1 0 12788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform -1 0 10396 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 26128 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 18676 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 9660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform -1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 20148 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform -1 0 21436 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 25944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output3
timestamp 1688980957
transform 1 0 25668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1688980957
transform -1 0 1932 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 26496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 26496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 26496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 26496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 26496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 26496 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 26496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 26496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 26496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 26496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 26496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 26496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 26496 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 26496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 26496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 26496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 26496 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 26496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 26496 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 26496 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 26496 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 26496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 26496 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 26496 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 26496 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 26496 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 26496 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 26496 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 26496 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 26496 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 26496 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 26496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 26496 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 26496 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 26496 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 26496 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 26496 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 26496 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 26496 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 26496 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 26496 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 26496 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 26496 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 26496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 8832 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 13984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 19136 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 24288 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire6
timestamp 1688980957
transform -1 0 15088 0 1 7616
box -38 -48 314 592
<< labels >>
flabel metal3 s 26841 19728 27641 19848 0 FreeSans 480 0 0 0 audio_sample[0]
port 0 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 audio_sample[10]
port 1 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 audio_sample[11]
port 2 nsew signal input
flabel metal3 s 26841 16328 27641 16448 0 FreeSans 480 0 0 0 audio_sample[12]
port 3 nsew signal input
flabel metal2 s 18050 28985 18106 29785 0 FreeSans 224 90 0 0 audio_sample[13]
port 4 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 audio_sample[14]
port 5 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 audio_sample[15]
port 6 nsew signal input
flabel metal3 s 26841 27888 27641 28008 0 FreeSans 480 0 0 0 audio_sample[1]
port 7 nsew signal input
flabel metal2 s 21914 28985 21970 29785 0 FreeSans 224 90 0 0 audio_sample[2]
port 8 nsew signal input
flabel metal3 s 26841 8848 27641 8968 0 FreeSans 480 0 0 0 audio_sample[3]
port 9 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 audio_sample[4]
port 10 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 audio_sample[5]
port 11 nsew signal input
flabel metal2 s 25778 28985 25834 29785 0 FreeSans 224 90 0 0 audio_sample[6]
port 12 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 audio_sample[7]
port 13 nsew signal input
flabel metal2 s 7746 28985 7802 29785 0 FreeSans 224 90 0 0 audio_sample[8]
port 14 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 audio_sample[9]
port 15 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 clk
port 16 nsew signal input
flabel metal3 s 26841 688 27641 808 0 FreeSans 480 0 0 0 done
port 17 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 psram_ce_n
port 18 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 psram_d[0]
port 19 nsew signal bidirectional
flabel metal2 s 3882 28985 3938 29785 0 FreeSans 224 90 0 0 psram_d[1]
port 20 nsew signal bidirectional
flabel metal3 s 26841 4768 27641 4888 0 FreeSans 480 0 0 0 psram_d[2]
port 21 nsew signal bidirectional
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 psram_d[3]
port 22 nsew signal bidirectional
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 psram_douten[0]
port 23 nsew signal tristate
flabel metal3 s 26841 23808 27641 23928 0 FreeSans 480 0 0 0 psram_douten[1]
port 24 nsew signal tristate
flabel metal2 s 10966 28985 11022 29785 0 FreeSans 224 90 0 0 psram_douten[2]
port 25 nsew signal tristate
flabel metal2 s 14830 28985 14886 29785 0 FreeSans 224 90 0 0 psram_douten[3]
port 26 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 psram_sck
port 27 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 rst_n
port 28 nsew signal input
flabel metal2 s 18 28985 74 29785 0 FreeSans 224 90 0 0 sample_valid
port 29 nsew signal input
flabel metal3 s 26841 12248 27641 12368 0 FreeSans 480 0 0 0 start
port 30 nsew signal input
flabel metal4 s 4118 2128 4438 27248 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 10466 2128 10786 27248 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 16814 2128 17134 27248 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 23162 2128 23482 27248 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 7292 2128 7612 27248 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 13640 2128 13960 27248 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 19988 2128 20308 27248 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 26336 2128 26656 27248 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
rlabel metal1 13800 26656 13800 26656 0 vccd1
rlabel via1 13880 27200 13880 27200 0 vssd1
rlabel metal1 9568 5882 9568 5882 0 _0000_
rlabel metal1 9936 4182 9936 4182 0 _0001_
rlabel metal1 9108 12954 9108 12954 0 _0002_
rlabel metal1 6808 15402 6808 15402 0 _0003_
rlabel metal1 19182 13838 19182 13838 0 _0004_
rlabel metal1 17703 16762 17703 16762 0 _0005_
rlabel via1 12367 14586 12367 14586 0 _0006_
rlabel metal1 15088 16626 15088 16626 0 _0007_
rlabel metal1 16774 22678 16774 22678 0 _0008_
rlabel metal1 14842 21930 14842 21930 0 _0009_
rlabel metal1 9476 8942 9476 8942 0 _0010_
rlabel metal1 9936 2482 9936 2482 0 _0011_
rlabel metal1 10810 9044 10810 9044 0 _0012_
rlabel metal1 10764 11662 10764 11662 0 _0013_
rlabel metal2 10442 15351 10442 15351 0 _0014_
rlabel metal1 10442 12750 10442 12750 0 _0015_
rlabel metal1 16376 13838 16376 13838 0 _0016_
rlabel metal1 18216 17646 18216 17646 0 _0017_
rlabel metal1 18216 12750 18216 12750 0 _0018_
rlabel metal1 13110 13362 13110 13362 0 _0019_
rlabel metal1 12972 15674 12972 15674 0 _0020_
rlabel metal1 14904 12410 14904 12410 0 _0021_
rlabel viali 22494 22613 22494 22613 0 _0022_
rlabel metal2 19826 22406 19826 22406 0 _0023_
rlabel metal1 15410 22746 15410 22746 0 _0024_
rlabel metal2 9982 25670 9982 25670 0 _0025_
rlabel metal2 9338 26044 9338 26044 0 _0026_
rlabel metal2 12374 6154 12374 6154 0 _0027_
rlabel metal1 14858 20434 14858 20434 0 _0028_
rlabel metal1 19964 16558 19964 16558 0 _0029_
rlabel metal1 6624 15946 6624 15946 0 _0030_
rlabel metal2 7958 5712 7958 5712 0 _0031_
rlabel metal1 5658 7310 5658 7310 0 _0032_
rlabel metal2 7038 11900 7038 11900 0 _0033_
rlabel metal1 20286 13838 20286 13838 0 _0034_
rlabel metal1 11684 13362 11684 13362 0 _0035_
rlabel metal1 16100 6970 16100 6970 0 _0036_
rlabel metal1 20838 8534 20838 8534 0 _0037_
rlabel metal1 19642 19278 19642 19278 0 _0038_
rlabel metal1 21160 9690 21160 9690 0 _0039_
rlabel metal1 22898 23698 22898 23698 0 _0040_
rlabel metal1 22816 22134 22816 22134 0 _0041_
rlabel metal2 24886 22406 24886 22406 0 _0042_
rlabel metal2 22126 20910 22126 20910 0 _0043_
rlabel metal1 22627 19754 22627 19754 0 _0044_
rlabel metal1 24462 20910 24462 20910 0 _0045_
rlabel via1 18625 24854 18625 24854 0 _0046_
rlabel metal1 19320 24378 19320 24378 0 _0047_
rlabel metal1 19085 25942 19085 25942 0 _0048_
rlabel metal1 21482 26792 21482 26792 0 _0049_
rlabel metal1 21236 25194 21236 25194 0 _0050_
rlabel metal1 19672 19754 19672 19754 0 _0051_
rlabel metal1 17245 21930 17245 21930 0 _0052_
rlabel metal1 17199 19414 17199 19414 0 _0053_
rlabel via1 17337 18734 17337 18734 0 _0054_
rlabel via1 17705 19822 17705 19822 0 _0055_
rlabel metal2 11178 6698 11178 6698 0 _0056_
rlabel metal1 11730 5882 11730 5882 0 _0057_
rlabel metal1 19228 23154 19228 23154 0 _0058_
rlabel metal1 14076 22202 14076 22202 0 _0059_
rlabel metal1 14934 25194 14934 25194 0 _0060_
rlabel metal1 17342 24922 17342 24922 0 _0061_
rlabel viali 16785 25262 16785 25262 0 _0062_
rlabel metal2 14674 24582 14674 24582 0 _0063_
rlabel metal2 12650 25738 12650 25738 0 _0064_
rlabel metal1 11035 25194 11035 25194 0 _0065_
rlabel metal2 7774 23970 7774 23970 0 _0066_
rlabel metal1 8781 23698 8781 23698 0 _0067_
rlabel metal2 9338 22406 9338 22406 0 _0068_
rlabel metal1 12328 21658 12328 21658 0 _0069_
rlabel metal1 11955 22678 11955 22678 0 _0070_
rlabel metal1 15778 7752 15778 7752 0 _0071_
rlabel metal1 8924 5338 8924 5338 0 _0072_
rlabel metal1 1978 3162 1978 3162 0 _0073_
rlabel via1 5007 3706 5007 3706 0 _0074_
rlabel metal1 3082 3128 3082 3128 0 _0075_
rlabel metal1 2231 5134 2231 5134 0 _0076_
rlabel metal1 2484 6222 2484 6222 0 _0077_
rlabel metal1 1932 7514 1932 7514 0 _0078_
rlabel metal1 3588 8330 3588 8330 0 _0079_
rlabel metal1 4600 7446 4600 7446 0 _0080_
rlabel metal1 8142 13498 8142 13498 0 _0081_
rlabel metal1 2024 15674 2024 15674 0 _0082_
rlabel metal2 5014 13532 5014 13532 0 _0083_
rlabel metal1 2392 14042 2392 14042 0 _0084_
rlabel metal1 2024 12954 2024 12954 0 _0085_
rlabel metal1 1925 11322 1925 11322 0 _0086_
rlabel metal1 1971 10234 1971 10234 0 _0087_
rlabel metal1 4554 10166 4554 10166 0 _0088_
rlabel metal1 5375 10234 5375 10234 0 _0089_
rlabel metal2 7682 4284 7682 4284 0 _0090_
rlabel metal1 7176 7786 7176 7786 0 _0091_
rlabel metal1 18308 14382 18308 14382 0 _0092_
rlabel metal1 23368 18326 23368 18326 0 _0093_
rlabel metal1 22126 17306 22126 17306 0 _0094_
rlabel metal1 23368 16762 23368 16762 0 _0095_
rlabel metal1 25070 16762 25070 16762 0 _0096_
rlabel metal1 24564 15062 24564 15062 0 _0097_
rlabel metal1 23184 13158 23184 13158 0 _0098_
rlabel metal1 23322 11662 23322 11662 0 _0099_
rlabel metal1 24288 13158 24288 13158 0 _0100_
rlabel metal1 6256 16218 6256 16218 0 _0101_
rlabel metal2 3266 16932 3266 16932 0 _0102_
rlabel metal2 8326 10846 8326 10846 0 _0103_
rlabel metal1 19596 11186 19596 11186 0 _0104_
rlabel metal2 17894 10948 17894 10948 0 _0105_
rlabel metal1 18630 9146 18630 9146 0 _0106_
rlabel metal2 12742 16286 12742 16286 0 _0107_
rlabel metal1 11362 20808 11362 20808 0 _0108_
rlabel metal1 12972 18938 12972 18938 0 _0109_
rlabel metal1 11592 19414 11592 19414 0 _0110_
rlabel metal1 9016 18326 9016 18326 0 _0111_
rlabel metal1 8142 20366 8142 20366 0 _0112_
rlabel metal1 8004 20026 8004 20026 0 _0113_
rlabel metal1 6394 18632 6394 18632 0 _0114_
rlabel metal1 6624 18326 6624 18326 0 _0115_
rlabel metal2 18906 17476 18906 17476 0 _0116_
rlabel metal1 19596 18326 19596 18326 0 _0117_
rlabel metal1 20746 12750 20746 12750 0 _0118_
rlabel metal1 11914 8602 11914 8602 0 _0119_
rlabel metal1 11730 8330 11730 8330 0 _0120_
rlabel metal1 10350 10098 10350 10098 0 _0121_
rlabel metal1 11086 3162 11086 3162 0 _0122_
rlabel metal1 15180 4046 15180 4046 0 _0123_
rlabel metal1 12650 2958 12650 2958 0 _0124_
rlabel metal1 14766 2890 14766 2890 0 _0125_
rlabel metal1 16836 5338 16836 5338 0 _0126_
rlabel metal1 17526 4794 17526 4794 0 _0127_
rlabel metal1 18124 2618 18124 2618 0 _0128_
rlabel metal1 20102 3128 20102 3128 0 _0129_
rlabel metal1 14306 18258 14306 18258 0 _0130_
rlabel metal2 15962 19516 15962 19516 0 _0131_
rlabel metal1 12098 12410 12098 12410 0 _0132_
rlabel metal1 21850 6834 21850 6834 0 _0133_
rlabel metal1 19964 5338 19964 5338 0 _0134_
rlabel metal1 21114 3162 21114 3162 0 _0135_
rlabel metal1 21114 3570 21114 3570 0 _0136_
rlabel metal1 22494 3128 22494 3128 0 _0137_
rlabel metal1 24150 3706 24150 3706 0 _0138_
rlabel metal1 24472 6426 24472 6426 0 _0139_
rlabel metal1 22862 9656 22862 9656 0 _0140_
rlabel metal1 24288 8534 24288 8534 0 _0141_
rlabel metal1 25024 9010 25024 9010 0 _0142_
rlabel metal1 18952 7310 18952 7310 0 _0143_
rlabel metal1 17664 6698 17664 6698 0 _0144_
rlabel metal1 16744 15606 16744 15606 0 _0145_
rlabel metal1 13800 15674 13800 15674 0 _0146_
rlabel metal1 7728 14586 7728 14586 0 _0147_
rlabel metal2 8234 3264 8234 3264 0 _0148_
rlabel metal1 15502 14518 15502 14518 0 _0149_
rlabel metal1 15640 10030 15640 10030 0 _0150_
rlabel metal1 15272 9894 15272 9894 0 _0151_
rlabel metal2 11638 17442 11638 17442 0 _0152_
rlabel metal2 13110 18462 13110 18462 0 _0153_
rlabel metal1 11086 17646 11086 17646 0 _0154_
rlabel metal1 13386 18190 13386 18190 0 _0155_
rlabel metal1 8970 17680 8970 17680 0 _0156_
rlabel metal1 10764 17714 10764 17714 0 _0157_
rlabel metal1 12466 12274 12466 12274 0 _0158_
rlabel metal2 15410 13770 15410 13770 0 _0159_
rlabel metal1 20194 16116 20194 16116 0 _0160_
rlabel metal1 4508 12274 4508 12274 0 _0161_
rlabel metal1 5842 12342 5842 12342 0 _0162_
rlabel metal1 6210 13498 6210 13498 0 _0163_
rlabel metal1 6256 12682 6256 12682 0 _0164_
rlabel metal1 6164 12750 6164 12750 0 _0165_
rlabel metal1 6716 12206 6716 12206 0 _0166_
rlabel metal2 6670 16490 6670 16490 0 _0167_
rlabel metal1 16100 11118 16100 11118 0 _0168_
rlabel metal2 15318 11679 15318 11679 0 _0169_
rlabel via1 7866 9690 7866 9690 0 _0170_
rlabel metal1 4186 5678 4186 5678 0 _0171_
rlabel metal1 5704 5338 5704 5338 0 _0172_
rlabel metal1 5750 4794 5750 4794 0 _0173_
rlabel metal1 5382 6222 5382 6222 0 _0174_
rlabel metal1 5750 5882 5750 5882 0 _0175_
rlabel metal1 6210 6324 6210 6324 0 _0176_
rlabel metal1 5980 7378 5980 7378 0 _0177_
rlabel metal2 24058 17000 24058 17000 0 _0178_
rlabel metal1 23414 14960 23414 14960 0 _0179_
rlabel metal1 22954 15538 22954 15538 0 _0180_
rlabel metal1 23644 13906 23644 13906 0 _0181_
rlabel metal2 22678 15844 22678 15844 0 _0182_
rlabel metal1 23782 14416 23782 14416 0 _0183_
rlabel metal1 18860 16558 18860 16558 0 _0184_
rlabel metal1 22816 20910 22816 20910 0 _0185_
rlabel metal1 21758 24650 21758 24650 0 _0186_
rlabel metal1 21942 24684 21942 24684 0 _0187_
rlabel metal1 21574 21556 21574 21556 0 _0188_
rlabel metal1 24242 21658 24242 21658 0 _0189_
rlabel metal1 25438 21658 25438 21658 0 _0190_
rlabel metal1 24150 21998 24150 21998 0 _0191_
rlabel metal1 21712 21658 21712 21658 0 _0192_
rlabel metal2 10350 24191 10350 24191 0 _0193_
rlabel metal1 15962 22746 15962 22746 0 _0194_
rlabel metal2 18032 21522 18032 21522 0 _0195_
rlabel metal1 17526 21658 17526 21658 0 _0196_
rlabel metal1 18216 21658 18216 21658 0 _0197_
rlabel metal1 9752 23834 9752 23834 0 _0198_
rlabel metal1 22954 22746 22954 22746 0 _0199_
rlabel metal1 22783 22678 22783 22678 0 _0200_
rlabel metal1 21390 22576 21390 22576 0 _0201_
rlabel metal1 20424 21930 20424 21930 0 _0202_
rlabel metal1 10212 14518 10212 14518 0 _0203_
rlabel metal1 10856 23290 10856 23290 0 _0204_
rlabel metal1 10810 24242 10810 24242 0 _0205_
rlabel metal1 12098 24650 12098 24650 0 _0206_
rlabel metal1 10810 24820 10810 24820 0 _0207_
rlabel metal2 10626 25024 10626 25024 0 _0208_
rlabel metal2 9522 25908 9522 25908 0 _0209_
rlabel metal1 10580 24582 10580 24582 0 _0210_
rlabel metal1 7774 12886 7774 12886 0 _0211_
rlabel metal1 16560 14042 16560 14042 0 _0212_
rlabel metal1 11362 8330 11362 8330 0 _0213_
rlabel metal1 13018 7922 13018 7922 0 _0214_
rlabel metal2 9706 4998 9706 4998 0 _0215_
rlabel metal1 20194 10710 20194 10710 0 _0216_
rlabel metal1 22954 5644 22954 5644 0 _0217_
rlabel metal1 22678 5338 22678 5338 0 _0218_
rlabel metal1 22770 5712 22770 5712 0 _0219_
rlabel metal1 23184 5678 23184 5678 0 _0220_
rlabel metal1 21482 9554 21482 9554 0 _0221_
rlabel metal1 20194 8602 20194 8602 0 _0222_
rlabel metal1 19826 11866 19826 11866 0 _0223_
rlabel via1 15612 10642 15612 10642 0 _0224_
rlabel metal2 20930 12614 20930 12614 0 _0225_
rlabel metal2 19918 11356 19918 11356 0 _0226_
rlabel metal1 17158 10438 17158 10438 0 _0227_
rlabel metal1 14030 11764 14030 11764 0 _0228_
rlabel metal2 16146 8194 16146 8194 0 _0229_
rlabel metal2 13294 9146 13294 9146 0 _0230_
rlabel metal1 14076 9418 14076 9418 0 _0231_
rlabel metal1 19550 10642 19550 10642 0 _0232_
rlabel metal1 18216 10030 18216 10030 0 _0233_
rlabel viali 15315 10642 15315 10642 0 _0234_
rlabel metal2 15502 9894 15502 9894 0 _0235_
rlabel metal1 20470 12138 20470 12138 0 _0236_
rlabel metal1 15778 10676 15778 10676 0 _0237_
rlabel metal1 14950 10778 14950 10778 0 _0238_
rlabel metal1 14352 9010 14352 9010 0 _0239_
rlabel metal2 17158 3264 17158 3264 0 _0240_
rlabel metal1 15318 9418 15318 9418 0 _0241_
rlabel metal1 15594 12104 15594 12104 0 _0242_
rlabel metal1 15364 11118 15364 11118 0 _0243_
rlabel metal1 9430 11220 9430 11220 0 _0244_
rlabel metal1 8188 10778 8188 10778 0 _0245_
rlabel metal1 2553 18258 2553 18258 0 _0246_
rlabel metal1 5658 4250 5658 4250 0 _0247_
rlabel metal2 6394 3978 6394 3978 0 _0248_
rlabel metal1 5014 4794 5014 4794 0 _0249_
rlabel metal1 5888 5542 5888 5542 0 _0250_
rlabel metal1 13294 4692 13294 4692 0 _0251_
rlabel metal1 12926 4590 12926 4590 0 _0252_
rlabel metal1 13018 3400 13018 3400 0 _0253_
rlabel metal1 14030 4794 14030 4794 0 _0254_
rlabel metal1 14674 2618 14674 2618 0 _0255_
rlabel metal1 14030 4998 14030 4998 0 _0256_
rlabel metal2 15502 4624 15502 4624 0 _0257_
rlabel metal1 15088 4794 15088 4794 0 _0258_
rlabel metal1 16974 4250 16974 4250 0 _0259_
rlabel metal1 15042 5338 15042 5338 0 _0260_
rlabel metal1 24610 6222 24610 6222 0 _0261_
rlabel metal1 24380 6834 24380 6834 0 _0262_
rlabel metal2 17618 7072 17618 7072 0 _0263_
rlabel metal1 22862 5848 22862 5848 0 _0264_
rlabel metal1 22770 6222 22770 6222 0 _0265_
rlabel metal1 23046 6324 23046 6324 0 _0266_
rlabel metal1 18584 7514 18584 7514 0 _0267_
rlabel metal2 17802 7820 17802 7820 0 _0268_
rlabel metal2 14950 10166 14950 10166 0 _0269_
rlabel metal1 13662 18802 13662 18802 0 _0270_
rlabel metal1 13064 18802 13064 18802 0 _0271_
rlabel metal2 14260 15470 14260 15470 0 _0272_
rlabel metal1 14260 18054 14260 18054 0 _0273_
rlabel metal1 13386 18292 13386 18292 0 _0274_
rlabel metal2 13478 16524 13478 16524 0 _0275_
rlabel metal1 14858 11764 14858 11764 0 _0276_
rlabel metal2 21666 16983 21666 16983 0 _0277_
rlabel metal1 22540 16694 22540 16694 0 _0278_
rlabel metal1 22080 16626 22080 16626 0 _0279_
rlabel metal1 22466 16626 22466 16626 0 _0280_
rlabel metal1 21390 12784 21390 12784 0 _0281_
rlabel metal1 21206 12750 21206 12750 0 _0282_
rlabel metal2 20746 12517 20746 12517 0 _0283_
rlabel metal2 14674 11016 14674 11016 0 _0284_
rlabel metal1 5934 12206 5934 12206 0 _0285_
rlabel metal1 5106 12852 5106 12852 0 _0286_
rlabel metal1 4922 13974 4922 13974 0 _0287_
rlabel viali 4817 12818 4817 12818 0 _0288_
rlabel metal1 5474 12614 5474 12614 0 _0289_
rlabel metal2 7774 11186 7774 11186 0 _0290_
rlabel metal1 6486 8908 6486 8908 0 _0291_
rlabel metal1 8004 6766 8004 6766 0 _0292_
rlabel metal2 4462 16490 4462 16490 0 _0293_
rlabel metal1 19780 14586 19780 14586 0 _0294_
rlabel metal1 11316 14994 11316 14994 0 _0295_
rlabel metal2 16146 4896 16146 4896 0 _0296_
rlabel via2 14490 3349 14490 3349 0 _0297_
rlabel metal2 16698 3638 16698 3638 0 _0298_
rlabel metal1 16238 6800 16238 6800 0 _0299_
rlabel metal1 13892 5678 13892 5678 0 _0300_
rlabel metal2 20378 7990 20378 7990 0 _0301_
rlabel metal1 14214 17204 14214 17204 0 _0302_
rlabel metal2 12558 15776 12558 15776 0 _0303_
rlabel metal1 8142 5236 8142 5236 0 _0304_
rlabel metal1 10810 3162 10810 3162 0 _0305_
rlabel metal1 19826 16592 19826 16592 0 _0306_
rlabel metal2 18814 14858 18814 14858 0 _0307_
rlabel metal2 16192 22508 16192 22508 0 _0308_
rlabel metal1 16514 22610 16514 22610 0 _0309_
rlabel metal2 6486 15742 6486 15742 0 _0310_
rlabel metal1 9246 13294 9246 13294 0 _0311_
rlabel metal1 21252 9486 21252 9486 0 _0312_
rlabel metal1 21666 9350 21666 9350 0 _0313_
rlabel metal1 22034 23664 22034 23664 0 _0314_
rlabel metal2 19918 21835 19918 21835 0 _0315_
rlabel metal1 22218 23732 22218 23732 0 _0316_
rlabel metal1 23598 22066 23598 22066 0 _0317_
rlabel metal1 24610 21964 24610 21964 0 _0318_
rlabel metal2 22034 21318 22034 21318 0 _0319_
rlabel metal1 22770 19278 22770 19278 0 _0320_
rlabel metal1 23552 20502 23552 20502 0 _0321_
rlabel metal2 23966 21046 23966 21046 0 _0322_
rlabel metal2 20930 24276 20930 24276 0 _0323_
rlabel metal2 21114 26418 21114 26418 0 _0324_
rlabel viali 18829 25262 18829 25262 0 _0325_
rlabel metal1 19918 25738 19918 25738 0 _0326_
rlabel metal1 19274 24174 19274 24174 0 _0327_
rlabel metal1 19734 24378 19734 24378 0 _0328_
rlabel metal1 21298 26826 21298 26826 0 _0329_
rlabel metal1 21390 26962 21390 26962 0 _0330_
rlabel metal2 22494 26078 22494 26078 0 _0331_
rlabel metal1 20194 19822 20194 19822 0 _0332_
rlabel metal2 17710 22338 17710 22338 0 _0333_
rlabel via2 17250 21403 17250 21403 0 _0334_
rlabel metal1 17334 19686 17334 19686 0 _0335_
rlabel metal1 19274 19176 19274 19176 0 _0336_
rlabel metal1 17434 20910 17434 20910 0 _0337_
rlabel metal1 16974 20468 16974 20468 0 _0338_
rlabel metal1 11362 6324 11362 6324 0 _0339_
rlabel metal1 11684 5678 11684 5678 0 _0340_
rlabel metal1 18124 23222 18124 23222 0 _0341_
rlabel viali 12686 25874 12686 25874 0 _0342_
rlabel via2 14490 25789 14490 25789 0 _0343_
rlabel metal1 12351 24038 12351 24038 0 _0344_
rlabel metal1 16468 24582 16468 24582 0 _0345_
rlabel metal1 15640 25466 15640 25466 0 _0346_
rlabel metal1 16652 26554 16652 26554 0 _0347_
rlabel metal1 17204 24786 17204 24786 0 _0348_
rlabel metal2 17250 25908 17250 25908 0 _0349_
rlabel metal1 13846 25942 13846 25942 0 _0350_
rlabel metal1 14674 25364 14674 25364 0 _0351_
rlabel metal1 13938 25466 13938 25466 0 _0352_
rlabel metal1 14046 25194 14046 25194 0 _0353_
rlabel metal1 14444 24174 14444 24174 0 _0354_
rlabel metal1 12834 26350 12834 26350 0 _0355_
rlabel metal1 12512 24718 12512 24718 0 _0356_
rlabel metal1 12696 25942 12696 25942 0 _0357_
rlabel via1 12374 25891 12374 25891 0 _0358_
rlabel metal1 11592 24786 11592 24786 0 _0359_
rlabel metal2 11362 25398 11362 25398 0 _0360_
rlabel metal1 9890 24378 9890 24378 0 _0361_
rlabel metal1 9706 23528 9706 23528 0 _0362_
rlabel metal1 7958 23732 7958 23732 0 _0363_
rlabel metal1 10120 23698 10120 23698 0 _0364_
rlabel metal1 11270 23154 11270 23154 0 _0365_
rlabel metal1 10212 22678 10212 22678 0 _0366_
rlabel metal1 9752 21998 9752 21998 0 _0367_
rlabel metal1 11822 23120 11822 23120 0 _0368_
rlabel metal1 13432 23222 13432 23222 0 _0369_
rlabel metal2 12190 22916 12190 22916 0 _0370_
rlabel metal2 15318 8058 15318 8058 0 _0371_
rlabel metal1 15410 7956 15410 7956 0 _0372_
rlabel metal1 16054 4726 16054 4726 0 _0373_
rlabel metal2 3082 4454 3082 4454 0 _0374_
rlabel metal1 4048 6290 4048 6290 0 _0375_
rlabel metal1 5198 6766 5198 6766 0 _0376_
rlabel metal1 2530 3026 2530 3026 0 _0377_
rlabel metal1 5060 3162 5060 3162 0 _0378_
rlabel metal1 4002 3706 4002 3706 0 _0379_
rlabel metal1 2714 4556 2714 4556 0 _0380_
rlabel metal1 3680 4104 3680 4104 0 _0381_
rlabel metal1 3634 5134 3634 5134 0 _0382_
rlabel metal1 3220 4794 3220 4794 0 _0383_
rlabel viali 4520 6324 4520 6324 0 _0384_
rlabel metal1 3726 6324 3726 6324 0 _0385_
rlabel metal1 3726 5882 3726 5882 0 _0386_
rlabel metal1 3450 7514 3450 7514 0 _0387_
rlabel metal1 2530 7378 2530 7378 0 _0388_
rlabel metal1 4600 6426 4600 6426 0 _0389_
rlabel metal2 3634 7582 3634 7582 0 _0390_
rlabel metal1 3785 8534 3785 8534 0 _0391_
rlabel metal2 4002 8160 4002 8160 0 _0392_
rlabel metal2 2714 13158 2714 13158 0 _0393_
rlabel metal1 4784 11730 4784 11730 0 _0394_
rlabel via1 5395 13906 5395 13906 0 _0395_
rlabel metal2 2346 15028 2346 15028 0 _0396_
rlabel metal1 5106 13974 5106 13974 0 _0397_
rlabel metal1 2622 14008 2622 14008 0 _0398_
rlabel metal1 2392 13906 2392 13906 0 _0399_
rlabel metal1 2691 12886 2691 12886 0 _0400_
rlabel metal1 3818 12852 3818 12852 0 _0401_
rlabel metal1 2530 12716 2530 12716 0 _0402_
rlabel metal1 3802 11050 3802 11050 0 _0403_
rlabel metal1 3910 11798 3910 11798 0 _0404_
rlabel metal1 2990 11662 2990 11662 0 _0405_
rlabel metal1 3404 10778 3404 10778 0 _0406_
rlabel metal1 2484 10642 2484 10642 0 _0407_
rlabel metal1 4922 11322 4922 11322 0 _0408_
rlabel metal1 5060 11526 5060 11526 0 _0409_
rlabel metal1 5428 11118 5428 11118 0 _0410_
rlabel metal1 5198 11152 5198 11152 0 _0411_
rlabel metal1 7774 4556 7774 4556 0 _0412_
rlabel metal1 7912 8466 7912 8466 0 _0413_
rlabel metal2 7774 8908 7774 8908 0 _0414_
rlabel metal2 23828 15062 23828 15062 0 _0415_
rlabel metal2 24886 13311 24886 13311 0 _0416_
rlabel metal1 24104 14994 24104 14994 0 _0417_
rlabel metal1 23046 17850 23046 17850 0 _0418_
rlabel metal1 22632 17510 22632 17510 0 _0419_
rlabel metal1 23368 16218 23368 16218 0 _0420_
rlabel metal1 23414 16558 23414 16558 0 _0421_
rlabel metal1 25254 16218 25254 16218 0 _0422_
rlabel metal1 25576 15878 25576 15878 0 _0423_
rlabel metal1 25576 16558 25576 16558 0 _0424_
rlabel metal1 24794 13940 24794 13940 0 _0425_
rlabel metal1 23874 14994 23874 14994 0 _0426_
rlabel metal1 24610 15130 24610 15130 0 _0427_
rlabel metal1 24702 15504 24702 15504 0 _0428_
rlabel metal1 24472 14042 24472 14042 0 _0429_
rlabel metal1 23966 13294 23966 13294 0 _0430_
rlabel metal1 24978 13260 24978 13260 0 _0431_
rlabel metal2 25070 13056 25070 13056 0 _0432_
rlabel metal1 24656 13294 24656 13294 0 _0433_
rlabel metal1 25070 12954 25070 12954 0 _0434_
rlabel metal1 6026 15674 6026 15674 0 _0435_
rlabel metal1 3726 16558 3726 16558 0 _0436_
rlabel metal1 8694 11186 8694 11186 0 _0437_
rlabel metal1 8464 11050 8464 11050 0 _0438_
rlabel metal1 18308 11866 18308 11866 0 _0439_
rlabel metal1 19136 10234 19136 10234 0 _0440_
rlabel metal1 18860 8942 18860 8942 0 _0441_
rlabel metal1 12604 17306 12604 17306 0 _0442_
rlabel metal1 12137 19414 12137 19414 0 _0443_
rlabel metal1 8556 17646 8556 17646 0 _0444_
rlabel metal1 9121 18666 9121 18666 0 _0445_
rlabel metal1 11454 20570 11454 20570 0 _0446_
rlabel metal2 12190 18904 12190 18904 0 _0447_
rlabel metal1 11822 19312 11822 19312 0 _0448_
rlabel metal1 9890 19380 9890 19380 0 _0449_
rlabel metal1 9338 18836 9338 18836 0 _0450_
rlabel metal1 9108 19482 9108 19482 0 _0451_
rlabel metal2 9246 19380 9246 19380 0 _0452_
rlabel metal1 8786 20944 8786 20944 0 _0453_
rlabel metal1 7820 20434 7820 20434 0 _0454_
rlabel metal1 8740 19686 8740 19686 0 _0455_
rlabel metal2 8418 20332 8418 20332 0 _0456_
rlabel metal1 8510 18258 8510 18258 0 _0457_
rlabel metal1 8372 18802 8372 18802 0 _0458_
rlabel metal1 8050 19482 8050 19482 0 _0459_
rlabel metal1 8280 18394 8280 18394 0 _0460_
rlabel metal1 7544 18938 7544 18938 0 _0461_
rlabel metal2 19366 18037 19366 18037 0 _0462_
rlabel metal1 20424 16762 20424 16762 0 _0463_
rlabel metal1 20194 12852 20194 12852 0 _0464_
rlabel metal1 20332 12070 20332 12070 0 _0465_
rlabel metal1 13294 9894 13294 9894 0 _0466_
rlabel metal1 11914 8398 11914 8398 0 _0467_
rlabel metal1 12144 10438 12144 10438 0 _0468_
rlabel metal1 10948 8602 10948 8602 0 _0469_
rlabel metal1 19826 4046 19826 4046 0 _0470_
rlabel metal1 18170 4556 18170 4556 0 _0471_
rlabel metal1 11362 3060 11362 3060 0 _0472_
rlabel metal1 13432 4454 13432 4454 0 _0473_
rlabel metal1 13662 3094 13662 3094 0 _0474_
rlabel viali 14950 3025 14950 3025 0 _0475_
rlabel metal1 15558 4454 15558 4454 0 _0476_
rlabel metal1 16100 3026 16100 3026 0 _0477_
rlabel metal2 19826 4420 19826 4420 0 _0478_
rlabel metal1 18630 4590 18630 4590 0 _0479_
rlabel metal1 17526 4726 17526 4726 0 _0480_
rlabel metal2 15870 4998 15870 4998 0 _0481_
rlabel metal1 18630 4046 18630 4046 0 _0482_
rlabel metal1 17618 4624 17618 4624 0 _0483_
rlabel metal1 18998 4114 18998 4114 0 _0484_
rlabel metal2 18078 2587 18078 2587 0 _0485_
rlabel metal1 18768 2414 18768 2414 0 _0486_
rlabel metal1 19872 3502 19872 3502 0 _0487_
rlabel metal2 20010 3910 20010 3910 0 _0488_
rlabel metal1 14858 18326 14858 18326 0 _0489_
rlabel metal1 15548 20434 15548 20434 0 _0490_
rlabel metal1 12834 11866 12834 11866 0 _0491_
rlabel metal1 12742 12274 12742 12274 0 _0492_
rlabel metal1 19366 6358 19366 6358 0 _0493_
rlabel metal1 18860 7854 18860 7854 0 _0494_
rlabel metal1 20884 5202 20884 5202 0 _0495_
rlabel metal1 23644 4998 23644 4998 0 _0496_
rlabel metal1 23414 7888 23414 7888 0 _0497_
rlabel metal1 23460 7242 23460 7242 0 _0498_
rlabel metal1 21666 3026 21666 3026 0 _0499_
rlabel metal2 22034 4998 22034 4998 0 _0500_
rlabel metal2 23046 4318 23046 4318 0 _0501_
rlabel metal1 22916 4104 22916 4104 0 _0502_
rlabel metal1 24564 3434 24564 3434 0 _0503_
rlabel metal2 23966 4794 23966 4794 0 _0504_
rlabel metal1 24472 3502 24472 3502 0 _0505_
rlabel metal1 23322 8942 23322 8942 0 _0506_
rlabel metal1 24150 7174 24150 7174 0 _0507_
rlabel metal2 24334 8160 24334 8160 0 _0508_
rlabel metal2 23690 9418 23690 9418 0 _0509_
rlabel metal1 23184 9146 23184 9146 0 _0510_
rlabel metal1 23184 8058 23184 8058 0 _0511_
rlabel metal2 23598 8228 23598 8228 0 _0512_
rlabel metal1 24518 9554 24518 9554 0 _0513_
rlabel metal1 23782 8296 23782 8296 0 _0514_
rlabel metal1 23644 9078 23644 9078 0 _0515_
rlabel metal1 25392 9690 25392 9690 0 _0516_
rlabel metal1 16790 15470 16790 15470 0 _0517_
rlabel metal1 13984 15470 13984 15470 0 _0518_
rlabel metal1 8004 14382 8004 14382 0 _0519_
rlabel metal1 8372 3026 8372 3026 0 _0520_
rlabel metal2 13938 14314 13938 14314 0 clk
rlabel metal1 14628 9078 14628 9078 0 clknet_0_clk
rlabel metal1 1518 3434 1518 3434 0 clknet_4_0_0_clk
rlabel metal1 20516 8942 20516 8942 0 clknet_4_10_0_clk
rlabel metal1 19826 13838 19826 13838 0 clknet_4_11_0_clk
rlabel metal1 13846 15538 13846 15538 0 clknet_4_12_0_clk
rlabel metal1 13386 22066 13386 22066 0 clknet_4_13_0_clk
rlabel metal1 19320 19890 19320 19890 0 clknet_4_14_0_clk
rlabel metal1 19734 22644 19734 22644 0 clknet_4_15_0_clk
rlabel metal2 1886 8704 1886 8704 0 clknet_4_1_0_clk
rlabel metal1 8786 3978 8786 3978 0 clknet_4_2_0_clk
rlabel metal1 12926 12682 12926 12682 0 clknet_4_3_0_clk
rlabel metal1 1656 14926 1656 14926 0 clknet_4_4_0_clk
rlabel metal2 2438 16932 2438 16932 0 clknet_4_5_0_clk
rlabel metal1 14214 14348 14214 14348 0 clknet_4_6_0_clk
rlabel metal1 11362 25262 11362 25262 0 clknet_4_7_0_clk
rlabel metal2 17342 4352 17342 4352 0 clknet_4_8_0_clk
rlabel metal1 19366 13940 19366 13940 0 clknet_4_9_0_clk
rlabel metal1 6164 4114 6164 4114 0 conv1.addr\[8\]
rlabel metal1 12926 7854 12926 7854 0 conv1.done
rlabel metal1 7314 9486 7314 9486 0 conv1.psram_ce_n
rlabel metal1 3266 4012 3266 4012 0 conv1.psram_ctrl.counter\[0\]
rlabel viali 6669 4136 6669 4136 0 conv1.psram_ctrl.counter\[1\]
rlabel metal1 4462 3502 4462 3502 0 conv1.psram_ctrl.counter\[2\]
rlabel metal1 2622 4624 2622 4624 0 conv1.psram_ctrl.counter\[3\]
rlabel metal2 3174 6596 3174 6596 0 conv1.psram_ctrl.counter\[4\]
rlabel metal1 4002 8398 4002 8398 0 conv1.psram_ctrl.counter\[5\]
rlabel metal1 4646 7786 4646 7786 0 conv1.psram_ctrl.counter\[6\]
rlabel metal1 5474 7174 5474 7174 0 conv1.psram_ctrl.counter\[7\]
rlabel metal1 6900 5542 6900 5542 0 conv1.psram_ctrl.has_wait_states
rlabel metal1 8050 6868 8050 6868 0 conv1.psram_ctrl.nstate
rlabel via2 12926 8789 12926 8789 0 conv1.psram_ctrl.sck
rlabel metal1 8556 6426 8556 6426 0 conv1.psram_ctrl.start
rlabel metal1 7958 7242 7958 7242 0 conv1.psram_ctrl.state
rlabel metal1 8418 8874 8418 8874 0 conv1.state\[0\]
rlabel metal1 10304 4250 10304 4250 0 conv1.state\[1\]
rlabel metal1 8694 4590 8694 4590 0 conv1.state\[2\]
rlabel metal1 8004 8602 8004 8602 0 conv1.state\[3\]
rlabel metal1 8648 4250 8648 4250 0 conv1.state\[5\]
rlabel metal2 6394 15980 6394 15980 0 conv2.addr\[8\]
rlabel metal2 4922 16286 4922 16286 0 conv2.addr\[9\]
rlabel metal1 15640 14314 15640 14314 0 conv2.data_out_valid
rlabel metal1 8671 11526 8671 11526 0 conv2.psram_ce_n
rlabel metal1 2162 14416 2162 14416 0 conv2.psram_ctrl.counter\[0\]
rlabel metal1 2898 14314 2898 14314 0 conv2.psram_ctrl.counter\[1\]
rlabel metal1 1978 13940 1978 13940 0 conv2.psram_ctrl.counter\[2\]
rlabel metal1 5474 12716 5474 12716 0 conv2.psram_ctrl.counter\[3\]
rlabel metal2 3910 11968 3910 11968 0 conv2.psram_ctrl.counter\[4\]
rlabel metal1 5060 12206 5060 12206 0 conv2.psram_ctrl.counter\[5\]
rlabel metal1 5382 10676 5382 10676 0 conv2.psram_ctrl.counter\[6\]
rlabel metal1 6440 10574 6440 10574 0 conv2.psram_ctrl.counter\[7\]
rlabel metal1 7130 13702 7130 13702 0 conv2.psram_ctrl.has_wait_states
rlabel metal1 4830 16490 4830 16490 0 conv2.psram_ctrl.nstate
rlabel metal1 4186 13226 4186 13226 0 conv2.psram_ctrl.sck
rlabel metal1 5750 16218 5750 16218 0 conv2.psram_ctrl.start
rlabel metal1 6256 14382 6256 14382 0 conv2.psram_ctrl.state
rlabel metal1 11385 12138 11385 12138 0 conv2.state\[0\]
rlabel metal2 9706 15742 9706 15742 0 conv2.state\[1\]
rlabel metal2 8510 13821 8510 13821 0 conv2.state\[2\]
rlabel metal2 10350 13872 10350 13872 0 conv2.state\[3\]
rlabel metal1 8740 15538 8740 15538 0 conv2.state\[5\]
rlabel metal2 26174 1547 26174 1547 0 done
rlabel metal1 21160 17170 21160 17170 0 fc1.addr\[10\]
rlabel metal2 20746 18020 20746 18020 0 fc1.addr\[8\]
rlabel metal1 18446 13702 18446 13702 0 fc1.data_out_valid
rlabel metal1 21114 13328 21114 13328 0 fc1.psram_ce_n
rlabel metal1 23874 17646 23874 17646 0 fc1.psram_ctrl.counter\[0\]
rlabel metal1 24702 15980 24702 15980 0 fc1.psram_ctrl.counter\[1\]
rlabel metal1 24196 17646 24196 17646 0 fc1.psram_ctrl.counter\[2\]
rlabel metal2 24610 15980 24610 15980 0 fc1.psram_ctrl.counter\[3\]
rlabel metal1 22448 16558 22448 16558 0 fc1.psram_ctrl.counter\[4\]
rlabel metal1 24058 12920 24058 12920 0 fc1.psram_ctrl.counter\[5\]
rlabel metal1 24748 12750 24748 12750 0 fc1.psram_ctrl.counter\[6\]
rlabel metal1 25898 12818 25898 12818 0 fc1.psram_ctrl.counter\[7\]
rlabel metal1 19182 14926 19182 14926 0 fc1.psram_ctrl.has_wait_states
rlabel metal1 19734 15062 19734 15062 0 fc1.psram_ctrl.nstate
rlabel metal1 21712 12818 21712 12818 0 fc1.psram_ctrl.sck
rlabel metal1 21344 14382 21344 14382 0 fc1.psram_ctrl.start
rlabel metal2 21390 14620 21390 14620 0 fc1.psram_ctrl.state
rlabel metal1 17342 13294 17342 13294 0 fc1.state\[0\]
rlabel metal2 18446 17408 18446 17408 0 fc1.state\[1\]
rlabel metal1 19366 16116 19366 16116 0 fc1.state\[2\]
rlabel metal1 19274 13362 19274 13362 0 fc1.state\[3\]
rlabel metal1 18078 16626 18078 16626 0 fc1.state\[5\]
rlabel metal1 14812 19822 14812 19822 0 fc2.addr\[10\]
rlabel metal1 14996 19686 14996 19686 0 fc2.addr\[8\]
rlabel metal2 14122 13685 14122 13685 0 fc2.done
rlabel via1 13179 13158 13179 13158 0 fc2.psram_ce_n
rlabel metal2 13570 18496 13570 18496 0 fc2.psram_ctrl.counter\[0\]
rlabel metal1 13524 20434 13524 20434 0 fc2.psram_ctrl.counter\[1\]
rlabel metal2 12466 18632 12466 18632 0 fc2.psram_ctrl.counter\[2\]
rlabel metal2 11362 17952 11362 17952 0 fc2.psram_ctrl.counter\[3\]
rlabel metal1 9430 19856 9430 19856 0 fc2.psram_ctrl.counter\[4\]
rlabel metal1 11132 19142 11132 19142 0 fc2.psram_ctrl.counter\[5\]
rlabel metal1 9154 19312 9154 19312 0 fc2.psram_ctrl.counter\[6\]
rlabel metal1 8510 18768 8510 18768 0 fc2.psram_ctrl.counter\[7\]
rlabel metal1 10442 17102 10442 17102 0 fc2.psram_ctrl.has_wait_states
rlabel metal2 10902 15555 10902 15555 0 fc2.psram_ctrl.nstate
rlabel metal1 13202 12614 13202 12614 0 fc2.psram_ctrl.sck
rlabel metal1 12512 15538 12512 15538 0 fc2.psram_ctrl.start
rlabel metal1 12144 16694 12144 16694 0 fc2.psram_ctrl.state
rlabel metal1 14306 13702 14306 13702 0 fc2.state\[0\]
rlabel metal1 15456 15674 15456 15674 0 fc2.state\[1\]
rlabel metal2 15318 15164 15318 15164 0 fc2.state\[2\]
rlabel metal1 15548 14382 15548 14382 0 fc2.state\[3\]
rlabel metal1 14030 16626 14030 16626 0 fc2.state\[5\]
rlabel metal1 13064 6086 13064 6086 0 maxpool.addr\[11\]
rlabel metal2 12006 7412 12006 7412 0 maxpool.addr\[8\]
rlabel metal2 16054 9044 16054 9044 0 maxpool.psram_ce_n
rlabel metal2 14122 2992 14122 2992 0 maxpool.psram_ctrl.counter\[0\]
rlabel metal1 14536 2414 14536 2414 0 maxpool.psram_ctrl.counter\[1\]
rlabel metal2 13294 3196 13294 3196 0 maxpool.psram_ctrl.counter\[2\]
rlabel metal1 15686 4590 15686 4590 0 maxpool.psram_ctrl.counter\[3\]
rlabel metal1 16192 5134 16192 5134 0 maxpool.psram_ctrl.counter\[4\]
rlabel metal1 16698 4590 16698 4590 0 maxpool.psram_ctrl.counter\[5\]
rlabel metal2 19366 3706 19366 3706 0 maxpool.psram_ctrl.counter\[6\]
rlabel metal1 17848 2890 17848 2890 0 maxpool.psram_ctrl.counter\[7\]
rlabel metal1 13110 5814 13110 5814 0 maxpool.psram_ctrl.nstate
rlabel metal1 16330 4658 16330 4658 0 maxpool.psram_ctrl.sck
rlabel metal1 14122 6290 14122 6290 0 maxpool.psram_ctrl.start
rlabel metal1 14444 6834 14444 6834 0 maxpool.psram_ctrl.state
rlabel metal1 13110 10064 13110 10064 0 maxpool.state\[0\]
rlabel metal1 12926 9894 12926 9894 0 maxpool.state\[1\]
rlabel metal1 11454 9894 11454 9894 0 maxpool.state\[2\]
rlabel metal1 21436 21522 21436 21522 0 mfcc.dct.data_valid
rlabel metal1 21666 19924 21666 19924 0 mfcc.dct.dct_valid
rlabel metal2 21114 25092 21114 25092 0 mfcc.dct.input_counter\[0\]
rlabel metal1 20516 25126 20516 25126 0 mfcc.dct.input_counter\[1\]
rlabel metal1 19964 25670 19964 25670 0 mfcc.dct.input_counter\[2\]
rlabel metal2 21850 26452 21850 26452 0 mfcc.dct.input_counter\[3\]
rlabel metal1 22586 25466 22586 25466 0 mfcc.dct.input_counter\[4\]
rlabel metal2 23322 24004 23322 24004 0 mfcc.dct.output_counter\[0\]
rlabel metal1 24600 22610 24600 22610 0 mfcc.dct.output_counter\[1\]
rlabel via1 24518 22763 24518 22763 0 mfcc.dct.output_counter\[2\]
rlabel metal2 23414 20604 23414 20604 0 mfcc.dct.output_counter\[3\]
rlabel metal1 23690 20910 23690 20910 0 mfcc.dct.output_counter\[4\]
rlabel metal1 23138 20910 23138 20910 0 mfcc.dct.output_counter\[5\]
rlabel metal1 20654 23154 20654 23154 0 mfcc.dct.state\[0\]
rlabel metal1 20792 22746 20792 22746 0 mfcc.dct.state\[1\]
rlabel metal1 15778 21522 15778 21522 0 mfcc.log.data_valid
rlabel metal1 18308 22134 18308 22134 0 mfcc.log.shift_count\[0\]
rlabel metal1 16882 20026 16882 20026 0 mfcc.log.shift_count\[1\]
rlabel metal2 18446 19856 18446 19856 0 mfcc.log.shift_count\[2\]
rlabel metal1 18906 20434 18906 20434 0 mfcc.log.shift_count\[3\]
rlabel metal1 15916 21658 15916 21658 0 mfcc.log.state\[0\]
rlabel metal1 17894 21658 17894 21658 0 mfcc.log.state\[1\]
rlabel metal2 16192 21522 16192 21522 0 mfcc.log.state\[2\]
rlabel metal2 9614 24548 9614 24548 0 mfcc.mel.coeff_counter\[0\]
rlabel metal1 10166 23256 10166 23256 0 mfcc.mel.coeff_counter\[1\]
rlabel metal1 9706 23018 9706 23018 0 mfcc.mel.coeff_counter\[2\]
rlabel metal1 11362 22542 11362 22542 0 mfcc.mel.coeff_counter\[3\]
rlabel metal1 13386 23052 13386 23052 0 mfcc.mel.coeff_counter\[4\]
rlabel metal1 16192 26418 16192 26418 0 mfcc.mel.filter_counter\[0\]
rlabel metal1 16744 26010 16744 26010 0 mfcc.mel.filter_counter\[1\]
rlabel metal1 17986 25466 17986 25466 0 mfcc.mel.filter_counter\[2\]
rlabel metal1 15870 25942 15870 25942 0 mfcc.mel.filter_counter\[3\]
rlabel metal1 12834 24684 12834 24684 0 mfcc.mel.filter_counter\[4\]
rlabel metal1 12144 25126 12144 25126 0 mfcc.mel.filter_counter\[5\]
rlabel metal2 11822 24956 11822 24956 0 mfcc.mel.state\[0\]
rlabel metal2 9890 25432 9890 25432 0 mfcc.mel.state\[1\]
rlabel metal2 20148 16660 20148 16660 0 mfcc.mfcc_valid
rlabel metal1 14766 15368 14766 15368 0 net1
rlabel metal2 12926 4862 12926 4862 0 net10
rlabel metal1 24794 6324 24794 6324 0 net100
rlabel viali 14489 4182 14489 4182 0 net101
rlabel metal1 13386 4046 13386 4046 0 net102
rlabel metal1 3220 11730 3220 11730 0 net103
rlabel metal1 22632 23698 22632 23698 0 net104
rlabel metal1 16652 24786 16652 24786 0 net105
rlabel metal1 18584 14518 18584 14518 0 net106
rlabel metal1 17526 14586 17526 14586 0 net107
rlabel metal1 18170 13498 18170 13498 0 net108
rlabel metal1 7544 19482 7544 19482 0 net109
rlabel metal2 6946 17612 6946 17612 0 net11
rlabel metal1 22494 21556 22494 21556 0 net110
rlabel metal1 16238 13940 16238 13940 0 net111
rlabel metal1 17250 13362 17250 13362 0 net112
rlabel metal1 6670 15062 6670 15062 0 net113
rlabel metal1 7826 16762 7826 16762 0 net114
rlabel metal1 14398 25772 14398 25772 0 net115
rlabel metal1 12098 15130 12098 15130 0 net116
rlabel metal1 22356 14994 22356 14994 0 net117
rlabel metal2 22126 17714 22126 17714 0 net118
rlabel metal1 19964 26350 19964 26350 0 net119
rlabel metal1 10120 22610 10120 22610 0 net12
rlabel metal1 18768 23086 18768 23086 0 net120
rlabel metal1 18901 22610 18901 22610 0 net121
rlabel metal1 4186 16456 4186 16456 0 net122
rlabel metal1 16790 5270 16790 5270 0 net123
rlabel metal1 5704 17578 5704 17578 0 net124
rlabel metal1 18722 15504 18722 15504 0 net125
rlabel metal1 15226 20026 15226 20026 0 net126
rlabel metal1 13018 24174 13018 24174 0 net127
rlabel metal2 13386 5984 13386 5984 0 net128
rlabel metal1 10258 11730 10258 11730 0 net129
rlabel metal1 12611 19754 12611 19754 0 net13
rlabel metal1 13018 16626 13018 16626 0 net130
rlabel metal1 14674 6426 14674 6426 0 net131
rlabel metal1 12282 16694 12282 16694 0 net132
rlabel metal2 12926 19482 12926 19482 0 net133
rlabel metal1 5704 4046 5704 4046 0 net134
rlabel metal2 21850 6902 21850 6902 0 net135
rlabel metal1 16514 8466 16514 8466 0 net136
rlabel metal1 24104 3570 24104 3570 0 net137
rlabel metal1 12282 8500 12282 8500 0 net138
rlabel metal1 18676 2482 18676 2482 0 net139
rlabel metal2 12466 13566 12466 13566 0 net14
rlabel metal1 17710 3162 17710 3162 0 net140
rlabel metal1 25208 9622 25208 9622 0 net141
rlabel metal1 17526 11186 17526 11186 0 net142
rlabel metal1 20470 16558 20470 16558 0 net143
rlabel metal1 12466 18666 12466 18666 0 net144
rlabel metal1 9246 24378 9246 24378 0 net145
rlabel metal1 22356 5270 22356 5270 0 net146
rlabel metal1 7498 8976 7498 8976 0 net147
rlabel metal1 9844 8398 9844 8398 0 net148
rlabel metal1 9752 18734 9752 18734 0 net149
rlabel metal2 18722 3298 18722 3298 0 net15
rlabel metal1 8694 3060 8694 3060 0 net150
rlabel metal1 3082 12750 3082 12750 0 net151
rlabel metal1 15318 3060 15318 3060 0 net152
rlabel metal1 14214 3026 14214 3026 0 net153
rlabel metal1 7360 12954 7360 12954 0 net154
rlabel metal1 19090 9962 19090 9962 0 net155
rlabel viali 23782 16559 23782 16559 0 net156
rlabel metal1 4232 4046 4232 4046 0 net157
rlabel metal1 19734 24208 19734 24208 0 net158
rlabel metal1 25898 16626 25898 16626 0 net159
rlabel metal2 21942 4046 21942 4046 0 net16
rlabel metal1 24012 3638 24012 3638 0 net160
rlabel metal1 12052 7514 12052 7514 0 net161
rlabel metal1 9016 19754 9016 19754 0 net162
rlabel metal1 25162 15334 25162 15334 0 net163
rlabel metal1 17710 15334 17710 15334 0 net164
rlabel metal1 7682 20332 7682 20332 0 net165
rlabel metal1 8694 13498 8694 13498 0 net166
rlabel metal1 19366 6086 19366 6086 0 net167
rlabel metal1 20884 26554 20884 26554 0 net168
rlabel metal2 21942 12517 21942 12517 0 net17
rlabel metal1 14674 7888 14674 7888 0 net18
rlabel metal2 14858 17000 14858 17000 0 net19
rlabel metal1 21275 11798 21275 11798 0 net2
rlabel metal1 14911 19346 14911 19346 0 net20
rlabel metal2 20562 19346 20562 19346 0 net21
rlabel metal2 21206 16286 21206 16286 0 net22
rlabel metal1 3956 26962 3956 26962 0 net23
rlabel metal1 26358 4998 26358 4998 0 net24
rlabel metal2 10350 1027 10350 1027 0 net25
rlabel metal2 26174 23953 26174 23953 0 net26
rlabel metal2 11086 27251 11086 27251 0 net27
rlabel metal1 14904 26962 14904 26962 0 net28
rlabel metal3 820 26588 820 26588 0 net29
rlabel metal1 20286 9894 20286 9894 0 net3
rlabel metal1 21022 20026 21022 20026 0 net30
rlabel metal2 7314 14246 7314 14246 0 net31
rlabel metal1 21942 6732 21942 6732 0 net32
rlabel metal1 19780 6358 19780 6358 0 net33
rlabel metal1 10212 14994 10212 14994 0 net34
rlabel metal1 7958 16184 7958 16184 0 net35
rlabel metal1 18538 17646 18538 17646 0 net36
rlabel metal1 17112 17238 17112 17238 0 net37
rlabel metal1 13248 15470 13248 15470 0 net38
rlabel metal1 14306 15538 14306 15538 0 net39
rlabel metal1 1978 18394 1978 18394 0 net4
rlabel metal2 10350 4318 10350 4318 0 net40
rlabel metal1 9108 2618 9108 2618 0 net41
rlabel metal1 20746 13294 20746 13294 0 net42
rlabel metal1 11868 13906 11868 13906 0 net43
rlabel metal1 15824 6766 15824 6766 0 net44
rlabel metal1 13110 13940 13110 13940 0 net45
rlabel metal1 14076 12818 14076 12818 0 net46
rlabel metal1 6808 7378 6808 7378 0 net47
rlabel metal1 10580 26214 10580 26214 0 net48
rlabel metal2 21758 26112 21758 26112 0 net49
rlabel metal1 18630 2346 18630 2346 0 net5
rlabel metal1 23874 20502 23874 20502 0 net50
rlabel metal1 17342 20332 17342 20332 0 net51
rlabel metal1 21436 8466 21436 8466 0 net52
rlabel via1 16414 21930 16414 21930 0 net53
rlabel metal1 14899 21522 14899 21522 0 net54
rlabel metal2 10074 8432 10074 8432 0 net55
rlabel metal1 9936 9146 9936 9146 0 net56
rlabel metal1 25070 21998 25070 21998 0 net57
rlabel metal2 11638 8670 11638 8670 0 net58
rlabel metal1 12742 23086 12742 23086 0 net59
rlabel metal1 13294 10064 13294 10064 0 net6
rlabel metal1 4324 7922 4324 7922 0 net60
rlabel metal2 2898 8364 2898 8364 0 net61
rlabel metal1 24380 12750 24380 12750 0 net62
rlabel metal1 24610 21522 24610 21522 0 net63
rlabel metal1 4784 10574 4784 10574 0 net64
rlabel metal1 3864 9486 3864 9486 0 net65
rlabel metal2 17526 26792 17526 26792 0 net66
rlabel via2 18538 20587 18538 20587 0 net67
rlabel metal1 19596 24922 19596 24922 0 net68
rlabel metal1 10442 14994 10442 14994 0 net69
rlabel metal1 6263 3434 6263 3434 0 net7
rlabel metal1 15548 14246 15548 14246 0 net70
rlabel metal1 14536 13498 14536 13498 0 net71
rlabel metal1 21206 26996 21206 26996 0 net72
rlabel metal1 14720 23630 14720 23630 0 net73
rlabel metal1 9016 13430 9016 13430 0 net74
rlabel metal1 8740 13974 8740 13974 0 net75
rlabel metal1 13662 22202 13662 22202 0 net76
rlabel metal1 19734 16082 19734 16082 0 net77
rlabel metal1 19366 17272 19366 17272 0 net78
rlabel metal1 13018 13192 13018 13192 0 net79
rlabel metal1 6723 9962 6723 9962 0 net8
rlabel metal1 9844 11866 9844 11866 0 net80
rlabel metal1 20654 7514 20654 7514 0 net81
rlabel metal1 18630 21624 18630 21624 0 net82
rlabel metal1 5428 11050 5428 11050 0 net83
rlabel metal1 7360 4250 7360 4250 0 net84
rlabel metal1 7912 3094 7912 3094 0 net85
rlabel metal1 25116 12886 25116 12886 0 net86
rlabel metal1 16192 17170 16192 17170 0 net87
rlabel metal1 15318 18394 15318 18394 0 net88
rlabel metal1 9062 6698 9062 6698 0 net89
rlabel metal1 8694 4073 8694 4073 0 net9
rlabel metal1 7820 5134 7820 5134 0 net90
rlabel metal1 8556 5610 8556 5610 0 net91
rlabel metal1 20792 14314 20792 14314 0 net92
rlabel metal1 3726 6426 3726 6426 0 net93
rlabel metal1 10626 3094 10626 3094 0 net94
rlabel metal1 4462 8602 4462 8602 0 net95
rlabel metal1 17434 19482 17434 19482 0 net96
rlabel metal1 17020 20366 17020 20366 0 net97
rlabel viali 21758 23086 21758 23086 0 net98
rlabel via1 21026 21998 21026 21998 0 net99
rlabel metal3 820 19108 820 19108 0 psram_ce_n
rlabel metal1 4738 2822 4738 2822 0 psram_d[0]
rlabel metal2 18078 1520 18078 1520 0 psram_sck
rlabel metal3 751 15028 751 15028 0 rst_n
rlabel metal1 21528 5814 21528 5814 0 softmax.addr\[11\]
rlabel metal1 21574 6358 21574 6358 0 softmax.addr\[8\]
rlabel metal1 19872 6834 19872 6834 0 softmax.data_valid
rlabel metal1 21022 9588 21022 9588 0 softmax.psram_ce_n
rlabel metal1 23690 4012 23690 4012 0 softmax.psram_ctrl.counter\[0\]
rlabel metal1 24334 5270 24334 5270 0 softmax.psram_ctrl.counter\[1\]
rlabel metal2 23506 6426 23506 6426 0 softmax.psram_ctrl.counter\[2\]
rlabel metal1 25116 5882 25116 5882 0 softmax.psram_ctrl.counter\[3\]
rlabel metal1 24932 7378 24932 7378 0 softmax.psram_ctrl.counter\[4\]
rlabel metal1 24150 9010 24150 9010 0 softmax.psram_ctrl.counter\[5\]
rlabel metal1 25760 8602 25760 8602 0 softmax.psram_ctrl.counter\[6\]
rlabel metal1 25024 7174 25024 7174 0 softmax.psram_ctrl.counter\[7\]
rlabel metal1 20884 7786 20884 7786 0 softmax.psram_ctrl.nstate
rlabel metal1 17894 8976 17894 8976 0 softmax.psram_ctrl.sck
rlabel metal2 19918 8126 19918 8126 0 softmax.psram_ctrl.start
rlabel metal2 22402 7514 22402 7514 0 softmax.psram_ctrl.state
rlabel metal3 26550 12308 26550 12308 0 start
rlabel metal1 21022 11662 21022 11662 0 state\[0\]
rlabel metal2 19642 11968 19642 11968 0 state\[1\]
rlabel metal1 18952 11118 18952 11118 0 state\[2\]
<< properties >>
string FIXED_BBOX 0 0 27641 29785
<< end >>
