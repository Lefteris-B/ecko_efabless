VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cnn_kws_accel
  CLASS BLOCK ;
  FOREIGN cnn_kws_accel ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN audio_sample[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 231.240 350.000 231.840 ;
    END
  END audio_sample[0]
  PIN audio_sample[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END audio_sample[10]
  PIN audio_sample[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END audio_sample[11]
  PIN audio_sample[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 187.040 350.000 187.640 ;
    END
  END audio_sample[12]
  PIN audio_sample[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 346.000 238.650 350.000 ;
    END
  END audio_sample[13]
  PIN audio_sample[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END audio_sample[14]
  PIN audio_sample[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END audio_sample[15]
  PIN audio_sample[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 326.440 350.000 327.040 ;
    END
  END audio_sample[1]
  PIN audio_sample[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 346.000 283.730 350.000 ;
    END
  END audio_sample[2]
  PIN audio_sample[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 91.840 350.000 92.440 ;
    END
  END audio_sample[3]
  PIN audio_sample[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END audio_sample[4]
  PIN audio_sample[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END audio_sample[5]
  PIN audio_sample[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 346.000 328.810 350.000 ;
    END
  END audio_sample[6]
  PIN audio_sample[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END audio_sample[7]
  PIN audio_sample[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 346.000 106.630 350.000 ;
    END
  END audio_sample[8]
  PIN audio_sample[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END audio_sample[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 0.040 350.000 0.640 ;
    END
  END done
  PIN psram_ce_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END psram_ce_n
  PIN psram_d[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END psram_d[0]
  PIN psram_d[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 346.000 64.770 350.000 ;
    END
  END psram_d[1]
  PIN psram_d[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 47.640 350.000 48.240 ;
    END
  END psram_d[2]
  PIN psram_d[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END psram_d[3]
  PIN psram_douten[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END psram_douten[0]
  PIN psram_douten[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 278.840 350.000 279.440 ;
    END
  END psram_douten[1]
  PIN psram_douten[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 346.000 151.710 350.000 ;
    END
  END psram_douten[2]
  PIN psram_douten[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 346.000 196.790 350.000 ;
    END
  END psram_douten[3]
  PIN psram_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END psram_sck
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END rst
  PIN sample_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 346.000 19.690 350.000 ;
    END
  END sample_valid
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 346.000 139.440 350.000 140.040 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 4.670 10.640 344.470 337.520 ;
      LAYER met2 ;
        RECT 4.690 345.720 19.130 346.530 ;
        RECT 19.970 345.720 64.210 346.530 ;
        RECT 65.050 345.720 106.070 346.530 ;
        RECT 106.910 345.720 151.150 346.530 ;
        RECT 151.990 345.720 196.230 346.530 ;
        RECT 197.070 345.720 238.090 346.530 ;
        RECT 238.930 345.720 283.170 346.530 ;
        RECT 284.010 345.720 328.250 346.530 ;
        RECT 329.090 345.720 344.450 346.530 ;
        RECT 4.690 4.280 344.450 345.720 ;
        RECT 4.690 0.155 41.670 4.280 ;
        RECT 42.510 0.155 86.750 4.280 ;
        RECT 87.590 0.155 131.830 4.280 ;
        RECT 132.670 0.155 173.690 4.280 ;
        RECT 174.530 0.155 218.770 4.280 ;
        RECT 219.610 0.155 263.850 4.280 ;
        RECT 264.690 0.155 305.710 4.280 ;
        RECT 306.550 0.155 344.450 4.280 ;
      LAYER met3 ;
        RECT 3.990 327.440 346.000 337.445 ;
        RECT 3.990 326.040 345.600 327.440 ;
        RECT 3.990 324.040 346.000 326.040 ;
        RECT 4.400 322.640 346.000 324.040 ;
        RECT 3.990 279.840 346.000 322.640 ;
        RECT 4.400 278.440 345.600 279.840 ;
        RECT 3.990 232.240 346.000 278.440 ;
        RECT 4.400 230.840 345.600 232.240 ;
        RECT 3.990 188.040 346.000 230.840 ;
        RECT 3.990 186.640 345.600 188.040 ;
        RECT 3.990 184.640 346.000 186.640 ;
        RECT 4.400 183.240 346.000 184.640 ;
        RECT 3.990 140.440 346.000 183.240 ;
        RECT 4.400 139.040 345.600 140.440 ;
        RECT 3.990 92.840 346.000 139.040 ;
        RECT 4.400 91.440 345.600 92.840 ;
        RECT 3.990 48.640 346.000 91.440 ;
        RECT 3.990 47.240 345.600 48.640 ;
        RECT 3.990 45.240 346.000 47.240 ;
        RECT 4.400 43.840 346.000 45.240 ;
        RECT 3.990 1.040 346.000 43.840 ;
        RECT 3.990 0.175 345.600 1.040 ;
  END
END cnn_kws_accel
END LIBRARY

